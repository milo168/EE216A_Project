`define CLOG2(x) \
(x <= 2) ? 1 : \
(x <= 4) ? 2 : \
(x <= 8) ? 3 : \
(x <= 16) ? 4 : \
(x <= 32) ? 5 : \
(x <= 64) ? 6 : \
(x <= 128) ? 7 : \
(x <= 256) ? 8 : \
(x <= 512) ? 9 : \
(x <= 1024) ? 10 : \
-1

module Image_Classifier
(
	clk,
	GlobalReset,
	Input_Valid,
	Wgt_0_0,Wgt_0_1,Wgt_0_2,Wgt_0_3,Wgt_0_4,Wgt_0_5,Wgt_0_6,Wgt_0_7,Wgt_0_8,Wgt_0_9,Wgt_0_10,Wgt_0_11,Wgt_0_12,Wgt_0_13,Wgt_0_14,Wgt_0_15,Wgt_0_16,Wgt_0_17,Wgt_0_18,Wgt_0_19,Wgt_0_20,Wgt_0_21,Wgt_0_22,Wgt_0_23,Wgt_0_24,Wgt_0_25,Wgt_0_26,Wgt_0_27,Wgt_0_28,Wgt_0_29,Wgt_0_30,Wgt_0_31,Wgt_0_32,Wgt_0_33,Wgt_0_34,Wgt_0_35,Wgt_0_36,Wgt_0_37,Wgt_0_38,Wgt_0_39,Wgt_0_40,Wgt_0_41,Wgt_0_42,Wgt_0_43,Wgt_0_44,Wgt_0_45,Wgt_0_46,Wgt_0_47,Wgt_0_48,Wgt_0_49,Wgt_0_50,Wgt_0_51,Wgt_0_52,Wgt_0_53,Wgt_0_54,Wgt_0_55,Wgt_0_56,Wgt_0_57,Wgt_0_58,Wgt_0_59,Wgt_0_60,Wgt_0_61,Wgt_0_62,Wgt_0_63,Wgt_0_64,Wgt_0_65,Wgt_0_66,Wgt_0_67,Wgt_0_68,Wgt_0_69,Wgt_0_70,Wgt_0_71,Wgt_0_72,Wgt_0_73,Wgt_0_74,Wgt_0_75,Wgt_0_76,Wgt_0_77,Wgt_0_78,Wgt_0_79,Wgt_0_80,Wgt_0_81,Wgt_0_82,Wgt_0_83,Wgt_0_84,Wgt_0_85,Wgt_0_86,Wgt_0_87,Wgt_0_88,Wgt_0_89,Wgt_0_90,Wgt_0_91,Wgt_0_92,Wgt_0_93,Wgt_0_94,Wgt_0_95,Wgt_0_96,Wgt_0_97,Wgt_0_98,Wgt_0_99,Wgt_0_100,Wgt_0_101,Wgt_0_102,Wgt_0_103,Wgt_0_104,Wgt_0_105,Wgt_0_106,Wgt_0_107,Wgt_0_108,Wgt_0_109,Wgt_0_110,Wgt_0_111,Wgt_0_112,Wgt_0_113,Wgt_0_114,Wgt_0_115,Wgt_0_116,Wgt_0_117,Wgt_0_118,Wgt_0_119,Wgt_0_120,Wgt_0_121,Wgt_0_122,Wgt_0_123,Wgt_0_124,Wgt_0_125,Wgt_0_126,Wgt_0_127,Wgt_0_128,Wgt_0_129,Wgt_0_130,Wgt_0_131,Wgt_0_132,Wgt_0_133,Wgt_0_134,Wgt_0_135,Wgt_0_136,Wgt_0_137,Wgt_0_138,Wgt_0_139,Wgt_0_140,Wgt_0_141,Wgt_0_142,Wgt_0_143,Wgt_0_144,Wgt_0_145,Wgt_0_146,Wgt_0_147,Wgt_0_148,Wgt_0_149,Wgt_0_150,Wgt_0_151,Wgt_0_152,Wgt_0_153,Wgt_0_154,Wgt_0_155,Wgt_0_156,Wgt_0_157,Wgt_0_158,Wgt_0_159,Wgt_0_160,Wgt_0_161,Wgt_0_162,Wgt_0_163,Wgt_0_164,Wgt_0_165,Wgt_0_166,Wgt_0_167,Wgt_0_168,Wgt_0_169,Wgt_0_170,Wgt_0_171,Wgt_0_172,Wgt_0_173,Wgt_0_174,Wgt_0_175,Wgt_0_176,Wgt_0_177,Wgt_0_178,Wgt_0_179,Wgt_0_180,Wgt_0_181,Wgt_0_182,Wgt_0_183,Wgt_0_184,Wgt_0_185,Wgt_0_186,Wgt_0_187,Wgt_0_188,Wgt_0_189,Wgt_0_190,Wgt_0_191,Wgt_0_192,Wgt_0_193,Wgt_0_194,Wgt_0_195,Wgt_0_196,Wgt_0_197,Wgt_0_198,Wgt_0_199,Wgt_0_200,Wgt_0_201,Wgt_0_202,Wgt_0_203,Wgt_0_204,Wgt_0_205,Wgt_0_206,Wgt_0_207,Wgt_0_208,Wgt_0_209,Wgt_0_210,Wgt_0_211,Wgt_0_212,Wgt_0_213,Wgt_0_214,Wgt_0_215,Wgt_0_216,Wgt_0_217,Wgt_0_218,Wgt_0_219,Wgt_0_220,Wgt_0_221,Wgt_0_222,Wgt_0_223,Wgt_0_224,Wgt_0_225,Wgt_0_226,Wgt_0_227,Wgt_0_228,Wgt_0_229,Wgt_0_230,Wgt_0_231,Wgt_0_232,Wgt_0_233,Wgt_0_234,Wgt_0_235,Wgt_0_236,Wgt_0_237,Wgt_0_238,Wgt_0_239,Wgt_0_240,Wgt_0_241,Wgt_0_242,Wgt_0_243,Wgt_0_244,Wgt_0_245,Wgt_0_246,Wgt_0_247,Wgt_0_248,Wgt_0_249,Wgt_0_250,Wgt_0_251,Wgt_0_252,Wgt_0_253,Wgt_0_254,Wgt_0_255,Wgt_0_256,Wgt_0_257,Wgt_0_258,Wgt_0_259,Wgt_0_260,Wgt_0_261,Wgt_0_262,Wgt_0_263,Wgt_0_264,Wgt_0_265,Wgt_0_266,Wgt_0_267,Wgt_0_268,Wgt_0_269,Wgt_0_270,Wgt_0_271,Wgt_0_272,Wgt_0_273,Wgt_0_274,Wgt_0_275,Wgt_0_276,Wgt_0_277,Wgt_0_278,Wgt_0_279,Wgt_0_280,Wgt_0_281,Wgt_0_282,Wgt_0_283,Wgt_0_284,Wgt_0_285,Wgt_0_286,Wgt_0_287,Wgt_0_288,Wgt_0_289,Wgt_0_290,Wgt_0_291,Wgt_0_292,Wgt_0_293,Wgt_0_294,Wgt_0_295,Wgt_0_296,Wgt_0_297,Wgt_0_298,Wgt_0_299,Wgt_0_300,Wgt_0_301,Wgt_0_302,Wgt_0_303,Wgt_0_304,Wgt_0_305,Wgt_0_306,Wgt_0_307,Wgt_0_308,Wgt_0_309,Wgt_0_310,Wgt_0_311,Wgt_0_312,Wgt_0_313,Wgt_0_314,Wgt_0_315,Wgt_0_316,Wgt_0_317,Wgt_0_318,Wgt_0_319,Wgt_0_320,Wgt_0_321,Wgt_0_322,Wgt_0_323,Wgt_0_324,Wgt_0_325,Wgt_0_326,Wgt_0_327,Wgt_0_328,Wgt_0_329,Wgt_0_330,Wgt_0_331,Wgt_0_332,Wgt_0_333,Wgt_0_334,Wgt_0_335,Wgt_0_336,Wgt_0_337,Wgt_0_338,Wgt_0_339,Wgt_0_340,Wgt_0_341,Wgt_0_342,Wgt_0_343,Wgt_0_344,Wgt_0_345,Wgt_0_346,Wgt_0_347,Wgt_0_348,Wgt_0_349,Wgt_0_350,Wgt_0_351,Wgt_0_352,Wgt_0_353,Wgt_0_354,Wgt_0_355,Wgt_0_356,Wgt_0_357,Wgt_0_358,Wgt_0_359,Wgt_0_360,Wgt_0_361,Wgt_0_362,Wgt_0_363,Wgt_0_364,Wgt_0_365,Wgt_0_366,Wgt_0_367,Wgt_0_368,Wgt_0_369,Wgt_0_370,Wgt_0_371,Wgt_0_372,Wgt_0_373,Wgt_0_374,Wgt_0_375,Wgt_0_376,Wgt_0_377,Wgt_0_378,Wgt_0_379,Wgt_0_380,Wgt_0_381,Wgt_0_382,Wgt_0_383,Wgt_0_384,Wgt_0_385,Wgt_0_386,Wgt_0_387,Wgt_0_388,Wgt_0_389,Wgt_0_390,Wgt_0_391,Wgt_0_392,Wgt_0_393,Wgt_0_394,Wgt_0_395,Wgt_0_396,Wgt_0_397,Wgt_0_398,Wgt_0_399,Wgt_0_400,Wgt_0_401,Wgt_0_402,Wgt_0_403,Wgt_0_404,Wgt_0_405,Wgt_0_406,Wgt_0_407,Wgt_0_408,Wgt_0_409,Wgt_0_410,Wgt_0_411,Wgt_0_412,Wgt_0_413,Wgt_0_414,Wgt_0_415,Wgt_0_416,Wgt_0_417,Wgt_0_418,Wgt_0_419,Wgt_0_420,Wgt_0_421,Wgt_0_422,Wgt_0_423,Wgt_0_424,Wgt_0_425,Wgt_0_426,Wgt_0_427,Wgt_0_428,Wgt_0_429,Wgt_0_430,Wgt_0_431,Wgt_0_432,Wgt_0_433,Wgt_0_434,Wgt_0_435,Wgt_0_436,Wgt_0_437,Wgt_0_438,Wgt_0_439,Wgt_0_440,Wgt_0_441,Wgt_0_442,Wgt_0_443,Wgt_0_444,Wgt_0_445,Wgt_0_446,Wgt_0_447,Wgt_0_448,Wgt_0_449,Wgt_0_450,Wgt_0_451,Wgt_0_452,Wgt_0_453,Wgt_0_454,Wgt_0_455,Wgt_0_456,Wgt_0_457,Wgt_0_458,Wgt_0_459,Wgt_0_460,Wgt_0_461,Wgt_0_462,Wgt_0_463,Wgt_0_464,Wgt_0_465,Wgt_0_466,Wgt_0_467,Wgt_0_468,Wgt_0_469,Wgt_0_470,Wgt_0_471,Wgt_0_472,Wgt_0_473,Wgt_0_474,Wgt_0_475,Wgt_0_476,Wgt_0_477,Wgt_0_478,Wgt_0_479,Wgt_0_480,Wgt_0_481,Wgt_0_482,Wgt_0_483,Wgt_0_484,Wgt_0_485,Wgt_0_486,Wgt_0_487,Wgt_0_488,Wgt_0_489,Wgt_0_490,Wgt_0_491,Wgt_0_492,Wgt_0_493,Wgt_0_494,Wgt_0_495,Wgt_0_496,Wgt_0_497,Wgt_0_498,Wgt_0_499,Wgt_0_500,Wgt_0_501,Wgt_0_502,Wgt_0_503,Wgt_0_504,Wgt_0_505,Wgt_0_506,Wgt_0_507,Wgt_0_508,Wgt_0_509,Wgt_0_510,Wgt_0_511,Wgt_0_512,Wgt_0_513,Wgt_0_514,Wgt_0_515,Wgt_0_516,Wgt_0_517,Wgt_0_518,Wgt_0_519,Wgt_0_520,Wgt_0_521,Wgt_0_522,Wgt_0_523,Wgt_0_524,Wgt_0_525,Wgt_0_526,Wgt_0_527,Wgt_0_528,Wgt_0_529,Wgt_0_530,Wgt_0_531,Wgt_0_532,Wgt_0_533,Wgt_0_534,Wgt_0_535,Wgt_0_536,Wgt_0_537,Wgt_0_538,Wgt_0_539,Wgt_0_540,Wgt_0_541,Wgt_0_542,Wgt_0_543,Wgt_0_544,Wgt_0_545,Wgt_0_546,Wgt_0_547,Wgt_0_548,Wgt_0_549,Wgt_0_550,Wgt_0_551,Wgt_0_552,Wgt_0_553,Wgt_0_554,Wgt_0_555,Wgt_0_556,Wgt_0_557,Wgt_0_558,Wgt_0_559,Wgt_0_560,Wgt_0_561,Wgt_0_562,Wgt_0_563,Wgt_0_564,Wgt_0_565,Wgt_0_566,Wgt_0_567,Wgt_0_568,Wgt_0_569,Wgt_0_570,Wgt_0_571,Wgt_0_572,Wgt_0_573,Wgt_0_574,Wgt_0_575,Wgt_0_576,Wgt_0_577,Wgt_0_578,Wgt_0_579,Wgt_0_580,Wgt_0_581,Wgt_0_582,Wgt_0_583,Wgt_0_584,Wgt_0_585,Wgt_0_586,Wgt_0_587,Wgt_0_588,Wgt_0_589,Wgt_0_590,Wgt_0_591,Wgt_0_592,Wgt_0_593,Wgt_0_594,Wgt_0_595,Wgt_0_596,Wgt_0_597,Wgt_0_598,Wgt_0_599,Wgt_0_600,Wgt_0_601,Wgt_0_602,Wgt_0_603,Wgt_0_604,Wgt_0_605,Wgt_0_606,Wgt_0_607,Wgt_0_608,Wgt_0_609,Wgt_0_610,Wgt_0_611,Wgt_0_612,Wgt_0_613,Wgt_0_614,Wgt_0_615,Wgt_0_616,Wgt_0_617,Wgt_0_618,Wgt_0_619,Wgt_0_620,Wgt_0_621,Wgt_0_622,Wgt_0_623,Wgt_0_624,Wgt_0_625,Wgt_0_626,Wgt_0_627,Wgt_0_628,Wgt_0_629,Wgt_0_630,Wgt_0_631,Wgt_0_632,Wgt_0_633,Wgt_0_634,Wgt_0_635,Wgt_0_636,Wgt_0_637,Wgt_0_638,Wgt_0_639,Wgt_0_640,Wgt_0_641,Wgt_0_642,Wgt_0_643,Wgt_0_644,Wgt_0_645,Wgt_0_646,Wgt_0_647,Wgt_0_648,Wgt_0_649,Wgt_0_650,Wgt_0_651,Wgt_0_652,Wgt_0_653,Wgt_0_654,Wgt_0_655,Wgt_0_656,Wgt_0_657,Wgt_0_658,Wgt_0_659,Wgt_0_660,Wgt_0_661,Wgt_0_662,Wgt_0_663,Wgt_0_664,Wgt_0_665,Wgt_0_666,Wgt_0_667,Wgt_0_668,Wgt_0_669,Wgt_0_670,Wgt_0_671,Wgt_0_672,Wgt_0_673,Wgt_0_674,Wgt_0_675,Wgt_0_676,Wgt_0_677,Wgt_0_678,Wgt_0_679,Wgt_0_680,Wgt_0_681,Wgt_0_682,Wgt_0_683,Wgt_0_684,Wgt_0_685,Wgt_0_686,Wgt_0_687,Wgt_0_688,Wgt_0_689,Wgt_0_690,Wgt_0_691,Wgt_0_692,Wgt_0_693,Wgt_0_694,Wgt_0_695,Wgt_0_696,Wgt_0_697,Wgt_0_698,Wgt_0_699,Wgt_0_700,Wgt_0_701,Wgt_0_702,Wgt_0_703,Wgt_0_704,Wgt_0_705,Wgt_0_706,Wgt_0_707,Wgt_0_708,Wgt_0_709,Wgt_0_710,Wgt_0_711,Wgt_0_712,Wgt_0_713,Wgt_0_714,Wgt_0_715,Wgt_0_716,Wgt_0_717,Wgt_0_718,Wgt_0_719,Wgt_0_720,Wgt_0_721,Wgt_0_722,Wgt_0_723,Wgt_0_724,Wgt_0_725,Wgt_0_726,Wgt_0_727,Wgt_0_728,Wgt_0_729,Wgt_0_730,Wgt_0_731,Wgt_0_732,Wgt_0_733,Wgt_0_734,Wgt_0_735,Wgt_0_736,Wgt_0_737,Wgt_0_738,Wgt_0_739,Wgt_0_740,Wgt_0_741,Wgt_0_742,Wgt_0_743,Wgt_0_744,Wgt_0_745,Wgt_0_746,Wgt_0_747,Wgt_0_748,Wgt_0_749,Wgt_0_750,Wgt_0_751,Wgt_0_752,Wgt_0_753,Wgt_0_754,Wgt_0_755,Wgt_0_756,Wgt_0_757,Wgt_0_758,Wgt_0_759,Wgt_0_760,Wgt_0_761,Wgt_0_762,Wgt_0_763,Wgt_0_764,Wgt_0_765,Wgt_0_766,Wgt_0_767,Wgt_0_768,Wgt_0_769,Wgt_0_770,Wgt_0_771,Wgt_0_772,Wgt_0_773,Wgt_0_774,Wgt_0_775,Wgt_0_776,Wgt_0_777,Wgt_0_778,Wgt_0_779,Wgt_0_780,Wgt_0_781,Wgt_0_782,Wgt_0_783,Wgt_0_784,Wgt_1_0,Wgt_1_1,Wgt_1_2,Wgt_1_3,Wgt_1_4,Wgt_1_5,Wgt_1_6,Wgt_1_7,Wgt_1_8,Wgt_1_9,Wgt_1_10,Wgt_1_11,Wgt_1_12,Wgt_1_13,Wgt_1_14,Wgt_1_15,Wgt_1_16,Wgt_1_17,Wgt_1_18,Wgt_1_19,Wgt_1_20,Wgt_1_21,Wgt_1_22,Wgt_1_23,Wgt_1_24,Wgt_1_25,Wgt_1_26,Wgt_1_27,Wgt_1_28,Wgt_1_29,Wgt_1_30,Wgt_1_31,Wgt_1_32,Wgt_1_33,Wgt_1_34,Wgt_1_35,Wgt_1_36,Wgt_1_37,Wgt_1_38,Wgt_1_39,Wgt_1_40,Wgt_1_41,Wgt_1_42,Wgt_1_43,Wgt_1_44,Wgt_1_45,Wgt_1_46,Wgt_1_47,Wgt_1_48,Wgt_1_49,Wgt_1_50,Wgt_1_51,Wgt_1_52,Wgt_1_53,Wgt_1_54,Wgt_1_55,Wgt_1_56,Wgt_1_57,Wgt_1_58,Wgt_1_59,Wgt_1_60,Wgt_1_61,Wgt_1_62,Wgt_1_63,Wgt_1_64,Wgt_1_65,Wgt_1_66,Wgt_1_67,Wgt_1_68,Wgt_1_69,Wgt_1_70,Wgt_1_71,Wgt_1_72,Wgt_1_73,Wgt_1_74,Wgt_1_75,Wgt_1_76,Wgt_1_77,Wgt_1_78,Wgt_1_79,Wgt_1_80,Wgt_1_81,Wgt_1_82,Wgt_1_83,Wgt_1_84,Wgt_1_85,Wgt_1_86,Wgt_1_87,Wgt_1_88,Wgt_1_89,Wgt_1_90,Wgt_1_91,Wgt_1_92,Wgt_1_93,Wgt_1_94,Wgt_1_95,Wgt_1_96,Wgt_1_97,Wgt_1_98,Wgt_1_99,Wgt_1_100,Wgt_1_101,Wgt_1_102,Wgt_1_103,Wgt_1_104,Wgt_1_105,Wgt_1_106,Wgt_1_107,Wgt_1_108,Wgt_1_109,Wgt_1_110,Wgt_1_111,Wgt_1_112,Wgt_1_113,Wgt_1_114,Wgt_1_115,Wgt_1_116,Wgt_1_117,Wgt_1_118,Wgt_1_119,Wgt_1_120,Wgt_1_121,Wgt_1_122,Wgt_1_123,Wgt_1_124,Wgt_1_125,Wgt_1_126,Wgt_1_127,Wgt_1_128,Wgt_1_129,Wgt_1_130,Wgt_1_131,Wgt_1_132,Wgt_1_133,Wgt_1_134,Wgt_1_135,Wgt_1_136,Wgt_1_137,Wgt_1_138,Wgt_1_139,Wgt_1_140,Wgt_1_141,Wgt_1_142,Wgt_1_143,Wgt_1_144,Wgt_1_145,Wgt_1_146,Wgt_1_147,Wgt_1_148,Wgt_1_149,Wgt_1_150,Wgt_1_151,Wgt_1_152,Wgt_1_153,Wgt_1_154,Wgt_1_155,Wgt_1_156,Wgt_1_157,Wgt_1_158,Wgt_1_159,Wgt_1_160,Wgt_1_161,Wgt_1_162,Wgt_1_163,Wgt_1_164,Wgt_1_165,Wgt_1_166,Wgt_1_167,Wgt_1_168,Wgt_1_169,Wgt_1_170,Wgt_1_171,Wgt_1_172,Wgt_1_173,Wgt_1_174,Wgt_1_175,Wgt_1_176,Wgt_1_177,Wgt_1_178,Wgt_1_179,Wgt_1_180,Wgt_1_181,Wgt_1_182,Wgt_1_183,Wgt_1_184,Wgt_1_185,Wgt_1_186,Wgt_1_187,Wgt_1_188,Wgt_1_189,Wgt_1_190,Wgt_1_191,Wgt_1_192,Wgt_1_193,Wgt_1_194,Wgt_1_195,Wgt_1_196,Wgt_1_197,Wgt_1_198,Wgt_1_199,Wgt_1_200,Wgt_1_201,Wgt_1_202,Wgt_1_203,Wgt_1_204,Wgt_1_205,Wgt_1_206,Wgt_1_207,Wgt_1_208,Wgt_1_209,Wgt_1_210,Wgt_1_211,Wgt_1_212,Wgt_1_213,Wgt_1_214,Wgt_1_215,Wgt_1_216,Wgt_1_217,Wgt_1_218,Wgt_1_219,Wgt_1_220,Wgt_1_221,Wgt_1_222,Wgt_1_223,Wgt_1_224,Wgt_1_225,Wgt_1_226,Wgt_1_227,Wgt_1_228,Wgt_1_229,Wgt_1_230,Wgt_1_231,Wgt_1_232,Wgt_1_233,Wgt_1_234,Wgt_1_235,Wgt_1_236,Wgt_1_237,Wgt_1_238,Wgt_1_239,Wgt_1_240,Wgt_1_241,Wgt_1_242,Wgt_1_243,Wgt_1_244,Wgt_1_245,Wgt_1_246,Wgt_1_247,Wgt_1_248,Wgt_1_249,Wgt_1_250,Wgt_1_251,Wgt_1_252,Wgt_1_253,Wgt_1_254,Wgt_1_255,Wgt_1_256,Wgt_1_257,Wgt_1_258,Wgt_1_259,Wgt_1_260,Wgt_1_261,Wgt_1_262,Wgt_1_263,Wgt_1_264,Wgt_1_265,Wgt_1_266,Wgt_1_267,Wgt_1_268,Wgt_1_269,Wgt_1_270,Wgt_1_271,Wgt_1_272,Wgt_1_273,Wgt_1_274,Wgt_1_275,Wgt_1_276,Wgt_1_277,Wgt_1_278,Wgt_1_279,Wgt_1_280,Wgt_1_281,Wgt_1_282,Wgt_1_283,Wgt_1_284,Wgt_1_285,Wgt_1_286,Wgt_1_287,Wgt_1_288,Wgt_1_289,Wgt_1_290,Wgt_1_291,Wgt_1_292,Wgt_1_293,Wgt_1_294,Wgt_1_295,Wgt_1_296,Wgt_1_297,Wgt_1_298,Wgt_1_299,Wgt_1_300,Wgt_1_301,Wgt_1_302,Wgt_1_303,Wgt_1_304,Wgt_1_305,Wgt_1_306,Wgt_1_307,Wgt_1_308,Wgt_1_309,Wgt_1_310,Wgt_1_311,Wgt_1_312,Wgt_1_313,Wgt_1_314,Wgt_1_315,Wgt_1_316,Wgt_1_317,Wgt_1_318,Wgt_1_319,Wgt_1_320,Wgt_1_321,Wgt_1_322,Wgt_1_323,Wgt_1_324,Wgt_1_325,Wgt_1_326,Wgt_1_327,Wgt_1_328,Wgt_1_329,Wgt_1_330,Wgt_1_331,Wgt_1_332,Wgt_1_333,Wgt_1_334,Wgt_1_335,Wgt_1_336,Wgt_1_337,Wgt_1_338,Wgt_1_339,Wgt_1_340,Wgt_1_341,Wgt_1_342,Wgt_1_343,Wgt_1_344,Wgt_1_345,Wgt_1_346,Wgt_1_347,Wgt_1_348,Wgt_1_349,Wgt_1_350,Wgt_1_351,Wgt_1_352,Wgt_1_353,Wgt_1_354,Wgt_1_355,Wgt_1_356,Wgt_1_357,Wgt_1_358,Wgt_1_359,Wgt_1_360,Wgt_1_361,Wgt_1_362,Wgt_1_363,Wgt_1_364,Wgt_1_365,Wgt_1_366,Wgt_1_367,Wgt_1_368,Wgt_1_369,Wgt_1_370,Wgt_1_371,Wgt_1_372,Wgt_1_373,Wgt_1_374,Wgt_1_375,Wgt_1_376,Wgt_1_377,Wgt_1_378,Wgt_1_379,Wgt_1_380,Wgt_1_381,Wgt_1_382,Wgt_1_383,Wgt_1_384,Wgt_1_385,Wgt_1_386,Wgt_1_387,Wgt_1_388,Wgt_1_389,Wgt_1_390,Wgt_1_391,Wgt_1_392,Wgt_1_393,Wgt_1_394,Wgt_1_395,Wgt_1_396,Wgt_1_397,Wgt_1_398,Wgt_1_399,Wgt_1_400,Wgt_1_401,Wgt_1_402,Wgt_1_403,Wgt_1_404,Wgt_1_405,Wgt_1_406,Wgt_1_407,Wgt_1_408,Wgt_1_409,Wgt_1_410,Wgt_1_411,Wgt_1_412,Wgt_1_413,Wgt_1_414,Wgt_1_415,Wgt_1_416,Wgt_1_417,Wgt_1_418,Wgt_1_419,Wgt_1_420,Wgt_1_421,Wgt_1_422,Wgt_1_423,Wgt_1_424,Wgt_1_425,Wgt_1_426,Wgt_1_427,Wgt_1_428,Wgt_1_429,Wgt_1_430,Wgt_1_431,Wgt_1_432,Wgt_1_433,Wgt_1_434,Wgt_1_435,Wgt_1_436,Wgt_1_437,Wgt_1_438,Wgt_1_439,Wgt_1_440,Wgt_1_441,Wgt_1_442,Wgt_1_443,Wgt_1_444,Wgt_1_445,Wgt_1_446,Wgt_1_447,Wgt_1_448,Wgt_1_449,Wgt_1_450,Wgt_1_451,Wgt_1_452,Wgt_1_453,Wgt_1_454,Wgt_1_455,Wgt_1_456,Wgt_1_457,Wgt_1_458,Wgt_1_459,Wgt_1_460,Wgt_1_461,Wgt_1_462,Wgt_1_463,Wgt_1_464,Wgt_1_465,Wgt_1_466,Wgt_1_467,Wgt_1_468,Wgt_1_469,Wgt_1_470,Wgt_1_471,Wgt_1_472,Wgt_1_473,Wgt_1_474,Wgt_1_475,Wgt_1_476,Wgt_1_477,Wgt_1_478,Wgt_1_479,Wgt_1_480,Wgt_1_481,Wgt_1_482,Wgt_1_483,Wgt_1_484,Wgt_1_485,Wgt_1_486,Wgt_1_487,Wgt_1_488,Wgt_1_489,Wgt_1_490,Wgt_1_491,Wgt_1_492,Wgt_1_493,Wgt_1_494,Wgt_1_495,Wgt_1_496,Wgt_1_497,Wgt_1_498,Wgt_1_499,Wgt_1_500,Wgt_1_501,Wgt_1_502,Wgt_1_503,Wgt_1_504,Wgt_1_505,Wgt_1_506,Wgt_1_507,Wgt_1_508,Wgt_1_509,Wgt_1_510,Wgt_1_511,Wgt_1_512,Wgt_1_513,Wgt_1_514,Wgt_1_515,Wgt_1_516,Wgt_1_517,Wgt_1_518,Wgt_1_519,Wgt_1_520,Wgt_1_521,Wgt_1_522,Wgt_1_523,Wgt_1_524,Wgt_1_525,Wgt_1_526,Wgt_1_527,Wgt_1_528,Wgt_1_529,Wgt_1_530,Wgt_1_531,Wgt_1_532,Wgt_1_533,Wgt_1_534,Wgt_1_535,Wgt_1_536,Wgt_1_537,Wgt_1_538,Wgt_1_539,Wgt_1_540,Wgt_1_541,Wgt_1_542,Wgt_1_543,Wgt_1_544,Wgt_1_545,Wgt_1_546,Wgt_1_547,Wgt_1_548,Wgt_1_549,Wgt_1_550,Wgt_1_551,Wgt_1_552,Wgt_1_553,Wgt_1_554,Wgt_1_555,Wgt_1_556,Wgt_1_557,Wgt_1_558,Wgt_1_559,Wgt_1_560,Wgt_1_561,Wgt_1_562,Wgt_1_563,Wgt_1_564,Wgt_1_565,Wgt_1_566,Wgt_1_567,Wgt_1_568,Wgt_1_569,Wgt_1_570,Wgt_1_571,Wgt_1_572,Wgt_1_573,Wgt_1_574,Wgt_1_575,Wgt_1_576,Wgt_1_577,Wgt_1_578,Wgt_1_579,Wgt_1_580,Wgt_1_581,Wgt_1_582,Wgt_1_583,Wgt_1_584,Wgt_1_585,Wgt_1_586,Wgt_1_587,Wgt_1_588,Wgt_1_589,Wgt_1_590,Wgt_1_591,Wgt_1_592,Wgt_1_593,Wgt_1_594,Wgt_1_595,Wgt_1_596,Wgt_1_597,Wgt_1_598,Wgt_1_599,Wgt_1_600,Wgt_1_601,Wgt_1_602,Wgt_1_603,Wgt_1_604,Wgt_1_605,Wgt_1_606,Wgt_1_607,Wgt_1_608,Wgt_1_609,Wgt_1_610,Wgt_1_611,Wgt_1_612,Wgt_1_613,Wgt_1_614,Wgt_1_615,Wgt_1_616,Wgt_1_617,Wgt_1_618,Wgt_1_619,Wgt_1_620,Wgt_1_621,Wgt_1_622,Wgt_1_623,Wgt_1_624,Wgt_1_625,Wgt_1_626,Wgt_1_627,Wgt_1_628,Wgt_1_629,Wgt_1_630,Wgt_1_631,Wgt_1_632,Wgt_1_633,Wgt_1_634,Wgt_1_635,Wgt_1_636,Wgt_1_637,Wgt_1_638,Wgt_1_639,Wgt_1_640,Wgt_1_641,Wgt_1_642,Wgt_1_643,Wgt_1_644,Wgt_1_645,Wgt_1_646,Wgt_1_647,Wgt_1_648,Wgt_1_649,Wgt_1_650,Wgt_1_651,Wgt_1_652,Wgt_1_653,Wgt_1_654,Wgt_1_655,Wgt_1_656,Wgt_1_657,Wgt_1_658,Wgt_1_659,Wgt_1_660,Wgt_1_661,Wgt_1_662,Wgt_1_663,Wgt_1_664,Wgt_1_665,Wgt_1_666,Wgt_1_667,Wgt_1_668,Wgt_1_669,Wgt_1_670,Wgt_1_671,Wgt_1_672,Wgt_1_673,Wgt_1_674,Wgt_1_675,Wgt_1_676,Wgt_1_677,Wgt_1_678,Wgt_1_679,Wgt_1_680,Wgt_1_681,Wgt_1_682,Wgt_1_683,Wgt_1_684,Wgt_1_685,Wgt_1_686,Wgt_1_687,Wgt_1_688,Wgt_1_689,Wgt_1_690,Wgt_1_691,Wgt_1_692,Wgt_1_693,Wgt_1_694,Wgt_1_695,Wgt_1_696,Wgt_1_697,Wgt_1_698,Wgt_1_699,Wgt_1_700,Wgt_1_701,Wgt_1_702,Wgt_1_703,Wgt_1_704,Wgt_1_705,Wgt_1_706,Wgt_1_707,Wgt_1_708,Wgt_1_709,Wgt_1_710,Wgt_1_711,Wgt_1_712,Wgt_1_713,Wgt_1_714,Wgt_1_715,Wgt_1_716,Wgt_1_717,Wgt_1_718,Wgt_1_719,Wgt_1_720,Wgt_1_721,Wgt_1_722,Wgt_1_723,Wgt_1_724,Wgt_1_725,Wgt_1_726,Wgt_1_727,Wgt_1_728,Wgt_1_729,Wgt_1_730,Wgt_1_731,Wgt_1_732,Wgt_1_733,Wgt_1_734,Wgt_1_735,Wgt_1_736,Wgt_1_737,Wgt_1_738,Wgt_1_739,Wgt_1_740,Wgt_1_741,Wgt_1_742,Wgt_1_743,Wgt_1_744,Wgt_1_745,Wgt_1_746,Wgt_1_747,Wgt_1_748,Wgt_1_749,Wgt_1_750,Wgt_1_751,Wgt_1_752,Wgt_1_753,Wgt_1_754,Wgt_1_755,Wgt_1_756,Wgt_1_757,Wgt_1_758,Wgt_1_759,Wgt_1_760,Wgt_1_761,Wgt_1_762,Wgt_1_763,Wgt_1_764,Wgt_1_765,Wgt_1_766,Wgt_1_767,Wgt_1_768,Wgt_1_769,Wgt_1_770,Wgt_1_771,Wgt_1_772,Wgt_1_773,Wgt_1_774,Wgt_1_775,Wgt_1_776,Wgt_1_777,Wgt_1_778,Wgt_1_779,Wgt_1_780,Wgt_1_781,Wgt_1_782,Wgt_1_783,Wgt_1_784,Wgt_2_0,Wgt_2_1,Wgt_2_2,Wgt_2_3,Wgt_2_4,Wgt_2_5,Wgt_2_6,Wgt_2_7,Wgt_2_8,Wgt_2_9,Wgt_2_10,Wgt_2_11,Wgt_2_12,Wgt_2_13,Wgt_2_14,Wgt_2_15,Wgt_2_16,Wgt_2_17,Wgt_2_18,Wgt_2_19,Wgt_2_20,Wgt_2_21,Wgt_2_22,Wgt_2_23,Wgt_2_24,Wgt_2_25,Wgt_2_26,Wgt_2_27,Wgt_2_28,Wgt_2_29,Wgt_2_30,Wgt_2_31,Wgt_2_32,Wgt_2_33,Wgt_2_34,Wgt_2_35,Wgt_2_36,Wgt_2_37,Wgt_2_38,Wgt_2_39,Wgt_2_40,Wgt_2_41,Wgt_2_42,Wgt_2_43,Wgt_2_44,Wgt_2_45,Wgt_2_46,Wgt_2_47,Wgt_2_48,Wgt_2_49,Wgt_2_50,Wgt_2_51,Wgt_2_52,Wgt_2_53,Wgt_2_54,Wgt_2_55,Wgt_2_56,Wgt_2_57,Wgt_2_58,Wgt_2_59,Wgt_2_60,Wgt_2_61,Wgt_2_62,Wgt_2_63,Wgt_2_64,Wgt_2_65,Wgt_2_66,Wgt_2_67,Wgt_2_68,Wgt_2_69,Wgt_2_70,Wgt_2_71,Wgt_2_72,Wgt_2_73,Wgt_2_74,Wgt_2_75,Wgt_2_76,Wgt_2_77,Wgt_2_78,Wgt_2_79,Wgt_2_80,Wgt_2_81,Wgt_2_82,Wgt_2_83,Wgt_2_84,Wgt_2_85,Wgt_2_86,Wgt_2_87,Wgt_2_88,Wgt_2_89,Wgt_2_90,Wgt_2_91,Wgt_2_92,Wgt_2_93,Wgt_2_94,Wgt_2_95,Wgt_2_96,Wgt_2_97,Wgt_2_98,Wgt_2_99,Wgt_2_100,Wgt_2_101,Wgt_2_102,Wgt_2_103,Wgt_2_104,Wgt_2_105,Wgt_2_106,Wgt_2_107,Wgt_2_108,Wgt_2_109,Wgt_2_110,Wgt_2_111,Wgt_2_112,Wgt_2_113,Wgt_2_114,Wgt_2_115,Wgt_2_116,Wgt_2_117,Wgt_2_118,Wgt_2_119,Wgt_2_120,Wgt_2_121,Wgt_2_122,Wgt_2_123,Wgt_2_124,Wgt_2_125,Wgt_2_126,Wgt_2_127,Wgt_2_128,Wgt_2_129,Wgt_2_130,Wgt_2_131,Wgt_2_132,Wgt_2_133,Wgt_2_134,Wgt_2_135,Wgt_2_136,Wgt_2_137,Wgt_2_138,Wgt_2_139,Wgt_2_140,Wgt_2_141,Wgt_2_142,Wgt_2_143,Wgt_2_144,Wgt_2_145,Wgt_2_146,Wgt_2_147,Wgt_2_148,Wgt_2_149,Wgt_2_150,Wgt_2_151,Wgt_2_152,Wgt_2_153,Wgt_2_154,Wgt_2_155,Wgt_2_156,Wgt_2_157,Wgt_2_158,Wgt_2_159,Wgt_2_160,Wgt_2_161,Wgt_2_162,Wgt_2_163,Wgt_2_164,Wgt_2_165,Wgt_2_166,Wgt_2_167,Wgt_2_168,Wgt_2_169,Wgt_2_170,Wgt_2_171,Wgt_2_172,Wgt_2_173,Wgt_2_174,Wgt_2_175,Wgt_2_176,Wgt_2_177,Wgt_2_178,Wgt_2_179,Wgt_2_180,Wgt_2_181,Wgt_2_182,Wgt_2_183,Wgt_2_184,Wgt_2_185,Wgt_2_186,Wgt_2_187,Wgt_2_188,Wgt_2_189,Wgt_2_190,Wgt_2_191,Wgt_2_192,Wgt_2_193,Wgt_2_194,Wgt_2_195,Wgt_2_196,Wgt_2_197,Wgt_2_198,Wgt_2_199,Wgt_2_200,Wgt_2_201,Wgt_2_202,Wgt_2_203,Wgt_2_204,Wgt_2_205,Wgt_2_206,Wgt_2_207,Wgt_2_208,Wgt_2_209,Wgt_2_210,Wgt_2_211,Wgt_2_212,Wgt_2_213,Wgt_2_214,Wgt_2_215,Wgt_2_216,Wgt_2_217,Wgt_2_218,Wgt_2_219,Wgt_2_220,Wgt_2_221,Wgt_2_222,Wgt_2_223,Wgt_2_224,Wgt_2_225,Wgt_2_226,Wgt_2_227,Wgt_2_228,Wgt_2_229,Wgt_2_230,Wgt_2_231,Wgt_2_232,Wgt_2_233,Wgt_2_234,Wgt_2_235,Wgt_2_236,Wgt_2_237,Wgt_2_238,Wgt_2_239,Wgt_2_240,Wgt_2_241,Wgt_2_242,Wgt_2_243,Wgt_2_244,Wgt_2_245,Wgt_2_246,Wgt_2_247,Wgt_2_248,Wgt_2_249,Wgt_2_250,Wgt_2_251,Wgt_2_252,Wgt_2_253,Wgt_2_254,Wgt_2_255,Wgt_2_256,Wgt_2_257,Wgt_2_258,Wgt_2_259,Wgt_2_260,Wgt_2_261,Wgt_2_262,Wgt_2_263,Wgt_2_264,Wgt_2_265,Wgt_2_266,Wgt_2_267,Wgt_2_268,Wgt_2_269,Wgt_2_270,Wgt_2_271,Wgt_2_272,Wgt_2_273,Wgt_2_274,Wgt_2_275,Wgt_2_276,Wgt_2_277,Wgt_2_278,Wgt_2_279,Wgt_2_280,Wgt_2_281,Wgt_2_282,Wgt_2_283,Wgt_2_284,Wgt_2_285,Wgt_2_286,Wgt_2_287,Wgt_2_288,Wgt_2_289,Wgt_2_290,Wgt_2_291,Wgt_2_292,Wgt_2_293,Wgt_2_294,Wgt_2_295,Wgt_2_296,Wgt_2_297,Wgt_2_298,Wgt_2_299,Wgt_2_300,Wgt_2_301,Wgt_2_302,Wgt_2_303,Wgt_2_304,Wgt_2_305,Wgt_2_306,Wgt_2_307,Wgt_2_308,Wgt_2_309,Wgt_2_310,Wgt_2_311,Wgt_2_312,Wgt_2_313,Wgt_2_314,Wgt_2_315,Wgt_2_316,Wgt_2_317,Wgt_2_318,Wgt_2_319,Wgt_2_320,Wgt_2_321,Wgt_2_322,Wgt_2_323,Wgt_2_324,Wgt_2_325,Wgt_2_326,Wgt_2_327,Wgt_2_328,Wgt_2_329,Wgt_2_330,Wgt_2_331,Wgt_2_332,Wgt_2_333,Wgt_2_334,Wgt_2_335,Wgt_2_336,Wgt_2_337,Wgt_2_338,Wgt_2_339,Wgt_2_340,Wgt_2_341,Wgt_2_342,Wgt_2_343,Wgt_2_344,Wgt_2_345,Wgt_2_346,Wgt_2_347,Wgt_2_348,Wgt_2_349,Wgt_2_350,Wgt_2_351,Wgt_2_352,Wgt_2_353,Wgt_2_354,Wgt_2_355,Wgt_2_356,Wgt_2_357,Wgt_2_358,Wgt_2_359,Wgt_2_360,Wgt_2_361,Wgt_2_362,Wgt_2_363,Wgt_2_364,Wgt_2_365,Wgt_2_366,Wgt_2_367,Wgt_2_368,Wgt_2_369,Wgt_2_370,Wgt_2_371,Wgt_2_372,Wgt_2_373,Wgt_2_374,Wgt_2_375,Wgt_2_376,Wgt_2_377,Wgt_2_378,Wgt_2_379,Wgt_2_380,Wgt_2_381,Wgt_2_382,Wgt_2_383,Wgt_2_384,Wgt_2_385,Wgt_2_386,Wgt_2_387,Wgt_2_388,Wgt_2_389,Wgt_2_390,Wgt_2_391,Wgt_2_392,Wgt_2_393,Wgt_2_394,Wgt_2_395,Wgt_2_396,Wgt_2_397,Wgt_2_398,Wgt_2_399,Wgt_2_400,Wgt_2_401,Wgt_2_402,Wgt_2_403,Wgt_2_404,Wgt_2_405,Wgt_2_406,Wgt_2_407,Wgt_2_408,Wgt_2_409,Wgt_2_410,Wgt_2_411,Wgt_2_412,Wgt_2_413,Wgt_2_414,Wgt_2_415,Wgt_2_416,Wgt_2_417,Wgt_2_418,Wgt_2_419,Wgt_2_420,Wgt_2_421,Wgt_2_422,Wgt_2_423,Wgt_2_424,Wgt_2_425,Wgt_2_426,Wgt_2_427,Wgt_2_428,Wgt_2_429,Wgt_2_430,Wgt_2_431,Wgt_2_432,Wgt_2_433,Wgt_2_434,Wgt_2_435,Wgt_2_436,Wgt_2_437,Wgt_2_438,Wgt_2_439,Wgt_2_440,Wgt_2_441,Wgt_2_442,Wgt_2_443,Wgt_2_444,Wgt_2_445,Wgt_2_446,Wgt_2_447,Wgt_2_448,Wgt_2_449,Wgt_2_450,Wgt_2_451,Wgt_2_452,Wgt_2_453,Wgt_2_454,Wgt_2_455,Wgt_2_456,Wgt_2_457,Wgt_2_458,Wgt_2_459,Wgt_2_460,Wgt_2_461,Wgt_2_462,Wgt_2_463,Wgt_2_464,Wgt_2_465,Wgt_2_466,Wgt_2_467,Wgt_2_468,Wgt_2_469,Wgt_2_470,Wgt_2_471,Wgt_2_472,Wgt_2_473,Wgt_2_474,Wgt_2_475,Wgt_2_476,Wgt_2_477,Wgt_2_478,Wgt_2_479,Wgt_2_480,Wgt_2_481,Wgt_2_482,Wgt_2_483,Wgt_2_484,Wgt_2_485,Wgt_2_486,Wgt_2_487,Wgt_2_488,Wgt_2_489,Wgt_2_490,Wgt_2_491,Wgt_2_492,Wgt_2_493,Wgt_2_494,Wgt_2_495,Wgt_2_496,Wgt_2_497,Wgt_2_498,Wgt_2_499,Wgt_2_500,Wgt_2_501,Wgt_2_502,Wgt_2_503,Wgt_2_504,Wgt_2_505,Wgt_2_506,Wgt_2_507,Wgt_2_508,Wgt_2_509,Wgt_2_510,Wgt_2_511,Wgt_2_512,Wgt_2_513,Wgt_2_514,Wgt_2_515,Wgt_2_516,Wgt_2_517,Wgt_2_518,Wgt_2_519,Wgt_2_520,Wgt_2_521,Wgt_2_522,Wgt_2_523,Wgt_2_524,Wgt_2_525,Wgt_2_526,Wgt_2_527,Wgt_2_528,Wgt_2_529,Wgt_2_530,Wgt_2_531,Wgt_2_532,Wgt_2_533,Wgt_2_534,Wgt_2_535,Wgt_2_536,Wgt_2_537,Wgt_2_538,Wgt_2_539,Wgt_2_540,Wgt_2_541,Wgt_2_542,Wgt_2_543,Wgt_2_544,Wgt_2_545,Wgt_2_546,Wgt_2_547,Wgt_2_548,Wgt_2_549,Wgt_2_550,Wgt_2_551,Wgt_2_552,Wgt_2_553,Wgt_2_554,Wgt_2_555,Wgt_2_556,Wgt_2_557,Wgt_2_558,Wgt_2_559,Wgt_2_560,Wgt_2_561,Wgt_2_562,Wgt_2_563,Wgt_2_564,Wgt_2_565,Wgt_2_566,Wgt_2_567,Wgt_2_568,Wgt_2_569,Wgt_2_570,Wgt_2_571,Wgt_2_572,Wgt_2_573,Wgt_2_574,Wgt_2_575,Wgt_2_576,Wgt_2_577,Wgt_2_578,Wgt_2_579,Wgt_2_580,Wgt_2_581,Wgt_2_582,Wgt_2_583,Wgt_2_584,Wgt_2_585,Wgt_2_586,Wgt_2_587,Wgt_2_588,Wgt_2_589,Wgt_2_590,Wgt_2_591,Wgt_2_592,Wgt_2_593,Wgt_2_594,Wgt_2_595,Wgt_2_596,Wgt_2_597,Wgt_2_598,Wgt_2_599,Wgt_2_600,Wgt_2_601,Wgt_2_602,Wgt_2_603,Wgt_2_604,Wgt_2_605,Wgt_2_606,Wgt_2_607,Wgt_2_608,Wgt_2_609,Wgt_2_610,Wgt_2_611,Wgt_2_612,Wgt_2_613,Wgt_2_614,Wgt_2_615,Wgt_2_616,Wgt_2_617,Wgt_2_618,Wgt_2_619,Wgt_2_620,Wgt_2_621,Wgt_2_622,Wgt_2_623,Wgt_2_624,Wgt_2_625,Wgt_2_626,Wgt_2_627,Wgt_2_628,Wgt_2_629,Wgt_2_630,Wgt_2_631,Wgt_2_632,Wgt_2_633,Wgt_2_634,Wgt_2_635,Wgt_2_636,Wgt_2_637,Wgt_2_638,Wgt_2_639,Wgt_2_640,Wgt_2_641,Wgt_2_642,Wgt_2_643,Wgt_2_644,Wgt_2_645,Wgt_2_646,Wgt_2_647,Wgt_2_648,Wgt_2_649,Wgt_2_650,Wgt_2_651,Wgt_2_652,Wgt_2_653,Wgt_2_654,Wgt_2_655,Wgt_2_656,Wgt_2_657,Wgt_2_658,Wgt_2_659,Wgt_2_660,Wgt_2_661,Wgt_2_662,Wgt_2_663,Wgt_2_664,Wgt_2_665,Wgt_2_666,Wgt_2_667,Wgt_2_668,Wgt_2_669,Wgt_2_670,Wgt_2_671,Wgt_2_672,Wgt_2_673,Wgt_2_674,Wgt_2_675,Wgt_2_676,Wgt_2_677,Wgt_2_678,Wgt_2_679,Wgt_2_680,Wgt_2_681,Wgt_2_682,Wgt_2_683,Wgt_2_684,Wgt_2_685,Wgt_2_686,Wgt_2_687,Wgt_2_688,Wgt_2_689,Wgt_2_690,Wgt_2_691,Wgt_2_692,Wgt_2_693,Wgt_2_694,Wgt_2_695,Wgt_2_696,Wgt_2_697,Wgt_2_698,Wgt_2_699,Wgt_2_700,Wgt_2_701,Wgt_2_702,Wgt_2_703,Wgt_2_704,Wgt_2_705,Wgt_2_706,Wgt_2_707,Wgt_2_708,Wgt_2_709,Wgt_2_710,Wgt_2_711,Wgt_2_712,Wgt_2_713,Wgt_2_714,Wgt_2_715,Wgt_2_716,Wgt_2_717,Wgt_2_718,Wgt_2_719,Wgt_2_720,Wgt_2_721,Wgt_2_722,Wgt_2_723,Wgt_2_724,Wgt_2_725,Wgt_2_726,Wgt_2_727,Wgt_2_728,Wgt_2_729,Wgt_2_730,Wgt_2_731,Wgt_2_732,Wgt_2_733,Wgt_2_734,Wgt_2_735,Wgt_2_736,Wgt_2_737,Wgt_2_738,Wgt_2_739,Wgt_2_740,Wgt_2_741,Wgt_2_742,Wgt_2_743,Wgt_2_744,Wgt_2_745,Wgt_2_746,Wgt_2_747,Wgt_2_748,Wgt_2_749,Wgt_2_750,Wgt_2_751,Wgt_2_752,Wgt_2_753,Wgt_2_754,Wgt_2_755,Wgt_2_756,Wgt_2_757,Wgt_2_758,Wgt_2_759,Wgt_2_760,Wgt_2_761,Wgt_2_762,Wgt_2_763,Wgt_2_764,Wgt_2_765,Wgt_2_766,Wgt_2_767,Wgt_2_768,Wgt_2_769,Wgt_2_770,Wgt_2_771,Wgt_2_772,Wgt_2_773,Wgt_2_774,Wgt_2_775,Wgt_2_776,Wgt_2_777,Wgt_2_778,Wgt_2_779,Wgt_2_780,Wgt_2_781,Wgt_2_782,Wgt_2_783,Wgt_2_784,Wgt_3_0,Wgt_3_1,Wgt_3_2,Wgt_3_3,Wgt_3_4,Wgt_3_5,Wgt_3_6,Wgt_3_7,Wgt_3_8,Wgt_3_9,Wgt_3_10,Wgt_3_11,Wgt_3_12,Wgt_3_13,Wgt_3_14,Wgt_3_15,Wgt_3_16,Wgt_3_17,Wgt_3_18,Wgt_3_19,Wgt_3_20,Wgt_3_21,Wgt_3_22,Wgt_3_23,Wgt_3_24,Wgt_3_25,Wgt_3_26,Wgt_3_27,Wgt_3_28,Wgt_3_29,Wgt_3_30,Wgt_3_31,Wgt_3_32,Wgt_3_33,Wgt_3_34,Wgt_3_35,Wgt_3_36,Wgt_3_37,Wgt_3_38,Wgt_3_39,Wgt_3_40,Wgt_3_41,Wgt_3_42,Wgt_3_43,Wgt_3_44,Wgt_3_45,Wgt_3_46,Wgt_3_47,Wgt_3_48,Wgt_3_49,Wgt_3_50,Wgt_3_51,Wgt_3_52,Wgt_3_53,Wgt_3_54,Wgt_3_55,Wgt_3_56,Wgt_3_57,Wgt_3_58,Wgt_3_59,Wgt_3_60,Wgt_3_61,Wgt_3_62,Wgt_3_63,Wgt_3_64,Wgt_3_65,Wgt_3_66,Wgt_3_67,Wgt_3_68,Wgt_3_69,Wgt_3_70,Wgt_3_71,Wgt_3_72,Wgt_3_73,Wgt_3_74,Wgt_3_75,Wgt_3_76,Wgt_3_77,Wgt_3_78,Wgt_3_79,Wgt_3_80,Wgt_3_81,Wgt_3_82,Wgt_3_83,Wgt_3_84,Wgt_3_85,Wgt_3_86,Wgt_3_87,Wgt_3_88,Wgt_3_89,Wgt_3_90,Wgt_3_91,Wgt_3_92,Wgt_3_93,Wgt_3_94,Wgt_3_95,Wgt_3_96,Wgt_3_97,Wgt_3_98,Wgt_3_99,Wgt_3_100,Wgt_3_101,Wgt_3_102,Wgt_3_103,Wgt_3_104,Wgt_3_105,Wgt_3_106,Wgt_3_107,Wgt_3_108,Wgt_3_109,Wgt_3_110,Wgt_3_111,Wgt_3_112,Wgt_3_113,Wgt_3_114,Wgt_3_115,Wgt_3_116,Wgt_3_117,Wgt_3_118,Wgt_3_119,Wgt_3_120,Wgt_3_121,Wgt_3_122,Wgt_3_123,Wgt_3_124,Wgt_3_125,Wgt_3_126,Wgt_3_127,Wgt_3_128,Wgt_3_129,Wgt_3_130,Wgt_3_131,Wgt_3_132,Wgt_3_133,Wgt_3_134,Wgt_3_135,Wgt_3_136,Wgt_3_137,Wgt_3_138,Wgt_3_139,Wgt_3_140,Wgt_3_141,Wgt_3_142,Wgt_3_143,Wgt_3_144,Wgt_3_145,Wgt_3_146,Wgt_3_147,Wgt_3_148,Wgt_3_149,Wgt_3_150,Wgt_3_151,Wgt_3_152,Wgt_3_153,Wgt_3_154,Wgt_3_155,Wgt_3_156,Wgt_3_157,Wgt_3_158,Wgt_3_159,Wgt_3_160,Wgt_3_161,Wgt_3_162,Wgt_3_163,Wgt_3_164,Wgt_3_165,Wgt_3_166,Wgt_3_167,Wgt_3_168,Wgt_3_169,Wgt_3_170,Wgt_3_171,Wgt_3_172,Wgt_3_173,Wgt_3_174,Wgt_3_175,Wgt_3_176,Wgt_3_177,Wgt_3_178,Wgt_3_179,Wgt_3_180,Wgt_3_181,Wgt_3_182,Wgt_3_183,Wgt_3_184,Wgt_3_185,Wgt_3_186,Wgt_3_187,Wgt_3_188,Wgt_3_189,Wgt_3_190,Wgt_3_191,Wgt_3_192,Wgt_3_193,Wgt_3_194,Wgt_3_195,Wgt_3_196,Wgt_3_197,Wgt_3_198,Wgt_3_199,Wgt_3_200,Wgt_3_201,Wgt_3_202,Wgt_3_203,Wgt_3_204,Wgt_3_205,Wgt_3_206,Wgt_3_207,Wgt_3_208,Wgt_3_209,Wgt_3_210,Wgt_3_211,Wgt_3_212,Wgt_3_213,Wgt_3_214,Wgt_3_215,Wgt_3_216,Wgt_3_217,Wgt_3_218,Wgt_3_219,Wgt_3_220,Wgt_3_221,Wgt_3_222,Wgt_3_223,Wgt_3_224,Wgt_3_225,Wgt_3_226,Wgt_3_227,Wgt_3_228,Wgt_3_229,Wgt_3_230,Wgt_3_231,Wgt_3_232,Wgt_3_233,Wgt_3_234,Wgt_3_235,Wgt_3_236,Wgt_3_237,Wgt_3_238,Wgt_3_239,Wgt_3_240,Wgt_3_241,Wgt_3_242,Wgt_3_243,Wgt_3_244,Wgt_3_245,Wgt_3_246,Wgt_3_247,Wgt_3_248,Wgt_3_249,Wgt_3_250,Wgt_3_251,Wgt_3_252,Wgt_3_253,Wgt_3_254,Wgt_3_255,Wgt_3_256,Wgt_3_257,Wgt_3_258,Wgt_3_259,Wgt_3_260,Wgt_3_261,Wgt_3_262,Wgt_3_263,Wgt_3_264,Wgt_3_265,Wgt_3_266,Wgt_3_267,Wgt_3_268,Wgt_3_269,Wgt_3_270,Wgt_3_271,Wgt_3_272,Wgt_3_273,Wgt_3_274,Wgt_3_275,Wgt_3_276,Wgt_3_277,Wgt_3_278,Wgt_3_279,Wgt_3_280,Wgt_3_281,Wgt_3_282,Wgt_3_283,Wgt_3_284,Wgt_3_285,Wgt_3_286,Wgt_3_287,Wgt_3_288,Wgt_3_289,Wgt_3_290,Wgt_3_291,Wgt_3_292,Wgt_3_293,Wgt_3_294,Wgt_3_295,Wgt_3_296,Wgt_3_297,Wgt_3_298,Wgt_3_299,Wgt_3_300,Wgt_3_301,Wgt_3_302,Wgt_3_303,Wgt_3_304,Wgt_3_305,Wgt_3_306,Wgt_3_307,Wgt_3_308,Wgt_3_309,Wgt_3_310,Wgt_3_311,Wgt_3_312,Wgt_3_313,Wgt_3_314,Wgt_3_315,Wgt_3_316,Wgt_3_317,Wgt_3_318,Wgt_3_319,Wgt_3_320,Wgt_3_321,Wgt_3_322,Wgt_3_323,Wgt_3_324,Wgt_3_325,Wgt_3_326,Wgt_3_327,Wgt_3_328,Wgt_3_329,Wgt_3_330,Wgt_3_331,Wgt_3_332,Wgt_3_333,Wgt_3_334,Wgt_3_335,Wgt_3_336,Wgt_3_337,Wgt_3_338,Wgt_3_339,Wgt_3_340,Wgt_3_341,Wgt_3_342,Wgt_3_343,Wgt_3_344,Wgt_3_345,Wgt_3_346,Wgt_3_347,Wgt_3_348,Wgt_3_349,Wgt_3_350,Wgt_3_351,Wgt_3_352,Wgt_3_353,Wgt_3_354,Wgt_3_355,Wgt_3_356,Wgt_3_357,Wgt_3_358,Wgt_3_359,Wgt_3_360,Wgt_3_361,Wgt_3_362,Wgt_3_363,Wgt_3_364,Wgt_3_365,Wgt_3_366,Wgt_3_367,Wgt_3_368,Wgt_3_369,Wgt_3_370,Wgt_3_371,Wgt_3_372,Wgt_3_373,Wgt_3_374,Wgt_3_375,Wgt_3_376,Wgt_3_377,Wgt_3_378,Wgt_3_379,Wgt_3_380,Wgt_3_381,Wgt_3_382,Wgt_3_383,Wgt_3_384,Wgt_3_385,Wgt_3_386,Wgt_3_387,Wgt_3_388,Wgt_3_389,Wgt_3_390,Wgt_3_391,Wgt_3_392,Wgt_3_393,Wgt_3_394,Wgt_3_395,Wgt_3_396,Wgt_3_397,Wgt_3_398,Wgt_3_399,Wgt_3_400,Wgt_3_401,Wgt_3_402,Wgt_3_403,Wgt_3_404,Wgt_3_405,Wgt_3_406,Wgt_3_407,Wgt_3_408,Wgt_3_409,Wgt_3_410,Wgt_3_411,Wgt_3_412,Wgt_3_413,Wgt_3_414,Wgt_3_415,Wgt_3_416,Wgt_3_417,Wgt_3_418,Wgt_3_419,Wgt_3_420,Wgt_3_421,Wgt_3_422,Wgt_3_423,Wgt_3_424,Wgt_3_425,Wgt_3_426,Wgt_3_427,Wgt_3_428,Wgt_3_429,Wgt_3_430,Wgt_3_431,Wgt_3_432,Wgt_3_433,Wgt_3_434,Wgt_3_435,Wgt_3_436,Wgt_3_437,Wgt_3_438,Wgt_3_439,Wgt_3_440,Wgt_3_441,Wgt_3_442,Wgt_3_443,Wgt_3_444,Wgt_3_445,Wgt_3_446,Wgt_3_447,Wgt_3_448,Wgt_3_449,Wgt_3_450,Wgt_3_451,Wgt_3_452,Wgt_3_453,Wgt_3_454,Wgt_3_455,Wgt_3_456,Wgt_3_457,Wgt_3_458,Wgt_3_459,Wgt_3_460,Wgt_3_461,Wgt_3_462,Wgt_3_463,Wgt_3_464,Wgt_3_465,Wgt_3_466,Wgt_3_467,Wgt_3_468,Wgt_3_469,Wgt_3_470,Wgt_3_471,Wgt_3_472,Wgt_3_473,Wgt_3_474,Wgt_3_475,Wgt_3_476,Wgt_3_477,Wgt_3_478,Wgt_3_479,Wgt_3_480,Wgt_3_481,Wgt_3_482,Wgt_3_483,Wgt_3_484,Wgt_3_485,Wgt_3_486,Wgt_3_487,Wgt_3_488,Wgt_3_489,Wgt_3_490,Wgt_3_491,Wgt_3_492,Wgt_3_493,Wgt_3_494,Wgt_3_495,Wgt_3_496,Wgt_3_497,Wgt_3_498,Wgt_3_499,Wgt_3_500,Wgt_3_501,Wgt_3_502,Wgt_3_503,Wgt_3_504,Wgt_3_505,Wgt_3_506,Wgt_3_507,Wgt_3_508,Wgt_3_509,Wgt_3_510,Wgt_3_511,Wgt_3_512,Wgt_3_513,Wgt_3_514,Wgt_3_515,Wgt_3_516,Wgt_3_517,Wgt_3_518,Wgt_3_519,Wgt_3_520,Wgt_3_521,Wgt_3_522,Wgt_3_523,Wgt_3_524,Wgt_3_525,Wgt_3_526,Wgt_3_527,Wgt_3_528,Wgt_3_529,Wgt_3_530,Wgt_3_531,Wgt_3_532,Wgt_3_533,Wgt_3_534,Wgt_3_535,Wgt_3_536,Wgt_3_537,Wgt_3_538,Wgt_3_539,Wgt_3_540,Wgt_3_541,Wgt_3_542,Wgt_3_543,Wgt_3_544,Wgt_3_545,Wgt_3_546,Wgt_3_547,Wgt_3_548,Wgt_3_549,Wgt_3_550,Wgt_3_551,Wgt_3_552,Wgt_3_553,Wgt_3_554,Wgt_3_555,Wgt_3_556,Wgt_3_557,Wgt_3_558,Wgt_3_559,Wgt_3_560,Wgt_3_561,Wgt_3_562,Wgt_3_563,Wgt_3_564,Wgt_3_565,Wgt_3_566,Wgt_3_567,Wgt_3_568,Wgt_3_569,Wgt_3_570,Wgt_3_571,Wgt_3_572,Wgt_3_573,Wgt_3_574,Wgt_3_575,Wgt_3_576,Wgt_3_577,Wgt_3_578,Wgt_3_579,Wgt_3_580,Wgt_3_581,Wgt_3_582,Wgt_3_583,Wgt_3_584,Wgt_3_585,Wgt_3_586,Wgt_3_587,Wgt_3_588,Wgt_3_589,Wgt_3_590,Wgt_3_591,Wgt_3_592,Wgt_3_593,Wgt_3_594,Wgt_3_595,Wgt_3_596,Wgt_3_597,Wgt_3_598,Wgt_3_599,Wgt_3_600,Wgt_3_601,Wgt_3_602,Wgt_3_603,Wgt_3_604,Wgt_3_605,Wgt_3_606,Wgt_3_607,Wgt_3_608,Wgt_3_609,Wgt_3_610,Wgt_3_611,Wgt_3_612,Wgt_3_613,Wgt_3_614,Wgt_3_615,Wgt_3_616,Wgt_3_617,Wgt_3_618,Wgt_3_619,Wgt_3_620,Wgt_3_621,Wgt_3_622,Wgt_3_623,Wgt_3_624,Wgt_3_625,Wgt_3_626,Wgt_3_627,Wgt_3_628,Wgt_3_629,Wgt_3_630,Wgt_3_631,Wgt_3_632,Wgt_3_633,Wgt_3_634,Wgt_3_635,Wgt_3_636,Wgt_3_637,Wgt_3_638,Wgt_3_639,Wgt_3_640,Wgt_3_641,Wgt_3_642,Wgt_3_643,Wgt_3_644,Wgt_3_645,Wgt_3_646,Wgt_3_647,Wgt_3_648,Wgt_3_649,Wgt_3_650,Wgt_3_651,Wgt_3_652,Wgt_3_653,Wgt_3_654,Wgt_3_655,Wgt_3_656,Wgt_3_657,Wgt_3_658,Wgt_3_659,Wgt_3_660,Wgt_3_661,Wgt_3_662,Wgt_3_663,Wgt_3_664,Wgt_3_665,Wgt_3_666,Wgt_3_667,Wgt_3_668,Wgt_3_669,Wgt_3_670,Wgt_3_671,Wgt_3_672,Wgt_3_673,Wgt_3_674,Wgt_3_675,Wgt_3_676,Wgt_3_677,Wgt_3_678,Wgt_3_679,Wgt_3_680,Wgt_3_681,Wgt_3_682,Wgt_3_683,Wgt_3_684,Wgt_3_685,Wgt_3_686,Wgt_3_687,Wgt_3_688,Wgt_3_689,Wgt_3_690,Wgt_3_691,Wgt_3_692,Wgt_3_693,Wgt_3_694,Wgt_3_695,Wgt_3_696,Wgt_3_697,Wgt_3_698,Wgt_3_699,Wgt_3_700,Wgt_3_701,Wgt_3_702,Wgt_3_703,Wgt_3_704,Wgt_3_705,Wgt_3_706,Wgt_3_707,Wgt_3_708,Wgt_3_709,Wgt_3_710,Wgt_3_711,Wgt_3_712,Wgt_3_713,Wgt_3_714,Wgt_3_715,Wgt_3_716,Wgt_3_717,Wgt_3_718,Wgt_3_719,Wgt_3_720,Wgt_3_721,Wgt_3_722,Wgt_3_723,Wgt_3_724,Wgt_3_725,Wgt_3_726,Wgt_3_727,Wgt_3_728,Wgt_3_729,Wgt_3_730,Wgt_3_731,Wgt_3_732,Wgt_3_733,Wgt_3_734,Wgt_3_735,Wgt_3_736,Wgt_3_737,Wgt_3_738,Wgt_3_739,Wgt_3_740,Wgt_3_741,Wgt_3_742,Wgt_3_743,Wgt_3_744,Wgt_3_745,Wgt_3_746,Wgt_3_747,Wgt_3_748,Wgt_3_749,Wgt_3_750,Wgt_3_751,Wgt_3_752,Wgt_3_753,Wgt_3_754,Wgt_3_755,Wgt_3_756,Wgt_3_757,Wgt_3_758,Wgt_3_759,Wgt_3_760,Wgt_3_761,Wgt_3_762,Wgt_3_763,Wgt_3_764,Wgt_3_765,Wgt_3_766,Wgt_3_767,Wgt_3_768,Wgt_3_769,Wgt_3_770,Wgt_3_771,Wgt_3_772,Wgt_3_773,Wgt_3_774,Wgt_3_775,Wgt_3_776,Wgt_3_777,Wgt_3_778,Wgt_3_779,Wgt_3_780,Wgt_3_781,Wgt_3_782,Wgt_3_783,Wgt_3_784,Wgt_4_0,Wgt_4_1,Wgt_4_2,Wgt_4_3,Wgt_4_4,Wgt_4_5,Wgt_4_6,Wgt_4_7,Wgt_4_8,Wgt_4_9,Wgt_4_10,Wgt_4_11,Wgt_4_12,Wgt_4_13,Wgt_4_14,Wgt_4_15,Wgt_4_16,Wgt_4_17,Wgt_4_18,Wgt_4_19,Wgt_4_20,Wgt_4_21,Wgt_4_22,Wgt_4_23,Wgt_4_24,Wgt_4_25,Wgt_4_26,Wgt_4_27,Wgt_4_28,Wgt_4_29,Wgt_4_30,Wgt_4_31,Wgt_4_32,Wgt_4_33,Wgt_4_34,Wgt_4_35,Wgt_4_36,Wgt_4_37,Wgt_4_38,Wgt_4_39,Wgt_4_40,Wgt_4_41,Wgt_4_42,Wgt_4_43,Wgt_4_44,Wgt_4_45,Wgt_4_46,Wgt_4_47,Wgt_4_48,Wgt_4_49,Wgt_4_50,Wgt_4_51,Wgt_4_52,Wgt_4_53,Wgt_4_54,Wgt_4_55,Wgt_4_56,Wgt_4_57,Wgt_4_58,Wgt_4_59,Wgt_4_60,Wgt_4_61,Wgt_4_62,Wgt_4_63,Wgt_4_64,Wgt_4_65,Wgt_4_66,Wgt_4_67,Wgt_4_68,Wgt_4_69,Wgt_4_70,Wgt_4_71,Wgt_4_72,Wgt_4_73,Wgt_4_74,Wgt_4_75,Wgt_4_76,Wgt_4_77,Wgt_4_78,Wgt_4_79,Wgt_4_80,Wgt_4_81,Wgt_4_82,Wgt_4_83,Wgt_4_84,Wgt_4_85,Wgt_4_86,Wgt_4_87,Wgt_4_88,Wgt_4_89,Wgt_4_90,Wgt_4_91,Wgt_4_92,Wgt_4_93,Wgt_4_94,Wgt_4_95,Wgt_4_96,Wgt_4_97,Wgt_4_98,Wgt_4_99,Wgt_4_100,Wgt_4_101,Wgt_4_102,Wgt_4_103,Wgt_4_104,Wgt_4_105,Wgt_4_106,Wgt_4_107,Wgt_4_108,Wgt_4_109,Wgt_4_110,Wgt_4_111,Wgt_4_112,Wgt_4_113,Wgt_4_114,Wgt_4_115,Wgt_4_116,Wgt_4_117,Wgt_4_118,Wgt_4_119,Wgt_4_120,Wgt_4_121,Wgt_4_122,Wgt_4_123,Wgt_4_124,Wgt_4_125,Wgt_4_126,Wgt_4_127,Wgt_4_128,Wgt_4_129,Wgt_4_130,Wgt_4_131,Wgt_4_132,Wgt_4_133,Wgt_4_134,Wgt_4_135,Wgt_4_136,Wgt_4_137,Wgt_4_138,Wgt_4_139,Wgt_4_140,Wgt_4_141,Wgt_4_142,Wgt_4_143,Wgt_4_144,Wgt_4_145,Wgt_4_146,Wgt_4_147,Wgt_4_148,Wgt_4_149,Wgt_4_150,Wgt_4_151,Wgt_4_152,Wgt_4_153,Wgt_4_154,Wgt_4_155,Wgt_4_156,Wgt_4_157,Wgt_4_158,Wgt_4_159,Wgt_4_160,Wgt_4_161,Wgt_4_162,Wgt_4_163,Wgt_4_164,Wgt_4_165,Wgt_4_166,Wgt_4_167,Wgt_4_168,Wgt_4_169,Wgt_4_170,Wgt_4_171,Wgt_4_172,Wgt_4_173,Wgt_4_174,Wgt_4_175,Wgt_4_176,Wgt_4_177,Wgt_4_178,Wgt_4_179,Wgt_4_180,Wgt_4_181,Wgt_4_182,Wgt_4_183,Wgt_4_184,Wgt_4_185,Wgt_4_186,Wgt_4_187,Wgt_4_188,Wgt_4_189,Wgt_4_190,Wgt_4_191,Wgt_4_192,Wgt_4_193,Wgt_4_194,Wgt_4_195,Wgt_4_196,Wgt_4_197,Wgt_4_198,Wgt_4_199,Wgt_4_200,Wgt_4_201,Wgt_4_202,Wgt_4_203,Wgt_4_204,Wgt_4_205,Wgt_4_206,Wgt_4_207,Wgt_4_208,Wgt_4_209,Wgt_4_210,Wgt_4_211,Wgt_4_212,Wgt_4_213,Wgt_4_214,Wgt_4_215,Wgt_4_216,Wgt_4_217,Wgt_4_218,Wgt_4_219,Wgt_4_220,Wgt_4_221,Wgt_4_222,Wgt_4_223,Wgt_4_224,Wgt_4_225,Wgt_4_226,Wgt_4_227,Wgt_4_228,Wgt_4_229,Wgt_4_230,Wgt_4_231,Wgt_4_232,Wgt_4_233,Wgt_4_234,Wgt_4_235,Wgt_4_236,Wgt_4_237,Wgt_4_238,Wgt_4_239,Wgt_4_240,Wgt_4_241,Wgt_4_242,Wgt_4_243,Wgt_4_244,Wgt_4_245,Wgt_4_246,Wgt_4_247,Wgt_4_248,Wgt_4_249,Wgt_4_250,Wgt_4_251,Wgt_4_252,Wgt_4_253,Wgt_4_254,Wgt_4_255,Wgt_4_256,Wgt_4_257,Wgt_4_258,Wgt_4_259,Wgt_4_260,Wgt_4_261,Wgt_4_262,Wgt_4_263,Wgt_4_264,Wgt_4_265,Wgt_4_266,Wgt_4_267,Wgt_4_268,Wgt_4_269,Wgt_4_270,Wgt_4_271,Wgt_4_272,Wgt_4_273,Wgt_4_274,Wgt_4_275,Wgt_4_276,Wgt_4_277,Wgt_4_278,Wgt_4_279,Wgt_4_280,Wgt_4_281,Wgt_4_282,Wgt_4_283,Wgt_4_284,Wgt_4_285,Wgt_4_286,Wgt_4_287,Wgt_4_288,Wgt_4_289,Wgt_4_290,Wgt_4_291,Wgt_4_292,Wgt_4_293,Wgt_4_294,Wgt_4_295,Wgt_4_296,Wgt_4_297,Wgt_4_298,Wgt_4_299,Wgt_4_300,Wgt_4_301,Wgt_4_302,Wgt_4_303,Wgt_4_304,Wgt_4_305,Wgt_4_306,Wgt_4_307,Wgt_4_308,Wgt_4_309,Wgt_4_310,Wgt_4_311,Wgt_4_312,Wgt_4_313,Wgt_4_314,Wgt_4_315,Wgt_4_316,Wgt_4_317,Wgt_4_318,Wgt_4_319,Wgt_4_320,Wgt_4_321,Wgt_4_322,Wgt_4_323,Wgt_4_324,Wgt_4_325,Wgt_4_326,Wgt_4_327,Wgt_4_328,Wgt_4_329,Wgt_4_330,Wgt_4_331,Wgt_4_332,Wgt_4_333,Wgt_4_334,Wgt_4_335,Wgt_4_336,Wgt_4_337,Wgt_4_338,Wgt_4_339,Wgt_4_340,Wgt_4_341,Wgt_4_342,Wgt_4_343,Wgt_4_344,Wgt_4_345,Wgt_4_346,Wgt_4_347,Wgt_4_348,Wgt_4_349,Wgt_4_350,Wgt_4_351,Wgt_4_352,Wgt_4_353,Wgt_4_354,Wgt_4_355,Wgt_4_356,Wgt_4_357,Wgt_4_358,Wgt_4_359,Wgt_4_360,Wgt_4_361,Wgt_4_362,Wgt_4_363,Wgt_4_364,Wgt_4_365,Wgt_4_366,Wgt_4_367,Wgt_4_368,Wgt_4_369,Wgt_4_370,Wgt_4_371,Wgt_4_372,Wgt_4_373,Wgt_4_374,Wgt_4_375,Wgt_4_376,Wgt_4_377,Wgt_4_378,Wgt_4_379,Wgt_4_380,Wgt_4_381,Wgt_4_382,Wgt_4_383,Wgt_4_384,Wgt_4_385,Wgt_4_386,Wgt_4_387,Wgt_4_388,Wgt_4_389,Wgt_4_390,Wgt_4_391,Wgt_4_392,Wgt_4_393,Wgt_4_394,Wgt_4_395,Wgt_4_396,Wgt_4_397,Wgt_4_398,Wgt_4_399,Wgt_4_400,Wgt_4_401,Wgt_4_402,Wgt_4_403,Wgt_4_404,Wgt_4_405,Wgt_4_406,Wgt_4_407,Wgt_4_408,Wgt_4_409,Wgt_4_410,Wgt_4_411,Wgt_4_412,Wgt_4_413,Wgt_4_414,Wgt_4_415,Wgt_4_416,Wgt_4_417,Wgt_4_418,Wgt_4_419,Wgt_4_420,Wgt_4_421,Wgt_4_422,Wgt_4_423,Wgt_4_424,Wgt_4_425,Wgt_4_426,Wgt_4_427,Wgt_4_428,Wgt_4_429,Wgt_4_430,Wgt_4_431,Wgt_4_432,Wgt_4_433,Wgt_4_434,Wgt_4_435,Wgt_4_436,Wgt_4_437,Wgt_4_438,Wgt_4_439,Wgt_4_440,Wgt_4_441,Wgt_4_442,Wgt_4_443,Wgt_4_444,Wgt_4_445,Wgt_4_446,Wgt_4_447,Wgt_4_448,Wgt_4_449,Wgt_4_450,Wgt_4_451,Wgt_4_452,Wgt_4_453,Wgt_4_454,Wgt_4_455,Wgt_4_456,Wgt_4_457,Wgt_4_458,Wgt_4_459,Wgt_4_460,Wgt_4_461,Wgt_4_462,Wgt_4_463,Wgt_4_464,Wgt_4_465,Wgt_4_466,Wgt_4_467,Wgt_4_468,Wgt_4_469,Wgt_4_470,Wgt_4_471,Wgt_4_472,Wgt_4_473,Wgt_4_474,Wgt_4_475,Wgt_4_476,Wgt_4_477,Wgt_4_478,Wgt_4_479,Wgt_4_480,Wgt_4_481,Wgt_4_482,Wgt_4_483,Wgt_4_484,Wgt_4_485,Wgt_4_486,Wgt_4_487,Wgt_4_488,Wgt_4_489,Wgt_4_490,Wgt_4_491,Wgt_4_492,Wgt_4_493,Wgt_4_494,Wgt_4_495,Wgt_4_496,Wgt_4_497,Wgt_4_498,Wgt_4_499,Wgt_4_500,Wgt_4_501,Wgt_4_502,Wgt_4_503,Wgt_4_504,Wgt_4_505,Wgt_4_506,Wgt_4_507,Wgt_4_508,Wgt_4_509,Wgt_4_510,Wgt_4_511,Wgt_4_512,Wgt_4_513,Wgt_4_514,Wgt_4_515,Wgt_4_516,Wgt_4_517,Wgt_4_518,Wgt_4_519,Wgt_4_520,Wgt_4_521,Wgt_4_522,Wgt_4_523,Wgt_4_524,Wgt_4_525,Wgt_4_526,Wgt_4_527,Wgt_4_528,Wgt_4_529,Wgt_4_530,Wgt_4_531,Wgt_4_532,Wgt_4_533,Wgt_4_534,Wgt_4_535,Wgt_4_536,Wgt_4_537,Wgt_4_538,Wgt_4_539,Wgt_4_540,Wgt_4_541,Wgt_4_542,Wgt_4_543,Wgt_4_544,Wgt_4_545,Wgt_4_546,Wgt_4_547,Wgt_4_548,Wgt_4_549,Wgt_4_550,Wgt_4_551,Wgt_4_552,Wgt_4_553,Wgt_4_554,Wgt_4_555,Wgt_4_556,Wgt_4_557,Wgt_4_558,Wgt_4_559,Wgt_4_560,Wgt_4_561,Wgt_4_562,Wgt_4_563,Wgt_4_564,Wgt_4_565,Wgt_4_566,Wgt_4_567,Wgt_4_568,Wgt_4_569,Wgt_4_570,Wgt_4_571,Wgt_4_572,Wgt_4_573,Wgt_4_574,Wgt_4_575,Wgt_4_576,Wgt_4_577,Wgt_4_578,Wgt_4_579,Wgt_4_580,Wgt_4_581,Wgt_4_582,Wgt_4_583,Wgt_4_584,Wgt_4_585,Wgt_4_586,Wgt_4_587,Wgt_4_588,Wgt_4_589,Wgt_4_590,Wgt_4_591,Wgt_4_592,Wgt_4_593,Wgt_4_594,Wgt_4_595,Wgt_4_596,Wgt_4_597,Wgt_4_598,Wgt_4_599,Wgt_4_600,Wgt_4_601,Wgt_4_602,Wgt_4_603,Wgt_4_604,Wgt_4_605,Wgt_4_606,Wgt_4_607,Wgt_4_608,Wgt_4_609,Wgt_4_610,Wgt_4_611,Wgt_4_612,Wgt_4_613,Wgt_4_614,Wgt_4_615,Wgt_4_616,Wgt_4_617,Wgt_4_618,Wgt_4_619,Wgt_4_620,Wgt_4_621,Wgt_4_622,Wgt_4_623,Wgt_4_624,Wgt_4_625,Wgt_4_626,Wgt_4_627,Wgt_4_628,Wgt_4_629,Wgt_4_630,Wgt_4_631,Wgt_4_632,Wgt_4_633,Wgt_4_634,Wgt_4_635,Wgt_4_636,Wgt_4_637,Wgt_4_638,Wgt_4_639,Wgt_4_640,Wgt_4_641,Wgt_4_642,Wgt_4_643,Wgt_4_644,Wgt_4_645,Wgt_4_646,Wgt_4_647,Wgt_4_648,Wgt_4_649,Wgt_4_650,Wgt_4_651,Wgt_4_652,Wgt_4_653,Wgt_4_654,Wgt_4_655,Wgt_4_656,Wgt_4_657,Wgt_4_658,Wgt_4_659,Wgt_4_660,Wgt_4_661,Wgt_4_662,Wgt_4_663,Wgt_4_664,Wgt_4_665,Wgt_4_666,Wgt_4_667,Wgt_4_668,Wgt_4_669,Wgt_4_670,Wgt_4_671,Wgt_4_672,Wgt_4_673,Wgt_4_674,Wgt_4_675,Wgt_4_676,Wgt_4_677,Wgt_4_678,Wgt_4_679,Wgt_4_680,Wgt_4_681,Wgt_4_682,Wgt_4_683,Wgt_4_684,Wgt_4_685,Wgt_4_686,Wgt_4_687,Wgt_4_688,Wgt_4_689,Wgt_4_690,Wgt_4_691,Wgt_4_692,Wgt_4_693,Wgt_4_694,Wgt_4_695,Wgt_4_696,Wgt_4_697,Wgt_4_698,Wgt_4_699,Wgt_4_700,Wgt_4_701,Wgt_4_702,Wgt_4_703,Wgt_4_704,Wgt_4_705,Wgt_4_706,Wgt_4_707,Wgt_4_708,Wgt_4_709,Wgt_4_710,Wgt_4_711,Wgt_4_712,Wgt_4_713,Wgt_4_714,Wgt_4_715,Wgt_4_716,Wgt_4_717,Wgt_4_718,Wgt_4_719,Wgt_4_720,Wgt_4_721,Wgt_4_722,Wgt_4_723,Wgt_4_724,Wgt_4_725,Wgt_4_726,Wgt_4_727,Wgt_4_728,Wgt_4_729,Wgt_4_730,Wgt_4_731,Wgt_4_732,Wgt_4_733,Wgt_4_734,Wgt_4_735,Wgt_4_736,Wgt_4_737,Wgt_4_738,Wgt_4_739,Wgt_4_740,Wgt_4_741,Wgt_4_742,Wgt_4_743,Wgt_4_744,Wgt_4_745,Wgt_4_746,Wgt_4_747,Wgt_4_748,Wgt_4_749,Wgt_4_750,Wgt_4_751,Wgt_4_752,Wgt_4_753,Wgt_4_754,Wgt_4_755,Wgt_4_756,Wgt_4_757,Wgt_4_758,Wgt_4_759,Wgt_4_760,Wgt_4_761,Wgt_4_762,Wgt_4_763,Wgt_4_764,Wgt_4_765,Wgt_4_766,Wgt_4_767,Wgt_4_768,Wgt_4_769,Wgt_4_770,Wgt_4_771,Wgt_4_772,Wgt_4_773,Wgt_4_774,Wgt_4_775,Wgt_4_776,Wgt_4_777,Wgt_4_778,Wgt_4_779,Wgt_4_780,Wgt_4_781,Wgt_4_782,Wgt_4_783,Wgt_4_784,Wgt_5_0,Wgt_5_1,Wgt_5_2,Wgt_5_3,Wgt_5_4,Wgt_5_5,Wgt_5_6,Wgt_5_7,Wgt_5_8,Wgt_5_9,Wgt_5_10,Wgt_5_11,Wgt_5_12,Wgt_5_13,Wgt_5_14,Wgt_5_15,Wgt_5_16,Wgt_5_17,Wgt_5_18,Wgt_5_19,Wgt_5_20,Wgt_5_21,Wgt_5_22,Wgt_5_23,Wgt_5_24,Wgt_5_25,Wgt_5_26,Wgt_5_27,Wgt_5_28,Wgt_5_29,Wgt_5_30,Wgt_5_31,Wgt_5_32,Wgt_5_33,Wgt_5_34,Wgt_5_35,Wgt_5_36,Wgt_5_37,Wgt_5_38,Wgt_5_39,Wgt_5_40,Wgt_5_41,Wgt_5_42,Wgt_5_43,Wgt_5_44,Wgt_5_45,Wgt_5_46,Wgt_5_47,Wgt_5_48,Wgt_5_49,Wgt_5_50,Wgt_5_51,Wgt_5_52,Wgt_5_53,Wgt_5_54,Wgt_5_55,Wgt_5_56,Wgt_5_57,Wgt_5_58,Wgt_5_59,Wgt_5_60,Wgt_5_61,Wgt_5_62,Wgt_5_63,Wgt_5_64,Wgt_5_65,Wgt_5_66,Wgt_5_67,Wgt_5_68,Wgt_5_69,Wgt_5_70,Wgt_5_71,Wgt_5_72,Wgt_5_73,Wgt_5_74,Wgt_5_75,Wgt_5_76,Wgt_5_77,Wgt_5_78,Wgt_5_79,Wgt_5_80,Wgt_5_81,Wgt_5_82,Wgt_5_83,Wgt_5_84,Wgt_5_85,Wgt_5_86,Wgt_5_87,Wgt_5_88,Wgt_5_89,Wgt_5_90,Wgt_5_91,Wgt_5_92,Wgt_5_93,Wgt_5_94,Wgt_5_95,Wgt_5_96,Wgt_5_97,Wgt_5_98,Wgt_5_99,Wgt_5_100,Wgt_5_101,Wgt_5_102,Wgt_5_103,Wgt_5_104,Wgt_5_105,Wgt_5_106,Wgt_5_107,Wgt_5_108,Wgt_5_109,Wgt_5_110,Wgt_5_111,Wgt_5_112,Wgt_5_113,Wgt_5_114,Wgt_5_115,Wgt_5_116,Wgt_5_117,Wgt_5_118,Wgt_5_119,Wgt_5_120,Wgt_5_121,Wgt_5_122,Wgt_5_123,Wgt_5_124,Wgt_5_125,Wgt_5_126,Wgt_5_127,Wgt_5_128,Wgt_5_129,Wgt_5_130,Wgt_5_131,Wgt_5_132,Wgt_5_133,Wgt_5_134,Wgt_5_135,Wgt_5_136,Wgt_5_137,Wgt_5_138,Wgt_5_139,Wgt_5_140,Wgt_5_141,Wgt_5_142,Wgt_5_143,Wgt_5_144,Wgt_5_145,Wgt_5_146,Wgt_5_147,Wgt_5_148,Wgt_5_149,Wgt_5_150,Wgt_5_151,Wgt_5_152,Wgt_5_153,Wgt_5_154,Wgt_5_155,Wgt_5_156,Wgt_5_157,Wgt_5_158,Wgt_5_159,Wgt_5_160,Wgt_5_161,Wgt_5_162,Wgt_5_163,Wgt_5_164,Wgt_5_165,Wgt_5_166,Wgt_5_167,Wgt_5_168,Wgt_5_169,Wgt_5_170,Wgt_5_171,Wgt_5_172,Wgt_5_173,Wgt_5_174,Wgt_5_175,Wgt_5_176,Wgt_5_177,Wgt_5_178,Wgt_5_179,Wgt_5_180,Wgt_5_181,Wgt_5_182,Wgt_5_183,Wgt_5_184,Wgt_5_185,Wgt_5_186,Wgt_5_187,Wgt_5_188,Wgt_5_189,Wgt_5_190,Wgt_5_191,Wgt_5_192,Wgt_5_193,Wgt_5_194,Wgt_5_195,Wgt_5_196,Wgt_5_197,Wgt_5_198,Wgt_5_199,Wgt_5_200,Wgt_5_201,Wgt_5_202,Wgt_5_203,Wgt_5_204,Wgt_5_205,Wgt_5_206,Wgt_5_207,Wgt_5_208,Wgt_5_209,Wgt_5_210,Wgt_5_211,Wgt_5_212,Wgt_5_213,Wgt_5_214,Wgt_5_215,Wgt_5_216,Wgt_5_217,Wgt_5_218,Wgt_5_219,Wgt_5_220,Wgt_5_221,Wgt_5_222,Wgt_5_223,Wgt_5_224,Wgt_5_225,Wgt_5_226,Wgt_5_227,Wgt_5_228,Wgt_5_229,Wgt_5_230,Wgt_5_231,Wgt_5_232,Wgt_5_233,Wgt_5_234,Wgt_5_235,Wgt_5_236,Wgt_5_237,Wgt_5_238,Wgt_5_239,Wgt_5_240,Wgt_5_241,Wgt_5_242,Wgt_5_243,Wgt_5_244,Wgt_5_245,Wgt_5_246,Wgt_5_247,Wgt_5_248,Wgt_5_249,Wgt_5_250,Wgt_5_251,Wgt_5_252,Wgt_5_253,Wgt_5_254,Wgt_5_255,Wgt_5_256,Wgt_5_257,Wgt_5_258,Wgt_5_259,Wgt_5_260,Wgt_5_261,Wgt_5_262,Wgt_5_263,Wgt_5_264,Wgt_5_265,Wgt_5_266,Wgt_5_267,Wgt_5_268,Wgt_5_269,Wgt_5_270,Wgt_5_271,Wgt_5_272,Wgt_5_273,Wgt_5_274,Wgt_5_275,Wgt_5_276,Wgt_5_277,Wgt_5_278,Wgt_5_279,Wgt_5_280,Wgt_5_281,Wgt_5_282,Wgt_5_283,Wgt_5_284,Wgt_5_285,Wgt_5_286,Wgt_5_287,Wgt_5_288,Wgt_5_289,Wgt_5_290,Wgt_5_291,Wgt_5_292,Wgt_5_293,Wgt_5_294,Wgt_5_295,Wgt_5_296,Wgt_5_297,Wgt_5_298,Wgt_5_299,Wgt_5_300,Wgt_5_301,Wgt_5_302,Wgt_5_303,Wgt_5_304,Wgt_5_305,Wgt_5_306,Wgt_5_307,Wgt_5_308,Wgt_5_309,Wgt_5_310,Wgt_5_311,Wgt_5_312,Wgt_5_313,Wgt_5_314,Wgt_5_315,Wgt_5_316,Wgt_5_317,Wgt_5_318,Wgt_5_319,Wgt_5_320,Wgt_5_321,Wgt_5_322,Wgt_5_323,Wgt_5_324,Wgt_5_325,Wgt_5_326,Wgt_5_327,Wgt_5_328,Wgt_5_329,Wgt_5_330,Wgt_5_331,Wgt_5_332,Wgt_5_333,Wgt_5_334,Wgt_5_335,Wgt_5_336,Wgt_5_337,Wgt_5_338,Wgt_5_339,Wgt_5_340,Wgt_5_341,Wgt_5_342,Wgt_5_343,Wgt_5_344,Wgt_5_345,Wgt_5_346,Wgt_5_347,Wgt_5_348,Wgt_5_349,Wgt_5_350,Wgt_5_351,Wgt_5_352,Wgt_5_353,Wgt_5_354,Wgt_5_355,Wgt_5_356,Wgt_5_357,Wgt_5_358,Wgt_5_359,Wgt_5_360,Wgt_5_361,Wgt_5_362,Wgt_5_363,Wgt_5_364,Wgt_5_365,Wgt_5_366,Wgt_5_367,Wgt_5_368,Wgt_5_369,Wgt_5_370,Wgt_5_371,Wgt_5_372,Wgt_5_373,Wgt_5_374,Wgt_5_375,Wgt_5_376,Wgt_5_377,Wgt_5_378,Wgt_5_379,Wgt_5_380,Wgt_5_381,Wgt_5_382,Wgt_5_383,Wgt_5_384,Wgt_5_385,Wgt_5_386,Wgt_5_387,Wgt_5_388,Wgt_5_389,Wgt_5_390,Wgt_5_391,Wgt_5_392,Wgt_5_393,Wgt_5_394,Wgt_5_395,Wgt_5_396,Wgt_5_397,Wgt_5_398,Wgt_5_399,Wgt_5_400,Wgt_5_401,Wgt_5_402,Wgt_5_403,Wgt_5_404,Wgt_5_405,Wgt_5_406,Wgt_5_407,Wgt_5_408,Wgt_5_409,Wgt_5_410,Wgt_5_411,Wgt_5_412,Wgt_5_413,Wgt_5_414,Wgt_5_415,Wgt_5_416,Wgt_5_417,Wgt_5_418,Wgt_5_419,Wgt_5_420,Wgt_5_421,Wgt_5_422,Wgt_5_423,Wgt_5_424,Wgt_5_425,Wgt_5_426,Wgt_5_427,Wgt_5_428,Wgt_5_429,Wgt_5_430,Wgt_5_431,Wgt_5_432,Wgt_5_433,Wgt_5_434,Wgt_5_435,Wgt_5_436,Wgt_5_437,Wgt_5_438,Wgt_5_439,Wgt_5_440,Wgt_5_441,Wgt_5_442,Wgt_5_443,Wgt_5_444,Wgt_5_445,Wgt_5_446,Wgt_5_447,Wgt_5_448,Wgt_5_449,Wgt_5_450,Wgt_5_451,Wgt_5_452,Wgt_5_453,Wgt_5_454,Wgt_5_455,Wgt_5_456,Wgt_5_457,Wgt_5_458,Wgt_5_459,Wgt_5_460,Wgt_5_461,Wgt_5_462,Wgt_5_463,Wgt_5_464,Wgt_5_465,Wgt_5_466,Wgt_5_467,Wgt_5_468,Wgt_5_469,Wgt_5_470,Wgt_5_471,Wgt_5_472,Wgt_5_473,Wgt_5_474,Wgt_5_475,Wgt_5_476,Wgt_5_477,Wgt_5_478,Wgt_5_479,Wgt_5_480,Wgt_5_481,Wgt_5_482,Wgt_5_483,Wgt_5_484,Wgt_5_485,Wgt_5_486,Wgt_5_487,Wgt_5_488,Wgt_5_489,Wgt_5_490,Wgt_5_491,Wgt_5_492,Wgt_5_493,Wgt_5_494,Wgt_5_495,Wgt_5_496,Wgt_5_497,Wgt_5_498,Wgt_5_499,Wgt_5_500,Wgt_5_501,Wgt_5_502,Wgt_5_503,Wgt_5_504,Wgt_5_505,Wgt_5_506,Wgt_5_507,Wgt_5_508,Wgt_5_509,Wgt_5_510,Wgt_5_511,Wgt_5_512,Wgt_5_513,Wgt_5_514,Wgt_5_515,Wgt_5_516,Wgt_5_517,Wgt_5_518,Wgt_5_519,Wgt_5_520,Wgt_5_521,Wgt_5_522,Wgt_5_523,Wgt_5_524,Wgt_5_525,Wgt_5_526,Wgt_5_527,Wgt_5_528,Wgt_5_529,Wgt_5_530,Wgt_5_531,Wgt_5_532,Wgt_5_533,Wgt_5_534,Wgt_5_535,Wgt_5_536,Wgt_5_537,Wgt_5_538,Wgt_5_539,Wgt_5_540,Wgt_5_541,Wgt_5_542,Wgt_5_543,Wgt_5_544,Wgt_5_545,Wgt_5_546,Wgt_5_547,Wgt_5_548,Wgt_5_549,Wgt_5_550,Wgt_5_551,Wgt_5_552,Wgt_5_553,Wgt_5_554,Wgt_5_555,Wgt_5_556,Wgt_5_557,Wgt_5_558,Wgt_5_559,Wgt_5_560,Wgt_5_561,Wgt_5_562,Wgt_5_563,Wgt_5_564,Wgt_5_565,Wgt_5_566,Wgt_5_567,Wgt_5_568,Wgt_5_569,Wgt_5_570,Wgt_5_571,Wgt_5_572,Wgt_5_573,Wgt_5_574,Wgt_5_575,Wgt_5_576,Wgt_5_577,Wgt_5_578,Wgt_5_579,Wgt_5_580,Wgt_5_581,Wgt_5_582,Wgt_5_583,Wgt_5_584,Wgt_5_585,Wgt_5_586,Wgt_5_587,Wgt_5_588,Wgt_5_589,Wgt_5_590,Wgt_5_591,Wgt_5_592,Wgt_5_593,Wgt_5_594,Wgt_5_595,Wgt_5_596,Wgt_5_597,Wgt_5_598,Wgt_5_599,Wgt_5_600,Wgt_5_601,Wgt_5_602,Wgt_5_603,Wgt_5_604,Wgt_5_605,Wgt_5_606,Wgt_5_607,Wgt_5_608,Wgt_5_609,Wgt_5_610,Wgt_5_611,Wgt_5_612,Wgt_5_613,Wgt_5_614,Wgt_5_615,Wgt_5_616,Wgt_5_617,Wgt_5_618,Wgt_5_619,Wgt_5_620,Wgt_5_621,Wgt_5_622,Wgt_5_623,Wgt_5_624,Wgt_5_625,Wgt_5_626,Wgt_5_627,Wgt_5_628,Wgt_5_629,Wgt_5_630,Wgt_5_631,Wgt_5_632,Wgt_5_633,Wgt_5_634,Wgt_5_635,Wgt_5_636,Wgt_5_637,Wgt_5_638,Wgt_5_639,Wgt_5_640,Wgt_5_641,Wgt_5_642,Wgt_5_643,Wgt_5_644,Wgt_5_645,Wgt_5_646,Wgt_5_647,Wgt_5_648,Wgt_5_649,Wgt_5_650,Wgt_5_651,Wgt_5_652,Wgt_5_653,Wgt_5_654,Wgt_5_655,Wgt_5_656,Wgt_5_657,Wgt_5_658,Wgt_5_659,Wgt_5_660,Wgt_5_661,Wgt_5_662,Wgt_5_663,Wgt_5_664,Wgt_5_665,Wgt_5_666,Wgt_5_667,Wgt_5_668,Wgt_5_669,Wgt_5_670,Wgt_5_671,Wgt_5_672,Wgt_5_673,Wgt_5_674,Wgt_5_675,Wgt_5_676,Wgt_5_677,Wgt_5_678,Wgt_5_679,Wgt_5_680,Wgt_5_681,Wgt_5_682,Wgt_5_683,Wgt_5_684,Wgt_5_685,Wgt_5_686,Wgt_5_687,Wgt_5_688,Wgt_5_689,Wgt_5_690,Wgt_5_691,Wgt_5_692,Wgt_5_693,Wgt_5_694,Wgt_5_695,Wgt_5_696,Wgt_5_697,Wgt_5_698,Wgt_5_699,Wgt_5_700,Wgt_5_701,Wgt_5_702,Wgt_5_703,Wgt_5_704,Wgt_5_705,Wgt_5_706,Wgt_5_707,Wgt_5_708,Wgt_5_709,Wgt_5_710,Wgt_5_711,Wgt_5_712,Wgt_5_713,Wgt_5_714,Wgt_5_715,Wgt_5_716,Wgt_5_717,Wgt_5_718,Wgt_5_719,Wgt_5_720,Wgt_5_721,Wgt_5_722,Wgt_5_723,Wgt_5_724,Wgt_5_725,Wgt_5_726,Wgt_5_727,Wgt_5_728,Wgt_5_729,Wgt_5_730,Wgt_5_731,Wgt_5_732,Wgt_5_733,Wgt_5_734,Wgt_5_735,Wgt_5_736,Wgt_5_737,Wgt_5_738,Wgt_5_739,Wgt_5_740,Wgt_5_741,Wgt_5_742,Wgt_5_743,Wgt_5_744,Wgt_5_745,Wgt_5_746,Wgt_5_747,Wgt_5_748,Wgt_5_749,Wgt_5_750,Wgt_5_751,Wgt_5_752,Wgt_5_753,Wgt_5_754,Wgt_5_755,Wgt_5_756,Wgt_5_757,Wgt_5_758,Wgt_5_759,Wgt_5_760,Wgt_5_761,Wgt_5_762,Wgt_5_763,Wgt_5_764,Wgt_5_765,Wgt_5_766,Wgt_5_767,Wgt_5_768,Wgt_5_769,Wgt_5_770,Wgt_5_771,Wgt_5_772,Wgt_5_773,Wgt_5_774,Wgt_5_775,Wgt_5_776,Wgt_5_777,Wgt_5_778,Wgt_5_779,Wgt_5_780,Wgt_5_781,Wgt_5_782,Wgt_5_783,Wgt_5_784,Wgt_6_0,Wgt_6_1,Wgt_6_2,Wgt_6_3,Wgt_6_4,Wgt_6_5,Wgt_6_6,Wgt_6_7,Wgt_6_8,Wgt_6_9,Wgt_6_10,Wgt_6_11,Wgt_6_12,Wgt_6_13,Wgt_6_14,Wgt_6_15,Wgt_6_16,Wgt_6_17,Wgt_6_18,Wgt_6_19,Wgt_6_20,Wgt_6_21,Wgt_6_22,Wgt_6_23,Wgt_6_24,Wgt_6_25,Wgt_6_26,Wgt_6_27,Wgt_6_28,Wgt_6_29,Wgt_6_30,Wgt_6_31,Wgt_6_32,Wgt_6_33,Wgt_6_34,Wgt_6_35,Wgt_6_36,Wgt_6_37,Wgt_6_38,Wgt_6_39,Wgt_6_40,Wgt_6_41,Wgt_6_42,Wgt_6_43,Wgt_6_44,Wgt_6_45,Wgt_6_46,Wgt_6_47,Wgt_6_48,Wgt_6_49,Wgt_6_50,Wgt_6_51,Wgt_6_52,Wgt_6_53,Wgt_6_54,Wgt_6_55,Wgt_6_56,Wgt_6_57,Wgt_6_58,Wgt_6_59,Wgt_6_60,Wgt_6_61,Wgt_6_62,Wgt_6_63,Wgt_6_64,Wgt_6_65,Wgt_6_66,Wgt_6_67,Wgt_6_68,Wgt_6_69,Wgt_6_70,Wgt_6_71,Wgt_6_72,Wgt_6_73,Wgt_6_74,Wgt_6_75,Wgt_6_76,Wgt_6_77,Wgt_6_78,Wgt_6_79,Wgt_6_80,Wgt_6_81,Wgt_6_82,Wgt_6_83,Wgt_6_84,Wgt_6_85,Wgt_6_86,Wgt_6_87,Wgt_6_88,Wgt_6_89,Wgt_6_90,Wgt_6_91,Wgt_6_92,Wgt_6_93,Wgt_6_94,Wgt_6_95,Wgt_6_96,Wgt_6_97,Wgt_6_98,Wgt_6_99,Wgt_6_100,Wgt_6_101,Wgt_6_102,Wgt_6_103,Wgt_6_104,Wgt_6_105,Wgt_6_106,Wgt_6_107,Wgt_6_108,Wgt_6_109,Wgt_6_110,Wgt_6_111,Wgt_6_112,Wgt_6_113,Wgt_6_114,Wgt_6_115,Wgt_6_116,Wgt_6_117,Wgt_6_118,Wgt_6_119,Wgt_6_120,Wgt_6_121,Wgt_6_122,Wgt_6_123,Wgt_6_124,Wgt_6_125,Wgt_6_126,Wgt_6_127,Wgt_6_128,Wgt_6_129,Wgt_6_130,Wgt_6_131,Wgt_6_132,Wgt_6_133,Wgt_6_134,Wgt_6_135,Wgt_6_136,Wgt_6_137,Wgt_6_138,Wgt_6_139,Wgt_6_140,Wgt_6_141,Wgt_6_142,Wgt_6_143,Wgt_6_144,Wgt_6_145,Wgt_6_146,Wgt_6_147,Wgt_6_148,Wgt_6_149,Wgt_6_150,Wgt_6_151,Wgt_6_152,Wgt_6_153,Wgt_6_154,Wgt_6_155,Wgt_6_156,Wgt_6_157,Wgt_6_158,Wgt_6_159,Wgt_6_160,Wgt_6_161,Wgt_6_162,Wgt_6_163,Wgt_6_164,Wgt_6_165,Wgt_6_166,Wgt_6_167,Wgt_6_168,Wgt_6_169,Wgt_6_170,Wgt_6_171,Wgt_6_172,Wgt_6_173,Wgt_6_174,Wgt_6_175,Wgt_6_176,Wgt_6_177,Wgt_6_178,Wgt_6_179,Wgt_6_180,Wgt_6_181,Wgt_6_182,Wgt_6_183,Wgt_6_184,Wgt_6_185,Wgt_6_186,Wgt_6_187,Wgt_6_188,Wgt_6_189,Wgt_6_190,Wgt_6_191,Wgt_6_192,Wgt_6_193,Wgt_6_194,Wgt_6_195,Wgt_6_196,Wgt_6_197,Wgt_6_198,Wgt_6_199,Wgt_6_200,Wgt_6_201,Wgt_6_202,Wgt_6_203,Wgt_6_204,Wgt_6_205,Wgt_6_206,Wgt_6_207,Wgt_6_208,Wgt_6_209,Wgt_6_210,Wgt_6_211,Wgt_6_212,Wgt_6_213,Wgt_6_214,Wgt_6_215,Wgt_6_216,Wgt_6_217,Wgt_6_218,Wgt_6_219,Wgt_6_220,Wgt_6_221,Wgt_6_222,Wgt_6_223,Wgt_6_224,Wgt_6_225,Wgt_6_226,Wgt_6_227,Wgt_6_228,Wgt_6_229,Wgt_6_230,Wgt_6_231,Wgt_6_232,Wgt_6_233,Wgt_6_234,Wgt_6_235,Wgt_6_236,Wgt_6_237,Wgt_6_238,Wgt_6_239,Wgt_6_240,Wgt_6_241,Wgt_6_242,Wgt_6_243,Wgt_6_244,Wgt_6_245,Wgt_6_246,Wgt_6_247,Wgt_6_248,Wgt_6_249,Wgt_6_250,Wgt_6_251,Wgt_6_252,Wgt_6_253,Wgt_6_254,Wgt_6_255,Wgt_6_256,Wgt_6_257,Wgt_6_258,Wgt_6_259,Wgt_6_260,Wgt_6_261,Wgt_6_262,Wgt_6_263,Wgt_6_264,Wgt_6_265,Wgt_6_266,Wgt_6_267,Wgt_6_268,Wgt_6_269,Wgt_6_270,Wgt_6_271,Wgt_6_272,Wgt_6_273,Wgt_6_274,Wgt_6_275,Wgt_6_276,Wgt_6_277,Wgt_6_278,Wgt_6_279,Wgt_6_280,Wgt_6_281,Wgt_6_282,Wgt_6_283,Wgt_6_284,Wgt_6_285,Wgt_6_286,Wgt_6_287,Wgt_6_288,Wgt_6_289,Wgt_6_290,Wgt_6_291,Wgt_6_292,Wgt_6_293,Wgt_6_294,Wgt_6_295,Wgt_6_296,Wgt_6_297,Wgt_6_298,Wgt_6_299,Wgt_6_300,Wgt_6_301,Wgt_6_302,Wgt_6_303,Wgt_6_304,Wgt_6_305,Wgt_6_306,Wgt_6_307,Wgt_6_308,Wgt_6_309,Wgt_6_310,Wgt_6_311,Wgt_6_312,Wgt_6_313,Wgt_6_314,Wgt_6_315,Wgt_6_316,Wgt_6_317,Wgt_6_318,Wgt_6_319,Wgt_6_320,Wgt_6_321,Wgt_6_322,Wgt_6_323,Wgt_6_324,Wgt_6_325,Wgt_6_326,Wgt_6_327,Wgt_6_328,Wgt_6_329,Wgt_6_330,Wgt_6_331,Wgt_6_332,Wgt_6_333,Wgt_6_334,Wgt_6_335,Wgt_6_336,Wgt_6_337,Wgt_6_338,Wgt_6_339,Wgt_6_340,Wgt_6_341,Wgt_6_342,Wgt_6_343,Wgt_6_344,Wgt_6_345,Wgt_6_346,Wgt_6_347,Wgt_6_348,Wgt_6_349,Wgt_6_350,Wgt_6_351,Wgt_6_352,Wgt_6_353,Wgt_6_354,Wgt_6_355,Wgt_6_356,Wgt_6_357,Wgt_6_358,Wgt_6_359,Wgt_6_360,Wgt_6_361,Wgt_6_362,Wgt_6_363,Wgt_6_364,Wgt_6_365,Wgt_6_366,Wgt_6_367,Wgt_6_368,Wgt_6_369,Wgt_6_370,Wgt_6_371,Wgt_6_372,Wgt_6_373,Wgt_6_374,Wgt_6_375,Wgt_6_376,Wgt_6_377,Wgt_6_378,Wgt_6_379,Wgt_6_380,Wgt_6_381,Wgt_6_382,Wgt_6_383,Wgt_6_384,Wgt_6_385,Wgt_6_386,Wgt_6_387,Wgt_6_388,Wgt_6_389,Wgt_6_390,Wgt_6_391,Wgt_6_392,Wgt_6_393,Wgt_6_394,Wgt_6_395,Wgt_6_396,Wgt_6_397,Wgt_6_398,Wgt_6_399,Wgt_6_400,Wgt_6_401,Wgt_6_402,Wgt_6_403,Wgt_6_404,Wgt_6_405,Wgt_6_406,Wgt_6_407,Wgt_6_408,Wgt_6_409,Wgt_6_410,Wgt_6_411,Wgt_6_412,Wgt_6_413,Wgt_6_414,Wgt_6_415,Wgt_6_416,Wgt_6_417,Wgt_6_418,Wgt_6_419,Wgt_6_420,Wgt_6_421,Wgt_6_422,Wgt_6_423,Wgt_6_424,Wgt_6_425,Wgt_6_426,Wgt_6_427,Wgt_6_428,Wgt_6_429,Wgt_6_430,Wgt_6_431,Wgt_6_432,Wgt_6_433,Wgt_6_434,Wgt_6_435,Wgt_6_436,Wgt_6_437,Wgt_6_438,Wgt_6_439,Wgt_6_440,Wgt_6_441,Wgt_6_442,Wgt_6_443,Wgt_6_444,Wgt_6_445,Wgt_6_446,Wgt_6_447,Wgt_6_448,Wgt_6_449,Wgt_6_450,Wgt_6_451,Wgt_6_452,Wgt_6_453,Wgt_6_454,Wgt_6_455,Wgt_6_456,Wgt_6_457,Wgt_6_458,Wgt_6_459,Wgt_6_460,Wgt_6_461,Wgt_6_462,Wgt_6_463,Wgt_6_464,Wgt_6_465,Wgt_6_466,Wgt_6_467,Wgt_6_468,Wgt_6_469,Wgt_6_470,Wgt_6_471,Wgt_6_472,Wgt_6_473,Wgt_6_474,Wgt_6_475,Wgt_6_476,Wgt_6_477,Wgt_6_478,Wgt_6_479,Wgt_6_480,Wgt_6_481,Wgt_6_482,Wgt_6_483,Wgt_6_484,Wgt_6_485,Wgt_6_486,Wgt_6_487,Wgt_6_488,Wgt_6_489,Wgt_6_490,Wgt_6_491,Wgt_6_492,Wgt_6_493,Wgt_6_494,Wgt_6_495,Wgt_6_496,Wgt_6_497,Wgt_6_498,Wgt_6_499,Wgt_6_500,Wgt_6_501,Wgt_6_502,Wgt_6_503,Wgt_6_504,Wgt_6_505,Wgt_6_506,Wgt_6_507,Wgt_6_508,Wgt_6_509,Wgt_6_510,Wgt_6_511,Wgt_6_512,Wgt_6_513,Wgt_6_514,Wgt_6_515,Wgt_6_516,Wgt_6_517,Wgt_6_518,Wgt_6_519,Wgt_6_520,Wgt_6_521,Wgt_6_522,Wgt_6_523,Wgt_6_524,Wgt_6_525,Wgt_6_526,Wgt_6_527,Wgt_6_528,Wgt_6_529,Wgt_6_530,Wgt_6_531,Wgt_6_532,Wgt_6_533,Wgt_6_534,Wgt_6_535,Wgt_6_536,Wgt_6_537,Wgt_6_538,Wgt_6_539,Wgt_6_540,Wgt_6_541,Wgt_6_542,Wgt_6_543,Wgt_6_544,Wgt_6_545,Wgt_6_546,Wgt_6_547,Wgt_6_548,Wgt_6_549,Wgt_6_550,Wgt_6_551,Wgt_6_552,Wgt_6_553,Wgt_6_554,Wgt_6_555,Wgt_6_556,Wgt_6_557,Wgt_6_558,Wgt_6_559,Wgt_6_560,Wgt_6_561,Wgt_6_562,Wgt_6_563,Wgt_6_564,Wgt_6_565,Wgt_6_566,Wgt_6_567,Wgt_6_568,Wgt_6_569,Wgt_6_570,Wgt_6_571,Wgt_6_572,Wgt_6_573,Wgt_6_574,Wgt_6_575,Wgt_6_576,Wgt_6_577,Wgt_6_578,Wgt_6_579,Wgt_6_580,Wgt_6_581,Wgt_6_582,Wgt_6_583,Wgt_6_584,Wgt_6_585,Wgt_6_586,Wgt_6_587,Wgt_6_588,Wgt_6_589,Wgt_6_590,Wgt_6_591,Wgt_6_592,Wgt_6_593,Wgt_6_594,Wgt_6_595,Wgt_6_596,Wgt_6_597,Wgt_6_598,Wgt_6_599,Wgt_6_600,Wgt_6_601,Wgt_6_602,Wgt_6_603,Wgt_6_604,Wgt_6_605,Wgt_6_606,Wgt_6_607,Wgt_6_608,Wgt_6_609,Wgt_6_610,Wgt_6_611,Wgt_6_612,Wgt_6_613,Wgt_6_614,Wgt_6_615,Wgt_6_616,Wgt_6_617,Wgt_6_618,Wgt_6_619,Wgt_6_620,Wgt_6_621,Wgt_6_622,Wgt_6_623,Wgt_6_624,Wgt_6_625,Wgt_6_626,Wgt_6_627,Wgt_6_628,Wgt_6_629,Wgt_6_630,Wgt_6_631,Wgt_6_632,Wgt_6_633,Wgt_6_634,Wgt_6_635,Wgt_6_636,Wgt_6_637,Wgt_6_638,Wgt_6_639,Wgt_6_640,Wgt_6_641,Wgt_6_642,Wgt_6_643,Wgt_6_644,Wgt_6_645,Wgt_6_646,Wgt_6_647,Wgt_6_648,Wgt_6_649,Wgt_6_650,Wgt_6_651,Wgt_6_652,Wgt_6_653,Wgt_6_654,Wgt_6_655,Wgt_6_656,Wgt_6_657,Wgt_6_658,Wgt_6_659,Wgt_6_660,Wgt_6_661,Wgt_6_662,Wgt_6_663,Wgt_6_664,Wgt_6_665,Wgt_6_666,Wgt_6_667,Wgt_6_668,Wgt_6_669,Wgt_6_670,Wgt_6_671,Wgt_6_672,Wgt_6_673,Wgt_6_674,Wgt_6_675,Wgt_6_676,Wgt_6_677,Wgt_6_678,Wgt_6_679,Wgt_6_680,Wgt_6_681,Wgt_6_682,Wgt_6_683,Wgt_6_684,Wgt_6_685,Wgt_6_686,Wgt_6_687,Wgt_6_688,Wgt_6_689,Wgt_6_690,Wgt_6_691,Wgt_6_692,Wgt_6_693,Wgt_6_694,Wgt_6_695,Wgt_6_696,Wgt_6_697,Wgt_6_698,Wgt_6_699,Wgt_6_700,Wgt_6_701,Wgt_6_702,Wgt_6_703,Wgt_6_704,Wgt_6_705,Wgt_6_706,Wgt_6_707,Wgt_6_708,Wgt_6_709,Wgt_6_710,Wgt_6_711,Wgt_6_712,Wgt_6_713,Wgt_6_714,Wgt_6_715,Wgt_6_716,Wgt_6_717,Wgt_6_718,Wgt_6_719,Wgt_6_720,Wgt_6_721,Wgt_6_722,Wgt_6_723,Wgt_6_724,Wgt_6_725,Wgt_6_726,Wgt_6_727,Wgt_6_728,Wgt_6_729,Wgt_6_730,Wgt_6_731,Wgt_6_732,Wgt_6_733,Wgt_6_734,Wgt_6_735,Wgt_6_736,Wgt_6_737,Wgt_6_738,Wgt_6_739,Wgt_6_740,Wgt_6_741,Wgt_6_742,Wgt_6_743,Wgt_6_744,Wgt_6_745,Wgt_6_746,Wgt_6_747,Wgt_6_748,Wgt_6_749,Wgt_6_750,Wgt_6_751,Wgt_6_752,Wgt_6_753,Wgt_6_754,Wgt_6_755,Wgt_6_756,Wgt_6_757,Wgt_6_758,Wgt_6_759,Wgt_6_760,Wgt_6_761,Wgt_6_762,Wgt_6_763,Wgt_6_764,Wgt_6_765,Wgt_6_766,Wgt_6_767,Wgt_6_768,Wgt_6_769,Wgt_6_770,Wgt_6_771,Wgt_6_772,Wgt_6_773,Wgt_6_774,Wgt_6_775,Wgt_6_776,Wgt_6_777,Wgt_6_778,Wgt_6_779,Wgt_6_780,Wgt_6_781,Wgt_6_782,Wgt_6_783,Wgt_6_784,Wgt_7_0,Wgt_7_1,Wgt_7_2,Wgt_7_3,Wgt_7_4,Wgt_7_5,Wgt_7_6,Wgt_7_7,Wgt_7_8,Wgt_7_9,Wgt_7_10,Wgt_7_11,Wgt_7_12,Wgt_7_13,Wgt_7_14,Wgt_7_15,Wgt_7_16,Wgt_7_17,Wgt_7_18,Wgt_7_19,Wgt_7_20,Wgt_7_21,Wgt_7_22,Wgt_7_23,Wgt_7_24,Wgt_7_25,Wgt_7_26,Wgt_7_27,Wgt_7_28,Wgt_7_29,Wgt_7_30,Wgt_7_31,Wgt_7_32,Wgt_7_33,Wgt_7_34,Wgt_7_35,Wgt_7_36,Wgt_7_37,Wgt_7_38,Wgt_7_39,Wgt_7_40,Wgt_7_41,Wgt_7_42,Wgt_7_43,Wgt_7_44,Wgt_7_45,Wgt_7_46,Wgt_7_47,Wgt_7_48,Wgt_7_49,Wgt_7_50,Wgt_7_51,Wgt_7_52,Wgt_7_53,Wgt_7_54,Wgt_7_55,Wgt_7_56,Wgt_7_57,Wgt_7_58,Wgt_7_59,Wgt_7_60,Wgt_7_61,Wgt_7_62,Wgt_7_63,Wgt_7_64,Wgt_7_65,Wgt_7_66,Wgt_7_67,Wgt_7_68,Wgt_7_69,Wgt_7_70,Wgt_7_71,Wgt_7_72,Wgt_7_73,Wgt_7_74,Wgt_7_75,Wgt_7_76,Wgt_7_77,Wgt_7_78,Wgt_7_79,Wgt_7_80,Wgt_7_81,Wgt_7_82,Wgt_7_83,Wgt_7_84,Wgt_7_85,Wgt_7_86,Wgt_7_87,Wgt_7_88,Wgt_7_89,Wgt_7_90,Wgt_7_91,Wgt_7_92,Wgt_7_93,Wgt_7_94,Wgt_7_95,Wgt_7_96,Wgt_7_97,Wgt_7_98,Wgt_7_99,Wgt_7_100,Wgt_7_101,Wgt_7_102,Wgt_7_103,Wgt_7_104,Wgt_7_105,Wgt_7_106,Wgt_7_107,Wgt_7_108,Wgt_7_109,Wgt_7_110,Wgt_7_111,Wgt_7_112,Wgt_7_113,Wgt_7_114,Wgt_7_115,Wgt_7_116,Wgt_7_117,Wgt_7_118,Wgt_7_119,Wgt_7_120,Wgt_7_121,Wgt_7_122,Wgt_7_123,Wgt_7_124,Wgt_7_125,Wgt_7_126,Wgt_7_127,Wgt_7_128,Wgt_7_129,Wgt_7_130,Wgt_7_131,Wgt_7_132,Wgt_7_133,Wgt_7_134,Wgt_7_135,Wgt_7_136,Wgt_7_137,Wgt_7_138,Wgt_7_139,Wgt_7_140,Wgt_7_141,Wgt_7_142,Wgt_7_143,Wgt_7_144,Wgt_7_145,Wgt_7_146,Wgt_7_147,Wgt_7_148,Wgt_7_149,Wgt_7_150,Wgt_7_151,Wgt_7_152,Wgt_7_153,Wgt_7_154,Wgt_7_155,Wgt_7_156,Wgt_7_157,Wgt_7_158,Wgt_7_159,Wgt_7_160,Wgt_7_161,Wgt_7_162,Wgt_7_163,Wgt_7_164,Wgt_7_165,Wgt_7_166,Wgt_7_167,Wgt_7_168,Wgt_7_169,Wgt_7_170,Wgt_7_171,Wgt_7_172,Wgt_7_173,Wgt_7_174,Wgt_7_175,Wgt_7_176,Wgt_7_177,Wgt_7_178,Wgt_7_179,Wgt_7_180,Wgt_7_181,Wgt_7_182,Wgt_7_183,Wgt_7_184,Wgt_7_185,Wgt_7_186,Wgt_7_187,Wgt_7_188,Wgt_7_189,Wgt_7_190,Wgt_7_191,Wgt_7_192,Wgt_7_193,Wgt_7_194,Wgt_7_195,Wgt_7_196,Wgt_7_197,Wgt_7_198,Wgt_7_199,Wgt_7_200,Wgt_7_201,Wgt_7_202,Wgt_7_203,Wgt_7_204,Wgt_7_205,Wgt_7_206,Wgt_7_207,Wgt_7_208,Wgt_7_209,Wgt_7_210,Wgt_7_211,Wgt_7_212,Wgt_7_213,Wgt_7_214,Wgt_7_215,Wgt_7_216,Wgt_7_217,Wgt_7_218,Wgt_7_219,Wgt_7_220,Wgt_7_221,Wgt_7_222,Wgt_7_223,Wgt_7_224,Wgt_7_225,Wgt_7_226,Wgt_7_227,Wgt_7_228,Wgt_7_229,Wgt_7_230,Wgt_7_231,Wgt_7_232,Wgt_7_233,Wgt_7_234,Wgt_7_235,Wgt_7_236,Wgt_7_237,Wgt_7_238,Wgt_7_239,Wgt_7_240,Wgt_7_241,Wgt_7_242,Wgt_7_243,Wgt_7_244,Wgt_7_245,Wgt_7_246,Wgt_7_247,Wgt_7_248,Wgt_7_249,Wgt_7_250,Wgt_7_251,Wgt_7_252,Wgt_7_253,Wgt_7_254,Wgt_7_255,Wgt_7_256,Wgt_7_257,Wgt_7_258,Wgt_7_259,Wgt_7_260,Wgt_7_261,Wgt_7_262,Wgt_7_263,Wgt_7_264,Wgt_7_265,Wgt_7_266,Wgt_7_267,Wgt_7_268,Wgt_7_269,Wgt_7_270,Wgt_7_271,Wgt_7_272,Wgt_7_273,Wgt_7_274,Wgt_7_275,Wgt_7_276,Wgt_7_277,Wgt_7_278,Wgt_7_279,Wgt_7_280,Wgt_7_281,Wgt_7_282,Wgt_7_283,Wgt_7_284,Wgt_7_285,Wgt_7_286,Wgt_7_287,Wgt_7_288,Wgt_7_289,Wgt_7_290,Wgt_7_291,Wgt_7_292,Wgt_7_293,Wgt_7_294,Wgt_7_295,Wgt_7_296,Wgt_7_297,Wgt_7_298,Wgt_7_299,Wgt_7_300,Wgt_7_301,Wgt_7_302,Wgt_7_303,Wgt_7_304,Wgt_7_305,Wgt_7_306,Wgt_7_307,Wgt_7_308,Wgt_7_309,Wgt_7_310,Wgt_7_311,Wgt_7_312,Wgt_7_313,Wgt_7_314,Wgt_7_315,Wgt_7_316,Wgt_7_317,Wgt_7_318,Wgt_7_319,Wgt_7_320,Wgt_7_321,Wgt_7_322,Wgt_7_323,Wgt_7_324,Wgt_7_325,Wgt_7_326,Wgt_7_327,Wgt_7_328,Wgt_7_329,Wgt_7_330,Wgt_7_331,Wgt_7_332,Wgt_7_333,Wgt_7_334,Wgt_7_335,Wgt_7_336,Wgt_7_337,Wgt_7_338,Wgt_7_339,Wgt_7_340,Wgt_7_341,Wgt_7_342,Wgt_7_343,Wgt_7_344,Wgt_7_345,Wgt_7_346,Wgt_7_347,Wgt_7_348,Wgt_7_349,Wgt_7_350,Wgt_7_351,Wgt_7_352,Wgt_7_353,Wgt_7_354,Wgt_7_355,Wgt_7_356,Wgt_7_357,Wgt_7_358,Wgt_7_359,Wgt_7_360,Wgt_7_361,Wgt_7_362,Wgt_7_363,Wgt_7_364,Wgt_7_365,Wgt_7_366,Wgt_7_367,Wgt_7_368,Wgt_7_369,Wgt_7_370,Wgt_7_371,Wgt_7_372,Wgt_7_373,Wgt_7_374,Wgt_7_375,Wgt_7_376,Wgt_7_377,Wgt_7_378,Wgt_7_379,Wgt_7_380,Wgt_7_381,Wgt_7_382,Wgt_7_383,Wgt_7_384,Wgt_7_385,Wgt_7_386,Wgt_7_387,Wgt_7_388,Wgt_7_389,Wgt_7_390,Wgt_7_391,Wgt_7_392,Wgt_7_393,Wgt_7_394,Wgt_7_395,Wgt_7_396,Wgt_7_397,Wgt_7_398,Wgt_7_399,Wgt_7_400,Wgt_7_401,Wgt_7_402,Wgt_7_403,Wgt_7_404,Wgt_7_405,Wgt_7_406,Wgt_7_407,Wgt_7_408,Wgt_7_409,Wgt_7_410,Wgt_7_411,Wgt_7_412,Wgt_7_413,Wgt_7_414,Wgt_7_415,Wgt_7_416,Wgt_7_417,Wgt_7_418,Wgt_7_419,Wgt_7_420,Wgt_7_421,Wgt_7_422,Wgt_7_423,Wgt_7_424,Wgt_7_425,Wgt_7_426,Wgt_7_427,Wgt_7_428,Wgt_7_429,Wgt_7_430,Wgt_7_431,Wgt_7_432,Wgt_7_433,Wgt_7_434,Wgt_7_435,Wgt_7_436,Wgt_7_437,Wgt_7_438,Wgt_7_439,Wgt_7_440,Wgt_7_441,Wgt_7_442,Wgt_7_443,Wgt_7_444,Wgt_7_445,Wgt_7_446,Wgt_7_447,Wgt_7_448,Wgt_7_449,Wgt_7_450,Wgt_7_451,Wgt_7_452,Wgt_7_453,Wgt_7_454,Wgt_7_455,Wgt_7_456,Wgt_7_457,Wgt_7_458,Wgt_7_459,Wgt_7_460,Wgt_7_461,Wgt_7_462,Wgt_7_463,Wgt_7_464,Wgt_7_465,Wgt_7_466,Wgt_7_467,Wgt_7_468,Wgt_7_469,Wgt_7_470,Wgt_7_471,Wgt_7_472,Wgt_7_473,Wgt_7_474,Wgt_7_475,Wgt_7_476,Wgt_7_477,Wgt_7_478,Wgt_7_479,Wgt_7_480,Wgt_7_481,Wgt_7_482,Wgt_7_483,Wgt_7_484,Wgt_7_485,Wgt_7_486,Wgt_7_487,Wgt_7_488,Wgt_7_489,Wgt_7_490,Wgt_7_491,Wgt_7_492,Wgt_7_493,Wgt_7_494,Wgt_7_495,Wgt_7_496,Wgt_7_497,Wgt_7_498,Wgt_7_499,Wgt_7_500,Wgt_7_501,Wgt_7_502,Wgt_7_503,Wgt_7_504,Wgt_7_505,Wgt_7_506,Wgt_7_507,Wgt_7_508,Wgt_7_509,Wgt_7_510,Wgt_7_511,Wgt_7_512,Wgt_7_513,Wgt_7_514,Wgt_7_515,Wgt_7_516,Wgt_7_517,Wgt_7_518,Wgt_7_519,Wgt_7_520,Wgt_7_521,Wgt_7_522,Wgt_7_523,Wgt_7_524,Wgt_7_525,Wgt_7_526,Wgt_7_527,Wgt_7_528,Wgt_7_529,Wgt_7_530,Wgt_7_531,Wgt_7_532,Wgt_7_533,Wgt_7_534,Wgt_7_535,Wgt_7_536,Wgt_7_537,Wgt_7_538,Wgt_7_539,Wgt_7_540,Wgt_7_541,Wgt_7_542,Wgt_7_543,Wgt_7_544,Wgt_7_545,Wgt_7_546,Wgt_7_547,Wgt_7_548,Wgt_7_549,Wgt_7_550,Wgt_7_551,Wgt_7_552,Wgt_7_553,Wgt_7_554,Wgt_7_555,Wgt_7_556,Wgt_7_557,Wgt_7_558,Wgt_7_559,Wgt_7_560,Wgt_7_561,Wgt_7_562,Wgt_7_563,Wgt_7_564,Wgt_7_565,Wgt_7_566,Wgt_7_567,Wgt_7_568,Wgt_7_569,Wgt_7_570,Wgt_7_571,Wgt_7_572,Wgt_7_573,Wgt_7_574,Wgt_7_575,Wgt_7_576,Wgt_7_577,Wgt_7_578,Wgt_7_579,Wgt_7_580,Wgt_7_581,Wgt_7_582,Wgt_7_583,Wgt_7_584,Wgt_7_585,Wgt_7_586,Wgt_7_587,Wgt_7_588,Wgt_7_589,Wgt_7_590,Wgt_7_591,Wgt_7_592,Wgt_7_593,Wgt_7_594,Wgt_7_595,Wgt_7_596,Wgt_7_597,Wgt_7_598,Wgt_7_599,Wgt_7_600,Wgt_7_601,Wgt_7_602,Wgt_7_603,Wgt_7_604,Wgt_7_605,Wgt_7_606,Wgt_7_607,Wgt_7_608,Wgt_7_609,Wgt_7_610,Wgt_7_611,Wgt_7_612,Wgt_7_613,Wgt_7_614,Wgt_7_615,Wgt_7_616,Wgt_7_617,Wgt_7_618,Wgt_7_619,Wgt_7_620,Wgt_7_621,Wgt_7_622,Wgt_7_623,Wgt_7_624,Wgt_7_625,Wgt_7_626,Wgt_7_627,Wgt_7_628,Wgt_7_629,Wgt_7_630,Wgt_7_631,Wgt_7_632,Wgt_7_633,Wgt_7_634,Wgt_7_635,Wgt_7_636,Wgt_7_637,Wgt_7_638,Wgt_7_639,Wgt_7_640,Wgt_7_641,Wgt_7_642,Wgt_7_643,Wgt_7_644,Wgt_7_645,Wgt_7_646,Wgt_7_647,Wgt_7_648,Wgt_7_649,Wgt_7_650,Wgt_7_651,Wgt_7_652,Wgt_7_653,Wgt_7_654,Wgt_7_655,Wgt_7_656,Wgt_7_657,Wgt_7_658,Wgt_7_659,Wgt_7_660,Wgt_7_661,Wgt_7_662,Wgt_7_663,Wgt_7_664,Wgt_7_665,Wgt_7_666,Wgt_7_667,Wgt_7_668,Wgt_7_669,Wgt_7_670,Wgt_7_671,Wgt_7_672,Wgt_7_673,Wgt_7_674,Wgt_7_675,Wgt_7_676,Wgt_7_677,Wgt_7_678,Wgt_7_679,Wgt_7_680,Wgt_7_681,Wgt_7_682,Wgt_7_683,Wgt_7_684,Wgt_7_685,Wgt_7_686,Wgt_7_687,Wgt_7_688,Wgt_7_689,Wgt_7_690,Wgt_7_691,Wgt_7_692,Wgt_7_693,Wgt_7_694,Wgt_7_695,Wgt_7_696,Wgt_7_697,Wgt_7_698,Wgt_7_699,Wgt_7_700,Wgt_7_701,Wgt_7_702,Wgt_7_703,Wgt_7_704,Wgt_7_705,Wgt_7_706,Wgt_7_707,Wgt_7_708,Wgt_7_709,Wgt_7_710,Wgt_7_711,Wgt_7_712,Wgt_7_713,Wgt_7_714,Wgt_7_715,Wgt_7_716,Wgt_7_717,Wgt_7_718,Wgt_7_719,Wgt_7_720,Wgt_7_721,Wgt_7_722,Wgt_7_723,Wgt_7_724,Wgt_7_725,Wgt_7_726,Wgt_7_727,Wgt_7_728,Wgt_7_729,Wgt_7_730,Wgt_7_731,Wgt_7_732,Wgt_7_733,Wgt_7_734,Wgt_7_735,Wgt_7_736,Wgt_7_737,Wgt_7_738,Wgt_7_739,Wgt_7_740,Wgt_7_741,Wgt_7_742,Wgt_7_743,Wgt_7_744,Wgt_7_745,Wgt_7_746,Wgt_7_747,Wgt_7_748,Wgt_7_749,Wgt_7_750,Wgt_7_751,Wgt_7_752,Wgt_7_753,Wgt_7_754,Wgt_7_755,Wgt_7_756,Wgt_7_757,Wgt_7_758,Wgt_7_759,Wgt_7_760,Wgt_7_761,Wgt_7_762,Wgt_7_763,Wgt_7_764,Wgt_7_765,Wgt_7_766,Wgt_7_767,Wgt_7_768,Wgt_7_769,Wgt_7_770,Wgt_7_771,Wgt_7_772,Wgt_7_773,Wgt_7_774,Wgt_7_775,Wgt_7_776,Wgt_7_777,Wgt_7_778,Wgt_7_779,Wgt_7_780,Wgt_7_781,Wgt_7_782,Wgt_7_783,Wgt_7_784,Wgt_8_0,Wgt_8_1,Wgt_8_2,Wgt_8_3,Wgt_8_4,Wgt_8_5,Wgt_8_6,Wgt_8_7,Wgt_8_8,Wgt_8_9,Wgt_8_10,Wgt_8_11,Wgt_8_12,Wgt_8_13,Wgt_8_14,Wgt_8_15,Wgt_8_16,Wgt_8_17,Wgt_8_18,Wgt_8_19,Wgt_8_20,Wgt_8_21,Wgt_8_22,Wgt_8_23,Wgt_8_24,Wgt_8_25,Wgt_8_26,Wgt_8_27,Wgt_8_28,Wgt_8_29,Wgt_8_30,Wgt_8_31,Wgt_8_32,Wgt_8_33,Wgt_8_34,Wgt_8_35,Wgt_8_36,Wgt_8_37,Wgt_8_38,Wgt_8_39,Wgt_8_40,Wgt_8_41,Wgt_8_42,Wgt_8_43,Wgt_8_44,Wgt_8_45,Wgt_8_46,Wgt_8_47,Wgt_8_48,Wgt_8_49,Wgt_8_50,Wgt_8_51,Wgt_8_52,Wgt_8_53,Wgt_8_54,Wgt_8_55,Wgt_8_56,Wgt_8_57,Wgt_8_58,Wgt_8_59,Wgt_8_60,Wgt_8_61,Wgt_8_62,Wgt_8_63,Wgt_8_64,Wgt_8_65,Wgt_8_66,Wgt_8_67,Wgt_8_68,Wgt_8_69,Wgt_8_70,Wgt_8_71,Wgt_8_72,Wgt_8_73,Wgt_8_74,Wgt_8_75,Wgt_8_76,Wgt_8_77,Wgt_8_78,Wgt_8_79,Wgt_8_80,Wgt_8_81,Wgt_8_82,Wgt_8_83,Wgt_8_84,Wgt_8_85,Wgt_8_86,Wgt_8_87,Wgt_8_88,Wgt_8_89,Wgt_8_90,Wgt_8_91,Wgt_8_92,Wgt_8_93,Wgt_8_94,Wgt_8_95,Wgt_8_96,Wgt_8_97,Wgt_8_98,Wgt_8_99,Wgt_8_100,Wgt_8_101,Wgt_8_102,Wgt_8_103,Wgt_8_104,Wgt_8_105,Wgt_8_106,Wgt_8_107,Wgt_8_108,Wgt_8_109,Wgt_8_110,Wgt_8_111,Wgt_8_112,Wgt_8_113,Wgt_8_114,Wgt_8_115,Wgt_8_116,Wgt_8_117,Wgt_8_118,Wgt_8_119,Wgt_8_120,Wgt_8_121,Wgt_8_122,Wgt_8_123,Wgt_8_124,Wgt_8_125,Wgt_8_126,Wgt_8_127,Wgt_8_128,Wgt_8_129,Wgt_8_130,Wgt_8_131,Wgt_8_132,Wgt_8_133,Wgt_8_134,Wgt_8_135,Wgt_8_136,Wgt_8_137,Wgt_8_138,Wgt_8_139,Wgt_8_140,Wgt_8_141,Wgt_8_142,Wgt_8_143,Wgt_8_144,Wgt_8_145,Wgt_8_146,Wgt_8_147,Wgt_8_148,Wgt_8_149,Wgt_8_150,Wgt_8_151,Wgt_8_152,Wgt_8_153,Wgt_8_154,Wgt_8_155,Wgt_8_156,Wgt_8_157,Wgt_8_158,Wgt_8_159,Wgt_8_160,Wgt_8_161,Wgt_8_162,Wgt_8_163,Wgt_8_164,Wgt_8_165,Wgt_8_166,Wgt_8_167,Wgt_8_168,Wgt_8_169,Wgt_8_170,Wgt_8_171,Wgt_8_172,Wgt_8_173,Wgt_8_174,Wgt_8_175,Wgt_8_176,Wgt_8_177,Wgt_8_178,Wgt_8_179,Wgt_8_180,Wgt_8_181,Wgt_8_182,Wgt_8_183,Wgt_8_184,Wgt_8_185,Wgt_8_186,Wgt_8_187,Wgt_8_188,Wgt_8_189,Wgt_8_190,Wgt_8_191,Wgt_8_192,Wgt_8_193,Wgt_8_194,Wgt_8_195,Wgt_8_196,Wgt_8_197,Wgt_8_198,Wgt_8_199,Wgt_8_200,Wgt_8_201,Wgt_8_202,Wgt_8_203,Wgt_8_204,Wgt_8_205,Wgt_8_206,Wgt_8_207,Wgt_8_208,Wgt_8_209,Wgt_8_210,Wgt_8_211,Wgt_8_212,Wgt_8_213,Wgt_8_214,Wgt_8_215,Wgt_8_216,Wgt_8_217,Wgt_8_218,Wgt_8_219,Wgt_8_220,Wgt_8_221,Wgt_8_222,Wgt_8_223,Wgt_8_224,Wgt_8_225,Wgt_8_226,Wgt_8_227,Wgt_8_228,Wgt_8_229,Wgt_8_230,Wgt_8_231,Wgt_8_232,Wgt_8_233,Wgt_8_234,Wgt_8_235,Wgt_8_236,Wgt_8_237,Wgt_8_238,Wgt_8_239,Wgt_8_240,Wgt_8_241,Wgt_8_242,Wgt_8_243,Wgt_8_244,Wgt_8_245,Wgt_8_246,Wgt_8_247,Wgt_8_248,Wgt_8_249,Wgt_8_250,Wgt_8_251,Wgt_8_252,Wgt_8_253,Wgt_8_254,Wgt_8_255,Wgt_8_256,Wgt_8_257,Wgt_8_258,Wgt_8_259,Wgt_8_260,Wgt_8_261,Wgt_8_262,Wgt_8_263,Wgt_8_264,Wgt_8_265,Wgt_8_266,Wgt_8_267,Wgt_8_268,Wgt_8_269,Wgt_8_270,Wgt_8_271,Wgt_8_272,Wgt_8_273,Wgt_8_274,Wgt_8_275,Wgt_8_276,Wgt_8_277,Wgt_8_278,Wgt_8_279,Wgt_8_280,Wgt_8_281,Wgt_8_282,Wgt_8_283,Wgt_8_284,Wgt_8_285,Wgt_8_286,Wgt_8_287,Wgt_8_288,Wgt_8_289,Wgt_8_290,Wgt_8_291,Wgt_8_292,Wgt_8_293,Wgt_8_294,Wgt_8_295,Wgt_8_296,Wgt_8_297,Wgt_8_298,Wgt_8_299,Wgt_8_300,Wgt_8_301,Wgt_8_302,Wgt_8_303,Wgt_8_304,Wgt_8_305,Wgt_8_306,Wgt_8_307,Wgt_8_308,Wgt_8_309,Wgt_8_310,Wgt_8_311,Wgt_8_312,Wgt_8_313,Wgt_8_314,Wgt_8_315,Wgt_8_316,Wgt_8_317,Wgt_8_318,Wgt_8_319,Wgt_8_320,Wgt_8_321,Wgt_8_322,Wgt_8_323,Wgt_8_324,Wgt_8_325,Wgt_8_326,Wgt_8_327,Wgt_8_328,Wgt_8_329,Wgt_8_330,Wgt_8_331,Wgt_8_332,Wgt_8_333,Wgt_8_334,Wgt_8_335,Wgt_8_336,Wgt_8_337,Wgt_8_338,Wgt_8_339,Wgt_8_340,Wgt_8_341,Wgt_8_342,Wgt_8_343,Wgt_8_344,Wgt_8_345,Wgt_8_346,Wgt_8_347,Wgt_8_348,Wgt_8_349,Wgt_8_350,Wgt_8_351,Wgt_8_352,Wgt_8_353,Wgt_8_354,Wgt_8_355,Wgt_8_356,Wgt_8_357,Wgt_8_358,Wgt_8_359,Wgt_8_360,Wgt_8_361,Wgt_8_362,Wgt_8_363,Wgt_8_364,Wgt_8_365,Wgt_8_366,Wgt_8_367,Wgt_8_368,Wgt_8_369,Wgt_8_370,Wgt_8_371,Wgt_8_372,Wgt_8_373,Wgt_8_374,Wgt_8_375,Wgt_8_376,Wgt_8_377,Wgt_8_378,Wgt_8_379,Wgt_8_380,Wgt_8_381,Wgt_8_382,Wgt_8_383,Wgt_8_384,Wgt_8_385,Wgt_8_386,Wgt_8_387,Wgt_8_388,Wgt_8_389,Wgt_8_390,Wgt_8_391,Wgt_8_392,Wgt_8_393,Wgt_8_394,Wgt_8_395,Wgt_8_396,Wgt_8_397,Wgt_8_398,Wgt_8_399,Wgt_8_400,Wgt_8_401,Wgt_8_402,Wgt_8_403,Wgt_8_404,Wgt_8_405,Wgt_8_406,Wgt_8_407,Wgt_8_408,Wgt_8_409,Wgt_8_410,Wgt_8_411,Wgt_8_412,Wgt_8_413,Wgt_8_414,Wgt_8_415,Wgt_8_416,Wgt_8_417,Wgt_8_418,Wgt_8_419,Wgt_8_420,Wgt_8_421,Wgt_8_422,Wgt_8_423,Wgt_8_424,Wgt_8_425,Wgt_8_426,Wgt_8_427,Wgt_8_428,Wgt_8_429,Wgt_8_430,Wgt_8_431,Wgt_8_432,Wgt_8_433,Wgt_8_434,Wgt_8_435,Wgt_8_436,Wgt_8_437,Wgt_8_438,Wgt_8_439,Wgt_8_440,Wgt_8_441,Wgt_8_442,Wgt_8_443,Wgt_8_444,Wgt_8_445,Wgt_8_446,Wgt_8_447,Wgt_8_448,Wgt_8_449,Wgt_8_450,Wgt_8_451,Wgt_8_452,Wgt_8_453,Wgt_8_454,Wgt_8_455,Wgt_8_456,Wgt_8_457,Wgt_8_458,Wgt_8_459,Wgt_8_460,Wgt_8_461,Wgt_8_462,Wgt_8_463,Wgt_8_464,Wgt_8_465,Wgt_8_466,Wgt_8_467,Wgt_8_468,Wgt_8_469,Wgt_8_470,Wgt_8_471,Wgt_8_472,Wgt_8_473,Wgt_8_474,Wgt_8_475,Wgt_8_476,Wgt_8_477,Wgt_8_478,Wgt_8_479,Wgt_8_480,Wgt_8_481,Wgt_8_482,Wgt_8_483,Wgt_8_484,Wgt_8_485,Wgt_8_486,Wgt_8_487,Wgt_8_488,Wgt_8_489,Wgt_8_490,Wgt_8_491,Wgt_8_492,Wgt_8_493,Wgt_8_494,Wgt_8_495,Wgt_8_496,Wgt_8_497,Wgt_8_498,Wgt_8_499,Wgt_8_500,Wgt_8_501,Wgt_8_502,Wgt_8_503,Wgt_8_504,Wgt_8_505,Wgt_8_506,Wgt_8_507,Wgt_8_508,Wgt_8_509,Wgt_8_510,Wgt_8_511,Wgt_8_512,Wgt_8_513,Wgt_8_514,Wgt_8_515,Wgt_8_516,Wgt_8_517,Wgt_8_518,Wgt_8_519,Wgt_8_520,Wgt_8_521,Wgt_8_522,Wgt_8_523,Wgt_8_524,Wgt_8_525,Wgt_8_526,Wgt_8_527,Wgt_8_528,Wgt_8_529,Wgt_8_530,Wgt_8_531,Wgt_8_532,Wgt_8_533,Wgt_8_534,Wgt_8_535,Wgt_8_536,Wgt_8_537,Wgt_8_538,Wgt_8_539,Wgt_8_540,Wgt_8_541,Wgt_8_542,Wgt_8_543,Wgt_8_544,Wgt_8_545,Wgt_8_546,Wgt_8_547,Wgt_8_548,Wgt_8_549,Wgt_8_550,Wgt_8_551,Wgt_8_552,Wgt_8_553,Wgt_8_554,Wgt_8_555,Wgt_8_556,Wgt_8_557,Wgt_8_558,Wgt_8_559,Wgt_8_560,Wgt_8_561,Wgt_8_562,Wgt_8_563,Wgt_8_564,Wgt_8_565,Wgt_8_566,Wgt_8_567,Wgt_8_568,Wgt_8_569,Wgt_8_570,Wgt_8_571,Wgt_8_572,Wgt_8_573,Wgt_8_574,Wgt_8_575,Wgt_8_576,Wgt_8_577,Wgt_8_578,Wgt_8_579,Wgt_8_580,Wgt_8_581,Wgt_8_582,Wgt_8_583,Wgt_8_584,Wgt_8_585,Wgt_8_586,Wgt_8_587,Wgt_8_588,Wgt_8_589,Wgt_8_590,Wgt_8_591,Wgt_8_592,Wgt_8_593,Wgt_8_594,Wgt_8_595,Wgt_8_596,Wgt_8_597,Wgt_8_598,Wgt_8_599,Wgt_8_600,Wgt_8_601,Wgt_8_602,Wgt_8_603,Wgt_8_604,Wgt_8_605,Wgt_8_606,Wgt_8_607,Wgt_8_608,Wgt_8_609,Wgt_8_610,Wgt_8_611,Wgt_8_612,Wgt_8_613,Wgt_8_614,Wgt_8_615,Wgt_8_616,Wgt_8_617,Wgt_8_618,Wgt_8_619,Wgt_8_620,Wgt_8_621,Wgt_8_622,Wgt_8_623,Wgt_8_624,Wgt_8_625,Wgt_8_626,Wgt_8_627,Wgt_8_628,Wgt_8_629,Wgt_8_630,Wgt_8_631,Wgt_8_632,Wgt_8_633,Wgt_8_634,Wgt_8_635,Wgt_8_636,Wgt_8_637,Wgt_8_638,Wgt_8_639,Wgt_8_640,Wgt_8_641,Wgt_8_642,Wgt_8_643,Wgt_8_644,Wgt_8_645,Wgt_8_646,Wgt_8_647,Wgt_8_648,Wgt_8_649,Wgt_8_650,Wgt_8_651,Wgt_8_652,Wgt_8_653,Wgt_8_654,Wgt_8_655,Wgt_8_656,Wgt_8_657,Wgt_8_658,Wgt_8_659,Wgt_8_660,Wgt_8_661,Wgt_8_662,Wgt_8_663,Wgt_8_664,Wgt_8_665,Wgt_8_666,Wgt_8_667,Wgt_8_668,Wgt_8_669,Wgt_8_670,Wgt_8_671,Wgt_8_672,Wgt_8_673,Wgt_8_674,Wgt_8_675,Wgt_8_676,Wgt_8_677,Wgt_8_678,Wgt_8_679,Wgt_8_680,Wgt_8_681,Wgt_8_682,Wgt_8_683,Wgt_8_684,Wgt_8_685,Wgt_8_686,Wgt_8_687,Wgt_8_688,Wgt_8_689,Wgt_8_690,Wgt_8_691,Wgt_8_692,Wgt_8_693,Wgt_8_694,Wgt_8_695,Wgt_8_696,Wgt_8_697,Wgt_8_698,Wgt_8_699,Wgt_8_700,Wgt_8_701,Wgt_8_702,Wgt_8_703,Wgt_8_704,Wgt_8_705,Wgt_8_706,Wgt_8_707,Wgt_8_708,Wgt_8_709,Wgt_8_710,Wgt_8_711,Wgt_8_712,Wgt_8_713,Wgt_8_714,Wgt_8_715,Wgt_8_716,Wgt_8_717,Wgt_8_718,Wgt_8_719,Wgt_8_720,Wgt_8_721,Wgt_8_722,Wgt_8_723,Wgt_8_724,Wgt_8_725,Wgt_8_726,Wgt_8_727,Wgt_8_728,Wgt_8_729,Wgt_8_730,Wgt_8_731,Wgt_8_732,Wgt_8_733,Wgt_8_734,Wgt_8_735,Wgt_8_736,Wgt_8_737,Wgt_8_738,Wgt_8_739,Wgt_8_740,Wgt_8_741,Wgt_8_742,Wgt_8_743,Wgt_8_744,Wgt_8_745,Wgt_8_746,Wgt_8_747,Wgt_8_748,Wgt_8_749,Wgt_8_750,Wgt_8_751,Wgt_8_752,Wgt_8_753,Wgt_8_754,Wgt_8_755,Wgt_8_756,Wgt_8_757,Wgt_8_758,Wgt_8_759,Wgt_8_760,Wgt_8_761,Wgt_8_762,Wgt_8_763,Wgt_8_764,Wgt_8_765,Wgt_8_766,Wgt_8_767,Wgt_8_768,Wgt_8_769,Wgt_8_770,Wgt_8_771,Wgt_8_772,Wgt_8_773,Wgt_8_774,Wgt_8_775,Wgt_8_776,Wgt_8_777,Wgt_8_778,Wgt_8_779,Wgt_8_780,Wgt_8_781,Wgt_8_782,Wgt_8_783,Wgt_8_784,Wgt_9_0,Wgt_9_1,Wgt_9_2,Wgt_9_3,Wgt_9_4,Wgt_9_5,Wgt_9_6,Wgt_9_7,Wgt_9_8,Wgt_9_9,Wgt_9_10,Wgt_9_11,Wgt_9_12,Wgt_9_13,Wgt_9_14,Wgt_9_15,Wgt_9_16,Wgt_9_17,Wgt_9_18,Wgt_9_19,Wgt_9_20,Wgt_9_21,Wgt_9_22,Wgt_9_23,Wgt_9_24,Wgt_9_25,Wgt_9_26,Wgt_9_27,Wgt_9_28,Wgt_9_29,Wgt_9_30,Wgt_9_31,Wgt_9_32,Wgt_9_33,Wgt_9_34,Wgt_9_35,Wgt_9_36,Wgt_9_37,Wgt_9_38,Wgt_9_39,Wgt_9_40,Wgt_9_41,Wgt_9_42,Wgt_9_43,Wgt_9_44,Wgt_9_45,Wgt_9_46,Wgt_9_47,Wgt_9_48,Wgt_9_49,Wgt_9_50,Wgt_9_51,Wgt_9_52,Wgt_9_53,Wgt_9_54,Wgt_9_55,Wgt_9_56,Wgt_9_57,Wgt_9_58,Wgt_9_59,Wgt_9_60,Wgt_9_61,Wgt_9_62,Wgt_9_63,Wgt_9_64,Wgt_9_65,Wgt_9_66,Wgt_9_67,Wgt_9_68,Wgt_9_69,Wgt_9_70,Wgt_9_71,Wgt_9_72,Wgt_9_73,Wgt_9_74,Wgt_9_75,Wgt_9_76,Wgt_9_77,Wgt_9_78,Wgt_9_79,Wgt_9_80,Wgt_9_81,Wgt_9_82,Wgt_9_83,Wgt_9_84,Wgt_9_85,Wgt_9_86,Wgt_9_87,Wgt_9_88,Wgt_9_89,Wgt_9_90,Wgt_9_91,Wgt_9_92,Wgt_9_93,Wgt_9_94,Wgt_9_95,Wgt_9_96,Wgt_9_97,Wgt_9_98,Wgt_9_99,Wgt_9_100,Wgt_9_101,Wgt_9_102,Wgt_9_103,Wgt_9_104,Wgt_9_105,Wgt_9_106,Wgt_9_107,Wgt_9_108,Wgt_9_109,Wgt_9_110,Wgt_9_111,Wgt_9_112,Wgt_9_113,Wgt_9_114,Wgt_9_115,Wgt_9_116,Wgt_9_117,Wgt_9_118,Wgt_9_119,Wgt_9_120,Wgt_9_121,Wgt_9_122,Wgt_9_123,Wgt_9_124,Wgt_9_125,Wgt_9_126,Wgt_9_127,Wgt_9_128,Wgt_9_129,Wgt_9_130,Wgt_9_131,Wgt_9_132,Wgt_9_133,Wgt_9_134,Wgt_9_135,Wgt_9_136,Wgt_9_137,Wgt_9_138,Wgt_9_139,Wgt_9_140,Wgt_9_141,Wgt_9_142,Wgt_9_143,Wgt_9_144,Wgt_9_145,Wgt_9_146,Wgt_9_147,Wgt_9_148,Wgt_9_149,Wgt_9_150,Wgt_9_151,Wgt_9_152,Wgt_9_153,Wgt_9_154,Wgt_9_155,Wgt_9_156,Wgt_9_157,Wgt_9_158,Wgt_9_159,Wgt_9_160,Wgt_9_161,Wgt_9_162,Wgt_9_163,Wgt_9_164,Wgt_9_165,Wgt_9_166,Wgt_9_167,Wgt_9_168,Wgt_9_169,Wgt_9_170,Wgt_9_171,Wgt_9_172,Wgt_9_173,Wgt_9_174,Wgt_9_175,Wgt_9_176,Wgt_9_177,Wgt_9_178,Wgt_9_179,Wgt_9_180,Wgt_9_181,Wgt_9_182,Wgt_9_183,Wgt_9_184,Wgt_9_185,Wgt_9_186,Wgt_9_187,Wgt_9_188,Wgt_9_189,Wgt_9_190,Wgt_9_191,Wgt_9_192,Wgt_9_193,Wgt_9_194,Wgt_9_195,Wgt_9_196,Wgt_9_197,Wgt_9_198,Wgt_9_199,Wgt_9_200,Wgt_9_201,Wgt_9_202,Wgt_9_203,Wgt_9_204,Wgt_9_205,Wgt_9_206,Wgt_9_207,Wgt_9_208,Wgt_9_209,Wgt_9_210,Wgt_9_211,Wgt_9_212,Wgt_9_213,Wgt_9_214,Wgt_9_215,Wgt_9_216,Wgt_9_217,Wgt_9_218,Wgt_9_219,Wgt_9_220,Wgt_9_221,Wgt_9_222,Wgt_9_223,Wgt_9_224,Wgt_9_225,Wgt_9_226,Wgt_9_227,Wgt_9_228,Wgt_9_229,Wgt_9_230,Wgt_9_231,Wgt_9_232,Wgt_9_233,Wgt_9_234,Wgt_9_235,Wgt_9_236,Wgt_9_237,Wgt_9_238,Wgt_9_239,Wgt_9_240,Wgt_9_241,Wgt_9_242,Wgt_9_243,Wgt_9_244,Wgt_9_245,Wgt_9_246,Wgt_9_247,Wgt_9_248,Wgt_9_249,Wgt_9_250,Wgt_9_251,Wgt_9_252,Wgt_9_253,Wgt_9_254,Wgt_9_255,Wgt_9_256,Wgt_9_257,Wgt_9_258,Wgt_9_259,Wgt_9_260,Wgt_9_261,Wgt_9_262,Wgt_9_263,Wgt_9_264,Wgt_9_265,Wgt_9_266,Wgt_9_267,Wgt_9_268,Wgt_9_269,Wgt_9_270,Wgt_9_271,Wgt_9_272,Wgt_9_273,Wgt_9_274,Wgt_9_275,Wgt_9_276,Wgt_9_277,Wgt_9_278,Wgt_9_279,Wgt_9_280,Wgt_9_281,Wgt_9_282,Wgt_9_283,Wgt_9_284,Wgt_9_285,Wgt_9_286,Wgt_9_287,Wgt_9_288,Wgt_9_289,Wgt_9_290,Wgt_9_291,Wgt_9_292,Wgt_9_293,Wgt_9_294,Wgt_9_295,Wgt_9_296,Wgt_9_297,Wgt_9_298,Wgt_9_299,Wgt_9_300,Wgt_9_301,Wgt_9_302,Wgt_9_303,Wgt_9_304,Wgt_9_305,Wgt_9_306,Wgt_9_307,Wgt_9_308,Wgt_9_309,Wgt_9_310,Wgt_9_311,Wgt_9_312,Wgt_9_313,Wgt_9_314,Wgt_9_315,Wgt_9_316,Wgt_9_317,Wgt_9_318,Wgt_9_319,Wgt_9_320,Wgt_9_321,Wgt_9_322,Wgt_9_323,Wgt_9_324,Wgt_9_325,Wgt_9_326,Wgt_9_327,Wgt_9_328,Wgt_9_329,Wgt_9_330,Wgt_9_331,Wgt_9_332,Wgt_9_333,Wgt_9_334,Wgt_9_335,Wgt_9_336,Wgt_9_337,Wgt_9_338,Wgt_9_339,Wgt_9_340,Wgt_9_341,Wgt_9_342,Wgt_9_343,Wgt_9_344,Wgt_9_345,Wgt_9_346,Wgt_9_347,Wgt_9_348,Wgt_9_349,Wgt_9_350,Wgt_9_351,Wgt_9_352,Wgt_9_353,Wgt_9_354,Wgt_9_355,Wgt_9_356,Wgt_9_357,Wgt_9_358,Wgt_9_359,Wgt_9_360,Wgt_9_361,Wgt_9_362,Wgt_9_363,Wgt_9_364,Wgt_9_365,Wgt_9_366,Wgt_9_367,Wgt_9_368,Wgt_9_369,Wgt_9_370,Wgt_9_371,Wgt_9_372,Wgt_9_373,Wgt_9_374,Wgt_9_375,Wgt_9_376,Wgt_9_377,Wgt_9_378,Wgt_9_379,Wgt_9_380,Wgt_9_381,Wgt_9_382,Wgt_9_383,Wgt_9_384,Wgt_9_385,Wgt_9_386,Wgt_9_387,Wgt_9_388,Wgt_9_389,Wgt_9_390,Wgt_9_391,Wgt_9_392,Wgt_9_393,Wgt_9_394,Wgt_9_395,Wgt_9_396,Wgt_9_397,Wgt_9_398,Wgt_9_399,Wgt_9_400,Wgt_9_401,Wgt_9_402,Wgt_9_403,Wgt_9_404,Wgt_9_405,Wgt_9_406,Wgt_9_407,Wgt_9_408,Wgt_9_409,Wgt_9_410,Wgt_9_411,Wgt_9_412,Wgt_9_413,Wgt_9_414,Wgt_9_415,Wgt_9_416,Wgt_9_417,Wgt_9_418,Wgt_9_419,Wgt_9_420,Wgt_9_421,Wgt_9_422,Wgt_9_423,Wgt_9_424,Wgt_9_425,Wgt_9_426,Wgt_9_427,Wgt_9_428,Wgt_9_429,Wgt_9_430,Wgt_9_431,Wgt_9_432,Wgt_9_433,Wgt_9_434,Wgt_9_435,Wgt_9_436,Wgt_9_437,Wgt_9_438,Wgt_9_439,Wgt_9_440,Wgt_9_441,Wgt_9_442,Wgt_9_443,Wgt_9_444,Wgt_9_445,Wgt_9_446,Wgt_9_447,Wgt_9_448,Wgt_9_449,Wgt_9_450,Wgt_9_451,Wgt_9_452,Wgt_9_453,Wgt_9_454,Wgt_9_455,Wgt_9_456,Wgt_9_457,Wgt_9_458,Wgt_9_459,Wgt_9_460,Wgt_9_461,Wgt_9_462,Wgt_9_463,Wgt_9_464,Wgt_9_465,Wgt_9_466,Wgt_9_467,Wgt_9_468,Wgt_9_469,Wgt_9_470,Wgt_9_471,Wgt_9_472,Wgt_9_473,Wgt_9_474,Wgt_9_475,Wgt_9_476,Wgt_9_477,Wgt_9_478,Wgt_9_479,Wgt_9_480,Wgt_9_481,Wgt_9_482,Wgt_9_483,Wgt_9_484,Wgt_9_485,Wgt_9_486,Wgt_9_487,Wgt_9_488,Wgt_9_489,Wgt_9_490,Wgt_9_491,Wgt_9_492,Wgt_9_493,Wgt_9_494,Wgt_9_495,Wgt_9_496,Wgt_9_497,Wgt_9_498,Wgt_9_499,Wgt_9_500,Wgt_9_501,Wgt_9_502,Wgt_9_503,Wgt_9_504,Wgt_9_505,Wgt_9_506,Wgt_9_507,Wgt_9_508,Wgt_9_509,Wgt_9_510,Wgt_9_511,Wgt_9_512,Wgt_9_513,Wgt_9_514,Wgt_9_515,Wgt_9_516,Wgt_9_517,Wgt_9_518,Wgt_9_519,Wgt_9_520,Wgt_9_521,Wgt_9_522,Wgt_9_523,Wgt_9_524,Wgt_9_525,Wgt_9_526,Wgt_9_527,Wgt_9_528,Wgt_9_529,Wgt_9_530,Wgt_9_531,Wgt_9_532,Wgt_9_533,Wgt_9_534,Wgt_9_535,Wgt_9_536,Wgt_9_537,Wgt_9_538,Wgt_9_539,Wgt_9_540,Wgt_9_541,Wgt_9_542,Wgt_9_543,Wgt_9_544,Wgt_9_545,Wgt_9_546,Wgt_9_547,Wgt_9_548,Wgt_9_549,Wgt_9_550,Wgt_9_551,Wgt_9_552,Wgt_9_553,Wgt_9_554,Wgt_9_555,Wgt_9_556,Wgt_9_557,Wgt_9_558,Wgt_9_559,Wgt_9_560,Wgt_9_561,Wgt_9_562,Wgt_9_563,Wgt_9_564,Wgt_9_565,Wgt_9_566,Wgt_9_567,Wgt_9_568,Wgt_9_569,Wgt_9_570,Wgt_9_571,Wgt_9_572,Wgt_9_573,Wgt_9_574,Wgt_9_575,Wgt_9_576,Wgt_9_577,Wgt_9_578,Wgt_9_579,Wgt_9_580,Wgt_9_581,Wgt_9_582,Wgt_9_583,Wgt_9_584,Wgt_9_585,Wgt_9_586,Wgt_9_587,Wgt_9_588,Wgt_9_589,Wgt_9_590,Wgt_9_591,Wgt_9_592,Wgt_9_593,Wgt_9_594,Wgt_9_595,Wgt_9_596,Wgt_9_597,Wgt_9_598,Wgt_9_599,Wgt_9_600,Wgt_9_601,Wgt_9_602,Wgt_9_603,Wgt_9_604,Wgt_9_605,Wgt_9_606,Wgt_9_607,Wgt_9_608,Wgt_9_609,Wgt_9_610,Wgt_9_611,Wgt_9_612,Wgt_9_613,Wgt_9_614,Wgt_9_615,Wgt_9_616,Wgt_9_617,Wgt_9_618,Wgt_9_619,Wgt_9_620,Wgt_9_621,Wgt_9_622,Wgt_9_623,Wgt_9_624,Wgt_9_625,Wgt_9_626,Wgt_9_627,Wgt_9_628,Wgt_9_629,Wgt_9_630,Wgt_9_631,Wgt_9_632,Wgt_9_633,Wgt_9_634,Wgt_9_635,Wgt_9_636,Wgt_9_637,Wgt_9_638,Wgt_9_639,Wgt_9_640,Wgt_9_641,Wgt_9_642,Wgt_9_643,Wgt_9_644,Wgt_9_645,Wgt_9_646,Wgt_9_647,Wgt_9_648,Wgt_9_649,Wgt_9_650,Wgt_9_651,Wgt_9_652,Wgt_9_653,Wgt_9_654,Wgt_9_655,Wgt_9_656,Wgt_9_657,Wgt_9_658,Wgt_9_659,Wgt_9_660,Wgt_9_661,Wgt_9_662,Wgt_9_663,Wgt_9_664,Wgt_9_665,Wgt_9_666,Wgt_9_667,Wgt_9_668,Wgt_9_669,Wgt_9_670,Wgt_9_671,Wgt_9_672,Wgt_9_673,Wgt_9_674,Wgt_9_675,Wgt_9_676,Wgt_9_677,Wgt_9_678,Wgt_9_679,Wgt_9_680,Wgt_9_681,Wgt_9_682,Wgt_9_683,Wgt_9_684,Wgt_9_685,Wgt_9_686,Wgt_9_687,Wgt_9_688,Wgt_9_689,Wgt_9_690,Wgt_9_691,Wgt_9_692,Wgt_9_693,Wgt_9_694,Wgt_9_695,Wgt_9_696,Wgt_9_697,Wgt_9_698,Wgt_9_699,Wgt_9_700,Wgt_9_701,Wgt_9_702,Wgt_9_703,Wgt_9_704,Wgt_9_705,Wgt_9_706,Wgt_9_707,Wgt_9_708,Wgt_9_709,Wgt_9_710,Wgt_9_711,Wgt_9_712,Wgt_9_713,Wgt_9_714,Wgt_9_715,Wgt_9_716,Wgt_9_717,Wgt_9_718,Wgt_9_719,Wgt_9_720,Wgt_9_721,Wgt_9_722,Wgt_9_723,Wgt_9_724,Wgt_9_725,Wgt_9_726,Wgt_9_727,Wgt_9_728,Wgt_9_729,Wgt_9_730,Wgt_9_731,Wgt_9_732,Wgt_9_733,Wgt_9_734,Wgt_9_735,Wgt_9_736,Wgt_9_737,Wgt_9_738,Wgt_9_739,Wgt_9_740,Wgt_9_741,Wgt_9_742,Wgt_9_743,Wgt_9_744,Wgt_9_745,Wgt_9_746,Wgt_9_747,Wgt_9_748,Wgt_9_749,Wgt_9_750,Wgt_9_751,Wgt_9_752,Wgt_9_753,Wgt_9_754,Wgt_9_755,Wgt_9_756,Wgt_9_757,Wgt_9_758,Wgt_9_759,Wgt_9_760,Wgt_9_761,Wgt_9_762,Wgt_9_763,Wgt_9_764,Wgt_9_765,Wgt_9_766,Wgt_9_767,Wgt_9_768,Wgt_9_769,Wgt_9_770,Wgt_9_771,Wgt_9_772,Wgt_9_773,Wgt_9_774,Wgt_9_775,Wgt_9_776,Wgt_9_777,Wgt_9_778,Wgt_9_779,Wgt_9_780,Wgt_9_781,Wgt_9_782,Wgt_9_783,Wgt_9_784,
	Pix_0,Pix_1,Pix_2,Pix_3,Pix_4,Pix_5,Pix_6,Pix_7,Pix_8,Pix_9,Pix_10,Pix_11,Pix_12,Pix_13,Pix_14,Pix_15,Pix_16,Pix_17,Pix_18,Pix_19,Pix_20,Pix_21,Pix_22,Pix_23,Pix_24,Pix_25,Pix_26,Pix_27,Pix_28,Pix_29,Pix_30,Pix_31,Pix_32,Pix_33,Pix_34,Pix_35,Pix_36,Pix_37,Pix_38,Pix_39,Pix_40,Pix_41,Pix_42,Pix_43,Pix_44,Pix_45,Pix_46,Pix_47,Pix_48,Pix_49,Pix_50,Pix_51,Pix_52,Pix_53,Pix_54,Pix_55,Pix_56,Pix_57,Pix_58,Pix_59,Pix_60,Pix_61,Pix_62,Pix_63,Pix_64,Pix_65,Pix_66,Pix_67,Pix_68,Pix_69,Pix_70,Pix_71,Pix_72,Pix_73,Pix_74,Pix_75,Pix_76,Pix_77,Pix_78,Pix_79,Pix_80,Pix_81,Pix_82,Pix_83,Pix_84,Pix_85,Pix_86,Pix_87,Pix_88,Pix_89,Pix_90,Pix_91,Pix_92,Pix_93,Pix_94,Pix_95,Pix_96,Pix_97,Pix_98,Pix_99,Pix_100,Pix_101,Pix_102,Pix_103,Pix_104,Pix_105,Pix_106,Pix_107,Pix_108,Pix_109,Pix_110,Pix_111,Pix_112,Pix_113,Pix_114,Pix_115,Pix_116,Pix_117,Pix_118,Pix_119,Pix_120,Pix_121,Pix_122,Pix_123,Pix_124,Pix_125,Pix_126,Pix_127,Pix_128,Pix_129,Pix_130,Pix_131,Pix_132,Pix_133,Pix_134,Pix_135,Pix_136,Pix_137,Pix_138,Pix_139,Pix_140,Pix_141,Pix_142,Pix_143,Pix_144,Pix_145,Pix_146,Pix_147,Pix_148,Pix_149,Pix_150,Pix_151,Pix_152,Pix_153,Pix_154,Pix_155,Pix_156,Pix_157,Pix_158,Pix_159,Pix_160,Pix_161,Pix_162,Pix_163,Pix_164,Pix_165,Pix_166,Pix_167,Pix_168,Pix_169,Pix_170,Pix_171,Pix_172,Pix_173,Pix_174,Pix_175,Pix_176,Pix_177,Pix_178,Pix_179,Pix_180,Pix_181,Pix_182,Pix_183,Pix_184,Pix_185,Pix_186,Pix_187,Pix_188,Pix_189,Pix_190,Pix_191,Pix_192,Pix_193,Pix_194,Pix_195,Pix_196,Pix_197,Pix_198,Pix_199,Pix_200,Pix_201,Pix_202,Pix_203,Pix_204,Pix_205,Pix_206,Pix_207,Pix_208,Pix_209,Pix_210,Pix_211,Pix_212,Pix_213,Pix_214,Pix_215,Pix_216,Pix_217,Pix_218,Pix_219,Pix_220,Pix_221,Pix_222,Pix_223,Pix_224,Pix_225,Pix_226,Pix_227,Pix_228,Pix_229,Pix_230,Pix_231,Pix_232,Pix_233,Pix_234,Pix_235,Pix_236,Pix_237,Pix_238,Pix_239,Pix_240,Pix_241,Pix_242,Pix_243,Pix_244,Pix_245,Pix_246,Pix_247,Pix_248,Pix_249,Pix_250,Pix_251,Pix_252,Pix_253,Pix_254,Pix_255,Pix_256,Pix_257,Pix_258,Pix_259,Pix_260,Pix_261,Pix_262,Pix_263,Pix_264,Pix_265,Pix_266,Pix_267,Pix_268,Pix_269,Pix_270,Pix_271,Pix_272,Pix_273,Pix_274,Pix_275,Pix_276,Pix_277,Pix_278,Pix_279,Pix_280,Pix_281,Pix_282,Pix_283,Pix_284,Pix_285,Pix_286,Pix_287,Pix_288,Pix_289,Pix_290,Pix_291,Pix_292,Pix_293,Pix_294,Pix_295,Pix_296,Pix_297,Pix_298,Pix_299,Pix_300,Pix_301,Pix_302,Pix_303,Pix_304,Pix_305,Pix_306,Pix_307,Pix_308,Pix_309,Pix_310,Pix_311,Pix_312,Pix_313,Pix_314,Pix_315,Pix_316,Pix_317,Pix_318,Pix_319,Pix_320,Pix_321,Pix_322,Pix_323,Pix_324,Pix_325,Pix_326,Pix_327,Pix_328,Pix_329,Pix_330,Pix_331,Pix_332,Pix_333,Pix_334,Pix_335,Pix_336,Pix_337,Pix_338,Pix_339,Pix_340,Pix_341,Pix_342,Pix_343,Pix_344,Pix_345,Pix_346,Pix_347,Pix_348,Pix_349,Pix_350,Pix_351,Pix_352,Pix_353,Pix_354,Pix_355,Pix_356,Pix_357,Pix_358,Pix_359,Pix_360,Pix_361,Pix_362,Pix_363,Pix_364,Pix_365,Pix_366,Pix_367,Pix_368,Pix_369,Pix_370,Pix_371,Pix_372,Pix_373,Pix_374,Pix_375,Pix_376,Pix_377,Pix_378,Pix_379,Pix_380,Pix_381,Pix_382,Pix_383,Pix_384,Pix_385,Pix_386,Pix_387,Pix_388,Pix_389,Pix_390,Pix_391,Pix_392,Pix_393,Pix_394,Pix_395,Pix_396,Pix_397,Pix_398,Pix_399,Pix_400,Pix_401,Pix_402,Pix_403,Pix_404,Pix_405,Pix_406,Pix_407,Pix_408,Pix_409,Pix_410,Pix_411,Pix_412,Pix_413,Pix_414,Pix_415,Pix_416,Pix_417,Pix_418,Pix_419,Pix_420,Pix_421,Pix_422,Pix_423,Pix_424,Pix_425,Pix_426,Pix_427,Pix_428,Pix_429,Pix_430,Pix_431,Pix_432,Pix_433,Pix_434,Pix_435,Pix_436,Pix_437,Pix_438,Pix_439,Pix_440,Pix_441,Pix_442,Pix_443,Pix_444,Pix_445,Pix_446,Pix_447,Pix_448,Pix_449,Pix_450,Pix_451,Pix_452,Pix_453,Pix_454,Pix_455,Pix_456,Pix_457,Pix_458,Pix_459,Pix_460,Pix_461,Pix_462,Pix_463,Pix_464,Pix_465,Pix_466,Pix_467,Pix_468,Pix_469,Pix_470,Pix_471,Pix_472,Pix_473,Pix_474,Pix_475,Pix_476,Pix_477,Pix_478,Pix_479,Pix_480,Pix_481,Pix_482,Pix_483,Pix_484,Pix_485,Pix_486,Pix_487,Pix_488,Pix_489,Pix_490,Pix_491,Pix_492,Pix_493,Pix_494,Pix_495,Pix_496,Pix_497,Pix_498,Pix_499,Pix_500,Pix_501,Pix_502,Pix_503,Pix_504,Pix_505,Pix_506,Pix_507,Pix_508,Pix_509,Pix_510,Pix_511,Pix_512,Pix_513,Pix_514,Pix_515,Pix_516,Pix_517,Pix_518,Pix_519,Pix_520,Pix_521,Pix_522,Pix_523,Pix_524,Pix_525,Pix_526,Pix_527,Pix_528,Pix_529,Pix_530,Pix_531,Pix_532,Pix_533,Pix_534,Pix_535,Pix_536,Pix_537,Pix_538,Pix_539,Pix_540,Pix_541,Pix_542,Pix_543,Pix_544,Pix_545,Pix_546,Pix_547,Pix_548,Pix_549,Pix_550,Pix_551,Pix_552,Pix_553,Pix_554,Pix_555,Pix_556,Pix_557,Pix_558,Pix_559,Pix_560,Pix_561,Pix_562,Pix_563,Pix_564,Pix_565,Pix_566,Pix_567,Pix_568,Pix_569,Pix_570,Pix_571,Pix_572,Pix_573,Pix_574,Pix_575,Pix_576,Pix_577,Pix_578,Pix_579,Pix_580,Pix_581,Pix_582,Pix_583,Pix_584,Pix_585,Pix_586,Pix_587,Pix_588,Pix_589,Pix_590,Pix_591,Pix_592,Pix_593,Pix_594,Pix_595,Pix_596,Pix_597,Pix_598,Pix_599,Pix_600,Pix_601,Pix_602,Pix_603,Pix_604,Pix_605,Pix_606,Pix_607,Pix_608,Pix_609,Pix_610,Pix_611,Pix_612,Pix_613,Pix_614,Pix_615,Pix_616,Pix_617,Pix_618,Pix_619,Pix_620,Pix_621,Pix_622,Pix_623,Pix_624,Pix_625,Pix_626,Pix_627,Pix_628,Pix_629,Pix_630,Pix_631,Pix_632,Pix_633,Pix_634,Pix_635,Pix_636,Pix_637,Pix_638,Pix_639,Pix_640,Pix_641,Pix_642,Pix_643,Pix_644,Pix_645,Pix_646,Pix_647,Pix_648,Pix_649,Pix_650,Pix_651,Pix_652,Pix_653,Pix_654,Pix_655,Pix_656,Pix_657,Pix_658,Pix_659,Pix_660,Pix_661,Pix_662,Pix_663,Pix_664,Pix_665,Pix_666,Pix_667,Pix_668,Pix_669,Pix_670,Pix_671,Pix_672,Pix_673,Pix_674,Pix_675,Pix_676,Pix_677,Pix_678,Pix_679,Pix_680,Pix_681,Pix_682,Pix_683,Pix_684,Pix_685,Pix_686,Pix_687,Pix_688,Pix_689,Pix_690,Pix_691,Pix_692,Pix_693,Pix_694,Pix_695,Pix_696,Pix_697,Pix_698,Pix_699,Pix_700,Pix_701,Pix_702,Pix_703,Pix_704,Pix_705,Pix_706,Pix_707,Pix_708,Pix_709,Pix_710,Pix_711,Pix_712,Pix_713,Pix_714,Pix_715,Pix_716,Pix_717,Pix_718,Pix_719,Pix_720,Pix_721,Pix_722,Pix_723,Pix_724,Pix_725,Pix_726,Pix_727,Pix_728,Pix_729,Pix_730,Pix_731,Pix_732,Pix_733,Pix_734,Pix_735,Pix_736,Pix_737,Pix_738,Pix_739,Pix_740,Pix_741,Pix_742,Pix_743,Pix_744,Pix_745,Pix_746,Pix_747,Pix_748,Pix_749,Pix_750,Pix_751,Pix_752,Pix_753,Pix_754,Pix_755,Pix_756,Pix_757,Pix_758,Pix_759,Pix_760,Pix_761,Pix_762,Pix_763,Pix_764,Pix_765,Pix_766,Pix_767,Pix_768,Pix_769,Pix_770,Pix_771,Pix_772,Pix_773,Pix_774,Pix_775,Pix_776,Pix_777,Pix_778,Pix_779,Pix_780,Pix_781,Pix_782,Pix_783,Pix_784,
	Image_Number,
	Output_Valid
);

parameter NEURONS = 10;
parameter PIXEL_N = 785;
parameter WEIGHT_SIZE = 19;
parameter PIXEL_SIZE = 10;
parameter FPM_DELAY = 6;
parameter FPA_DELAY = 2;
parameter PARALLEL = 4;
parameter BUS_WIDTH = PIXEL_N/PARALLEL;
parameter VAL_SIZE = 26;

input clk;
input GlobalReset;
input Input_Valid;
input [WEIGHT_SIZE-1:0] Wgt_0_0;input [WEIGHT_SIZE-1:0] Wgt_0_1;input [WEIGHT_SIZE-1:0] Wgt_0_2;input [WEIGHT_SIZE-1:0] Wgt_0_3;input [WEIGHT_SIZE-1:0] Wgt_0_4;input [WEIGHT_SIZE-1:0] Wgt_0_5;input [WEIGHT_SIZE-1:0] Wgt_0_6;input [WEIGHT_SIZE-1:0] Wgt_0_7;input [WEIGHT_SIZE-1:0] Wgt_0_8;input [WEIGHT_SIZE-1:0] Wgt_0_9;input [WEIGHT_SIZE-1:0] Wgt_0_10;input [WEIGHT_SIZE-1:0] Wgt_0_11;input [WEIGHT_SIZE-1:0] Wgt_0_12;input [WEIGHT_SIZE-1:0] Wgt_0_13;input [WEIGHT_SIZE-1:0] Wgt_0_14;input [WEIGHT_SIZE-1:0] Wgt_0_15;input [WEIGHT_SIZE-1:0] Wgt_0_16;input [WEIGHT_SIZE-1:0] Wgt_0_17;input [WEIGHT_SIZE-1:0] Wgt_0_18;input [WEIGHT_SIZE-1:0] Wgt_0_19;input [WEIGHT_SIZE-1:0] Wgt_0_20;input [WEIGHT_SIZE-1:0] Wgt_0_21;input [WEIGHT_SIZE-1:0] Wgt_0_22;input [WEIGHT_SIZE-1:0] Wgt_0_23;input [WEIGHT_SIZE-1:0] Wgt_0_24;input [WEIGHT_SIZE-1:0] Wgt_0_25;input [WEIGHT_SIZE-1:0] Wgt_0_26;input [WEIGHT_SIZE-1:0] Wgt_0_27;input [WEIGHT_SIZE-1:0] Wgt_0_28;input [WEIGHT_SIZE-1:0] Wgt_0_29;input [WEIGHT_SIZE-1:0] Wgt_0_30;input [WEIGHT_SIZE-1:0] Wgt_0_31;input [WEIGHT_SIZE-1:0] Wgt_0_32;input [WEIGHT_SIZE-1:0] Wgt_0_33;input [WEIGHT_SIZE-1:0] Wgt_0_34;input [WEIGHT_SIZE-1:0] Wgt_0_35;input [WEIGHT_SIZE-1:0] Wgt_0_36;input [WEIGHT_SIZE-1:0] Wgt_0_37;input [WEIGHT_SIZE-1:0] Wgt_0_38;input [WEIGHT_SIZE-1:0] Wgt_0_39;input [WEIGHT_SIZE-1:0] Wgt_0_40;input [WEIGHT_SIZE-1:0] Wgt_0_41;input [WEIGHT_SIZE-1:0] Wgt_0_42;input [WEIGHT_SIZE-1:0] Wgt_0_43;input [WEIGHT_SIZE-1:0] Wgt_0_44;input [WEIGHT_SIZE-1:0] Wgt_0_45;input [WEIGHT_SIZE-1:0] Wgt_0_46;input [WEIGHT_SIZE-1:0] Wgt_0_47;input [WEIGHT_SIZE-1:0] Wgt_0_48;input [WEIGHT_SIZE-1:0] Wgt_0_49;input [WEIGHT_SIZE-1:0] Wgt_0_50;input [WEIGHT_SIZE-1:0] Wgt_0_51;input [WEIGHT_SIZE-1:0] Wgt_0_52;input [WEIGHT_SIZE-1:0] Wgt_0_53;input [WEIGHT_SIZE-1:0] Wgt_0_54;input [WEIGHT_SIZE-1:0] Wgt_0_55;input [WEIGHT_SIZE-1:0] Wgt_0_56;input [WEIGHT_SIZE-1:0] Wgt_0_57;input [WEIGHT_SIZE-1:0] Wgt_0_58;input [WEIGHT_SIZE-1:0] Wgt_0_59;input [WEIGHT_SIZE-1:0] Wgt_0_60;input [WEIGHT_SIZE-1:0] Wgt_0_61;input [WEIGHT_SIZE-1:0] Wgt_0_62;input [WEIGHT_SIZE-1:0] Wgt_0_63;input [WEIGHT_SIZE-1:0] Wgt_0_64;input [WEIGHT_SIZE-1:0] Wgt_0_65;input [WEIGHT_SIZE-1:0] Wgt_0_66;input [WEIGHT_SIZE-1:0] Wgt_0_67;input [WEIGHT_SIZE-1:0] Wgt_0_68;input [WEIGHT_SIZE-1:0] Wgt_0_69;input [WEIGHT_SIZE-1:0] Wgt_0_70;input [WEIGHT_SIZE-1:0] Wgt_0_71;input [WEIGHT_SIZE-1:0] Wgt_0_72;input [WEIGHT_SIZE-1:0] Wgt_0_73;input [WEIGHT_SIZE-1:0] Wgt_0_74;input [WEIGHT_SIZE-1:0] Wgt_0_75;input [WEIGHT_SIZE-1:0] Wgt_0_76;input [WEIGHT_SIZE-1:0] Wgt_0_77;input [WEIGHT_SIZE-1:0] Wgt_0_78;input [WEIGHT_SIZE-1:0] Wgt_0_79;input [WEIGHT_SIZE-1:0] Wgt_0_80;input [WEIGHT_SIZE-1:0] Wgt_0_81;input [WEIGHT_SIZE-1:0] Wgt_0_82;input [WEIGHT_SIZE-1:0] Wgt_0_83;input [WEIGHT_SIZE-1:0] Wgt_0_84;input [WEIGHT_SIZE-1:0] Wgt_0_85;input [WEIGHT_SIZE-1:0] Wgt_0_86;input [WEIGHT_SIZE-1:0] Wgt_0_87;input [WEIGHT_SIZE-1:0] Wgt_0_88;input [WEIGHT_SIZE-1:0] Wgt_0_89;input [WEIGHT_SIZE-1:0] Wgt_0_90;input [WEIGHT_SIZE-1:0] Wgt_0_91;input [WEIGHT_SIZE-1:0] Wgt_0_92;input [WEIGHT_SIZE-1:0] Wgt_0_93;input [WEIGHT_SIZE-1:0] Wgt_0_94;input [WEIGHT_SIZE-1:0] Wgt_0_95;input [WEIGHT_SIZE-1:0] Wgt_0_96;input [WEIGHT_SIZE-1:0] Wgt_0_97;input [WEIGHT_SIZE-1:0] Wgt_0_98;input [WEIGHT_SIZE-1:0] Wgt_0_99;input [WEIGHT_SIZE-1:0] Wgt_0_100;input [WEIGHT_SIZE-1:0] Wgt_0_101;input [WEIGHT_SIZE-1:0] Wgt_0_102;input [WEIGHT_SIZE-1:0] Wgt_0_103;input [WEIGHT_SIZE-1:0] Wgt_0_104;input [WEIGHT_SIZE-1:0] Wgt_0_105;input [WEIGHT_SIZE-1:0] Wgt_0_106;input [WEIGHT_SIZE-1:0] Wgt_0_107;input [WEIGHT_SIZE-1:0] Wgt_0_108;input [WEIGHT_SIZE-1:0] Wgt_0_109;input [WEIGHT_SIZE-1:0] Wgt_0_110;input [WEIGHT_SIZE-1:0] Wgt_0_111;input [WEIGHT_SIZE-1:0] Wgt_0_112;input [WEIGHT_SIZE-1:0] Wgt_0_113;input [WEIGHT_SIZE-1:0] Wgt_0_114;input [WEIGHT_SIZE-1:0] Wgt_0_115;input [WEIGHT_SIZE-1:0] Wgt_0_116;input [WEIGHT_SIZE-1:0] Wgt_0_117;input [WEIGHT_SIZE-1:0] Wgt_0_118;input [WEIGHT_SIZE-1:0] Wgt_0_119;input [WEIGHT_SIZE-1:0] Wgt_0_120;input [WEIGHT_SIZE-1:0] Wgt_0_121;input [WEIGHT_SIZE-1:0] Wgt_0_122;input [WEIGHT_SIZE-1:0] Wgt_0_123;input [WEIGHT_SIZE-1:0] Wgt_0_124;input [WEIGHT_SIZE-1:0] Wgt_0_125;input [WEIGHT_SIZE-1:0] Wgt_0_126;input [WEIGHT_SIZE-1:0] Wgt_0_127;input [WEIGHT_SIZE-1:0] Wgt_0_128;input [WEIGHT_SIZE-1:0] Wgt_0_129;input [WEIGHT_SIZE-1:0] Wgt_0_130;input [WEIGHT_SIZE-1:0] Wgt_0_131;input [WEIGHT_SIZE-1:0] Wgt_0_132;input [WEIGHT_SIZE-1:0] Wgt_0_133;input [WEIGHT_SIZE-1:0] Wgt_0_134;input [WEIGHT_SIZE-1:0] Wgt_0_135;input [WEIGHT_SIZE-1:0] Wgt_0_136;input [WEIGHT_SIZE-1:0] Wgt_0_137;input [WEIGHT_SIZE-1:0] Wgt_0_138;input [WEIGHT_SIZE-1:0] Wgt_0_139;input [WEIGHT_SIZE-1:0] Wgt_0_140;input [WEIGHT_SIZE-1:0] Wgt_0_141;input [WEIGHT_SIZE-1:0] Wgt_0_142;input [WEIGHT_SIZE-1:0] Wgt_0_143;input [WEIGHT_SIZE-1:0] Wgt_0_144;input [WEIGHT_SIZE-1:0] Wgt_0_145;input [WEIGHT_SIZE-1:0] Wgt_0_146;input [WEIGHT_SIZE-1:0] Wgt_0_147;input [WEIGHT_SIZE-1:0] Wgt_0_148;input [WEIGHT_SIZE-1:0] Wgt_0_149;input [WEIGHT_SIZE-1:0] Wgt_0_150;input [WEIGHT_SIZE-1:0] Wgt_0_151;input [WEIGHT_SIZE-1:0] Wgt_0_152;input [WEIGHT_SIZE-1:0] Wgt_0_153;input [WEIGHT_SIZE-1:0] Wgt_0_154;input [WEIGHT_SIZE-1:0] Wgt_0_155;input [WEIGHT_SIZE-1:0] Wgt_0_156;input [WEIGHT_SIZE-1:0] Wgt_0_157;input [WEIGHT_SIZE-1:0] Wgt_0_158;input [WEIGHT_SIZE-1:0] Wgt_0_159;input [WEIGHT_SIZE-1:0] Wgt_0_160;input [WEIGHT_SIZE-1:0] Wgt_0_161;input [WEIGHT_SIZE-1:0] Wgt_0_162;input [WEIGHT_SIZE-1:0] Wgt_0_163;input [WEIGHT_SIZE-1:0] Wgt_0_164;input [WEIGHT_SIZE-1:0] Wgt_0_165;input [WEIGHT_SIZE-1:0] Wgt_0_166;input [WEIGHT_SIZE-1:0] Wgt_0_167;input [WEIGHT_SIZE-1:0] Wgt_0_168;input [WEIGHT_SIZE-1:0] Wgt_0_169;input [WEIGHT_SIZE-1:0] Wgt_0_170;input [WEIGHT_SIZE-1:0] Wgt_0_171;input [WEIGHT_SIZE-1:0] Wgt_0_172;input [WEIGHT_SIZE-1:0] Wgt_0_173;input [WEIGHT_SIZE-1:0] Wgt_0_174;input [WEIGHT_SIZE-1:0] Wgt_0_175;input [WEIGHT_SIZE-1:0] Wgt_0_176;input [WEIGHT_SIZE-1:0] Wgt_0_177;input [WEIGHT_SIZE-1:0] Wgt_0_178;input [WEIGHT_SIZE-1:0] Wgt_0_179;input [WEIGHT_SIZE-1:0] Wgt_0_180;input [WEIGHT_SIZE-1:0] Wgt_0_181;input [WEIGHT_SIZE-1:0] Wgt_0_182;input [WEIGHT_SIZE-1:0] Wgt_0_183;input [WEIGHT_SIZE-1:0] Wgt_0_184;input [WEIGHT_SIZE-1:0] Wgt_0_185;input [WEIGHT_SIZE-1:0] Wgt_0_186;input [WEIGHT_SIZE-1:0] Wgt_0_187;input [WEIGHT_SIZE-1:0] Wgt_0_188;input [WEIGHT_SIZE-1:0] Wgt_0_189;input [WEIGHT_SIZE-1:0] Wgt_0_190;input [WEIGHT_SIZE-1:0] Wgt_0_191;input [WEIGHT_SIZE-1:0] Wgt_0_192;input [WEIGHT_SIZE-1:0] Wgt_0_193;input [WEIGHT_SIZE-1:0] Wgt_0_194;input [WEIGHT_SIZE-1:0] Wgt_0_195;input [WEIGHT_SIZE-1:0] Wgt_0_196;input [WEIGHT_SIZE-1:0] Wgt_0_197;input [WEIGHT_SIZE-1:0] Wgt_0_198;input [WEIGHT_SIZE-1:0] Wgt_0_199;input [WEIGHT_SIZE-1:0] Wgt_0_200;input [WEIGHT_SIZE-1:0] Wgt_0_201;input [WEIGHT_SIZE-1:0] Wgt_0_202;input [WEIGHT_SIZE-1:0] Wgt_0_203;input [WEIGHT_SIZE-1:0] Wgt_0_204;input [WEIGHT_SIZE-1:0] Wgt_0_205;input [WEIGHT_SIZE-1:0] Wgt_0_206;input [WEIGHT_SIZE-1:0] Wgt_0_207;input [WEIGHT_SIZE-1:0] Wgt_0_208;input [WEIGHT_SIZE-1:0] Wgt_0_209;input [WEIGHT_SIZE-1:0] Wgt_0_210;input [WEIGHT_SIZE-1:0] Wgt_0_211;input [WEIGHT_SIZE-1:0] Wgt_0_212;input [WEIGHT_SIZE-1:0] Wgt_0_213;input [WEIGHT_SIZE-1:0] Wgt_0_214;input [WEIGHT_SIZE-1:0] Wgt_0_215;input [WEIGHT_SIZE-1:0] Wgt_0_216;input [WEIGHT_SIZE-1:0] Wgt_0_217;input [WEIGHT_SIZE-1:0] Wgt_0_218;input [WEIGHT_SIZE-1:0] Wgt_0_219;input [WEIGHT_SIZE-1:0] Wgt_0_220;input [WEIGHT_SIZE-1:0] Wgt_0_221;input [WEIGHT_SIZE-1:0] Wgt_0_222;input [WEIGHT_SIZE-1:0] Wgt_0_223;input [WEIGHT_SIZE-1:0] Wgt_0_224;input [WEIGHT_SIZE-1:0] Wgt_0_225;input [WEIGHT_SIZE-1:0] Wgt_0_226;input [WEIGHT_SIZE-1:0] Wgt_0_227;input [WEIGHT_SIZE-1:0] Wgt_0_228;input [WEIGHT_SIZE-1:0] Wgt_0_229;input [WEIGHT_SIZE-1:0] Wgt_0_230;input [WEIGHT_SIZE-1:0] Wgt_0_231;input [WEIGHT_SIZE-1:0] Wgt_0_232;input [WEIGHT_SIZE-1:0] Wgt_0_233;input [WEIGHT_SIZE-1:0] Wgt_0_234;input [WEIGHT_SIZE-1:0] Wgt_0_235;input [WEIGHT_SIZE-1:0] Wgt_0_236;input [WEIGHT_SIZE-1:0] Wgt_0_237;input [WEIGHT_SIZE-1:0] Wgt_0_238;input [WEIGHT_SIZE-1:0] Wgt_0_239;input [WEIGHT_SIZE-1:0] Wgt_0_240;input [WEIGHT_SIZE-1:0] Wgt_0_241;input [WEIGHT_SIZE-1:0] Wgt_0_242;input [WEIGHT_SIZE-1:0] Wgt_0_243;input [WEIGHT_SIZE-1:0] Wgt_0_244;input [WEIGHT_SIZE-1:0] Wgt_0_245;input [WEIGHT_SIZE-1:0] Wgt_0_246;input [WEIGHT_SIZE-1:0] Wgt_0_247;input [WEIGHT_SIZE-1:0] Wgt_0_248;input [WEIGHT_SIZE-1:0] Wgt_0_249;input [WEIGHT_SIZE-1:0] Wgt_0_250;input [WEIGHT_SIZE-1:0] Wgt_0_251;input [WEIGHT_SIZE-1:0] Wgt_0_252;input [WEIGHT_SIZE-1:0] Wgt_0_253;input [WEIGHT_SIZE-1:0] Wgt_0_254;input [WEIGHT_SIZE-1:0] Wgt_0_255;input [WEIGHT_SIZE-1:0] Wgt_0_256;input [WEIGHT_SIZE-1:0] Wgt_0_257;input [WEIGHT_SIZE-1:0] Wgt_0_258;input [WEIGHT_SIZE-1:0] Wgt_0_259;input [WEIGHT_SIZE-1:0] Wgt_0_260;input [WEIGHT_SIZE-1:0] Wgt_0_261;input [WEIGHT_SIZE-1:0] Wgt_0_262;input [WEIGHT_SIZE-1:0] Wgt_0_263;input [WEIGHT_SIZE-1:0] Wgt_0_264;input [WEIGHT_SIZE-1:0] Wgt_0_265;input [WEIGHT_SIZE-1:0] Wgt_0_266;input [WEIGHT_SIZE-1:0] Wgt_0_267;input [WEIGHT_SIZE-1:0] Wgt_0_268;input [WEIGHT_SIZE-1:0] Wgt_0_269;input [WEIGHT_SIZE-1:0] Wgt_0_270;input [WEIGHT_SIZE-1:0] Wgt_0_271;input [WEIGHT_SIZE-1:0] Wgt_0_272;input [WEIGHT_SIZE-1:0] Wgt_0_273;input [WEIGHT_SIZE-1:0] Wgt_0_274;input [WEIGHT_SIZE-1:0] Wgt_0_275;input [WEIGHT_SIZE-1:0] Wgt_0_276;input [WEIGHT_SIZE-1:0] Wgt_0_277;input [WEIGHT_SIZE-1:0] Wgt_0_278;input [WEIGHT_SIZE-1:0] Wgt_0_279;input [WEIGHT_SIZE-1:0] Wgt_0_280;input [WEIGHT_SIZE-1:0] Wgt_0_281;input [WEIGHT_SIZE-1:0] Wgt_0_282;input [WEIGHT_SIZE-1:0] Wgt_0_283;input [WEIGHT_SIZE-1:0] Wgt_0_284;input [WEIGHT_SIZE-1:0] Wgt_0_285;input [WEIGHT_SIZE-1:0] Wgt_0_286;input [WEIGHT_SIZE-1:0] Wgt_0_287;input [WEIGHT_SIZE-1:0] Wgt_0_288;input [WEIGHT_SIZE-1:0] Wgt_0_289;input [WEIGHT_SIZE-1:0] Wgt_0_290;input [WEIGHT_SIZE-1:0] Wgt_0_291;input [WEIGHT_SIZE-1:0] Wgt_0_292;input [WEIGHT_SIZE-1:0] Wgt_0_293;input [WEIGHT_SIZE-1:0] Wgt_0_294;input [WEIGHT_SIZE-1:0] Wgt_0_295;input [WEIGHT_SIZE-1:0] Wgt_0_296;input [WEIGHT_SIZE-1:0] Wgt_0_297;input [WEIGHT_SIZE-1:0] Wgt_0_298;input [WEIGHT_SIZE-1:0] Wgt_0_299;input [WEIGHT_SIZE-1:0] Wgt_0_300;input [WEIGHT_SIZE-1:0] Wgt_0_301;input [WEIGHT_SIZE-1:0] Wgt_0_302;input [WEIGHT_SIZE-1:0] Wgt_0_303;input [WEIGHT_SIZE-1:0] Wgt_0_304;input [WEIGHT_SIZE-1:0] Wgt_0_305;input [WEIGHT_SIZE-1:0] Wgt_0_306;input [WEIGHT_SIZE-1:0] Wgt_0_307;input [WEIGHT_SIZE-1:0] Wgt_0_308;input [WEIGHT_SIZE-1:0] Wgt_0_309;input [WEIGHT_SIZE-1:0] Wgt_0_310;input [WEIGHT_SIZE-1:0] Wgt_0_311;input [WEIGHT_SIZE-1:0] Wgt_0_312;input [WEIGHT_SIZE-1:0] Wgt_0_313;input [WEIGHT_SIZE-1:0] Wgt_0_314;input [WEIGHT_SIZE-1:0] Wgt_0_315;input [WEIGHT_SIZE-1:0] Wgt_0_316;input [WEIGHT_SIZE-1:0] Wgt_0_317;input [WEIGHT_SIZE-1:0] Wgt_0_318;input [WEIGHT_SIZE-1:0] Wgt_0_319;input [WEIGHT_SIZE-1:0] Wgt_0_320;input [WEIGHT_SIZE-1:0] Wgt_0_321;input [WEIGHT_SIZE-1:0] Wgt_0_322;input [WEIGHT_SIZE-1:0] Wgt_0_323;input [WEIGHT_SIZE-1:0] Wgt_0_324;input [WEIGHT_SIZE-1:0] Wgt_0_325;input [WEIGHT_SIZE-1:0] Wgt_0_326;input [WEIGHT_SIZE-1:0] Wgt_0_327;input [WEIGHT_SIZE-1:0] Wgt_0_328;input [WEIGHT_SIZE-1:0] Wgt_0_329;input [WEIGHT_SIZE-1:0] Wgt_0_330;input [WEIGHT_SIZE-1:0] Wgt_0_331;input [WEIGHT_SIZE-1:0] Wgt_0_332;input [WEIGHT_SIZE-1:0] Wgt_0_333;input [WEIGHT_SIZE-1:0] Wgt_0_334;input [WEIGHT_SIZE-1:0] Wgt_0_335;input [WEIGHT_SIZE-1:0] Wgt_0_336;input [WEIGHT_SIZE-1:0] Wgt_0_337;input [WEIGHT_SIZE-1:0] Wgt_0_338;input [WEIGHT_SIZE-1:0] Wgt_0_339;input [WEIGHT_SIZE-1:0] Wgt_0_340;input [WEIGHT_SIZE-1:0] Wgt_0_341;input [WEIGHT_SIZE-1:0] Wgt_0_342;input [WEIGHT_SIZE-1:0] Wgt_0_343;input [WEIGHT_SIZE-1:0] Wgt_0_344;input [WEIGHT_SIZE-1:0] Wgt_0_345;input [WEIGHT_SIZE-1:0] Wgt_0_346;input [WEIGHT_SIZE-1:0] Wgt_0_347;input [WEIGHT_SIZE-1:0] Wgt_0_348;input [WEIGHT_SIZE-1:0] Wgt_0_349;input [WEIGHT_SIZE-1:0] Wgt_0_350;input [WEIGHT_SIZE-1:0] Wgt_0_351;input [WEIGHT_SIZE-1:0] Wgt_0_352;input [WEIGHT_SIZE-1:0] Wgt_0_353;input [WEIGHT_SIZE-1:0] Wgt_0_354;input [WEIGHT_SIZE-1:0] Wgt_0_355;input [WEIGHT_SIZE-1:0] Wgt_0_356;input [WEIGHT_SIZE-1:0] Wgt_0_357;input [WEIGHT_SIZE-1:0] Wgt_0_358;input [WEIGHT_SIZE-1:0] Wgt_0_359;input [WEIGHT_SIZE-1:0] Wgt_0_360;input [WEIGHT_SIZE-1:0] Wgt_0_361;input [WEIGHT_SIZE-1:0] Wgt_0_362;input [WEIGHT_SIZE-1:0] Wgt_0_363;input [WEIGHT_SIZE-1:0] Wgt_0_364;input [WEIGHT_SIZE-1:0] Wgt_0_365;input [WEIGHT_SIZE-1:0] Wgt_0_366;input [WEIGHT_SIZE-1:0] Wgt_0_367;input [WEIGHT_SIZE-1:0] Wgt_0_368;input [WEIGHT_SIZE-1:0] Wgt_0_369;input [WEIGHT_SIZE-1:0] Wgt_0_370;input [WEIGHT_SIZE-1:0] Wgt_0_371;input [WEIGHT_SIZE-1:0] Wgt_0_372;input [WEIGHT_SIZE-1:0] Wgt_0_373;input [WEIGHT_SIZE-1:0] Wgt_0_374;input [WEIGHT_SIZE-1:0] Wgt_0_375;input [WEIGHT_SIZE-1:0] Wgt_0_376;input [WEIGHT_SIZE-1:0] Wgt_0_377;input [WEIGHT_SIZE-1:0] Wgt_0_378;input [WEIGHT_SIZE-1:0] Wgt_0_379;input [WEIGHT_SIZE-1:0] Wgt_0_380;input [WEIGHT_SIZE-1:0] Wgt_0_381;input [WEIGHT_SIZE-1:0] Wgt_0_382;input [WEIGHT_SIZE-1:0] Wgt_0_383;input [WEIGHT_SIZE-1:0] Wgt_0_384;input [WEIGHT_SIZE-1:0] Wgt_0_385;input [WEIGHT_SIZE-1:0] Wgt_0_386;input [WEIGHT_SIZE-1:0] Wgt_0_387;input [WEIGHT_SIZE-1:0] Wgt_0_388;input [WEIGHT_SIZE-1:0] Wgt_0_389;input [WEIGHT_SIZE-1:0] Wgt_0_390;input [WEIGHT_SIZE-1:0] Wgt_0_391;input [WEIGHT_SIZE-1:0] Wgt_0_392;input [WEIGHT_SIZE-1:0] Wgt_0_393;input [WEIGHT_SIZE-1:0] Wgt_0_394;input [WEIGHT_SIZE-1:0] Wgt_0_395;input [WEIGHT_SIZE-1:0] Wgt_0_396;input [WEIGHT_SIZE-1:0] Wgt_0_397;input [WEIGHT_SIZE-1:0] Wgt_0_398;input [WEIGHT_SIZE-1:0] Wgt_0_399;input [WEIGHT_SIZE-1:0] Wgt_0_400;input [WEIGHT_SIZE-1:0] Wgt_0_401;input [WEIGHT_SIZE-1:0] Wgt_0_402;input [WEIGHT_SIZE-1:0] Wgt_0_403;input [WEIGHT_SIZE-1:0] Wgt_0_404;input [WEIGHT_SIZE-1:0] Wgt_0_405;input [WEIGHT_SIZE-1:0] Wgt_0_406;input [WEIGHT_SIZE-1:0] Wgt_0_407;input [WEIGHT_SIZE-1:0] Wgt_0_408;input [WEIGHT_SIZE-1:0] Wgt_0_409;input [WEIGHT_SIZE-1:0] Wgt_0_410;input [WEIGHT_SIZE-1:0] Wgt_0_411;input [WEIGHT_SIZE-1:0] Wgt_0_412;input [WEIGHT_SIZE-1:0] Wgt_0_413;input [WEIGHT_SIZE-1:0] Wgt_0_414;input [WEIGHT_SIZE-1:0] Wgt_0_415;input [WEIGHT_SIZE-1:0] Wgt_0_416;input [WEIGHT_SIZE-1:0] Wgt_0_417;input [WEIGHT_SIZE-1:0] Wgt_0_418;input [WEIGHT_SIZE-1:0] Wgt_0_419;input [WEIGHT_SIZE-1:0] Wgt_0_420;input [WEIGHT_SIZE-1:0] Wgt_0_421;input [WEIGHT_SIZE-1:0] Wgt_0_422;input [WEIGHT_SIZE-1:0] Wgt_0_423;input [WEIGHT_SIZE-1:0] Wgt_0_424;input [WEIGHT_SIZE-1:0] Wgt_0_425;input [WEIGHT_SIZE-1:0] Wgt_0_426;input [WEIGHT_SIZE-1:0] Wgt_0_427;input [WEIGHT_SIZE-1:0] Wgt_0_428;input [WEIGHT_SIZE-1:0] Wgt_0_429;input [WEIGHT_SIZE-1:0] Wgt_0_430;input [WEIGHT_SIZE-1:0] Wgt_0_431;input [WEIGHT_SIZE-1:0] Wgt_0_432;input [WEIGHT_SIZE-1:0] Wgt_0_433;input [WEIGHT_SIZE-1:0] Wgt_0_434;input [WEIGHT_SIZE-1:0] Wgt_0_435;input [WEIGHT_SIZE-1:0] Wgt_0_436;input [WEIGHT_SIZE-1:0] Wgt_0_437;input [WEIGHT_SIZE-1:0] Wgt_0_438;input [WEIGHT_SIZE-1:0] Wgt_0_439;input [WEIGHT_SIZE-1:0] Wgt_0_440;input [WEIGHT_SIZE-1:0] Wgt_0_441;input [WEIGHT_SIZE-1:0] Wgt_0_442;input [WEIGHT_SIZE-1:0] Wgt_0_443;input [WEIGHT_SIZE-1:0] Wgt_0_444;input [WEIGHT_SIZE-1:0] Wgt_0_445;input [WEIGHT_SIZE-1:0] Wgt_0_446;input [WEIGHT_SIZE-1:0] Wgt_0_447;input [WEIGHT_SIZE-1:0] Wgt_0_448;input [WEIGHT_SIZE-1:0] Wgt_0_449;input [WEIGHT_SIZE-1:0] Wgt_0_450;input [WEIGHT_SIZE-1:0] Wgt_0_451;input [WEIGHT_SIZE-1:0] Wgt_0_452;input [WEIGHT_SIZE-1:0] Wgt_0_453;input [WEIGHT_SIZE-1:0] Wgt_0_454;input [WEIGHT_SIZE-1:0] Wgt_0_455;input [WEIGHT_SIZE-1:0] Wgt_0_456;input [WEIGHT_SIZE-1:0] Wgt_0_457;input [WEIGHT_SIZE-1:0] Wgt_0_458;input [WEIGHT_SIZE-1:0] Wgt_0_459;input [WEIGHT_SIZE-1:0] Wgt_0_460;input [WEIGHT_SIZE-1:0] Wgt_0_461;input [WEIGHT_SIZE-1:0] Wgt_0_462;input [WEIGHT_SIZE-1:0] Wgt_0_463;input [WEIGHT_SIZE-1:0] Wgt_0_464;input [WEIGHT_SIZE-1:0] Wgt_0_465;input [WEIGHT_SIZE-1:0] Wgt_0_466;input [WEIGHT_SIZE-1:0] Wgt_0_467;input [WEIGHT_SIZE-1:0] Wgt_0_468;input [WEIGHT_SIZE-1:0] Wgt_0_469;input [WEIGHT_SIZE-1:0] Wgt_0_470;input [WEIGHT_SIZE-1:0] Wgt_0_471;input [WEIGHT_SIZE-1:0] Wgt_0_472;input [WEIGHT_SIZE-1:0] Wgt_0_473;input [WEIGHT_SIZE-1:0] Wgt_0_474;input [WEIGHT_SIZE-1:0] Wgt_0_475;input [WEIGHT_SIZE-1:0] Wgt_0_476;input [WEIGHT_SIZE-1:0] Wgt_0_477;input [WEIGHT_SIZE-1:0] Wgt_0_478;input [WEIGHT_SIZE-1:0] Wgt_0_479;input [WEIGHT_SIZE-1:0] Wgt_0_480;input [WEIGHT_SIZE-1:0] Wgt_0_481;input [WEIGHT_SIZE-1:0] Wgt_0_482;input [WEIGHT_SIZE-1:0] Wgt_0_483;input [WEIGHT_SIZE-1:0] Wgt_0_484;input [WEIGHT_SIZE-1:0] Wgt_0_485;input [WEIGHT_SIZE-1:0] Wgt_0_486;input [WEIGHT_SIZE-1:0] Wgt_0_487;input [WEIGHT_SIZE-1:0] Wgt_0_488;input [WEIGHT_SIZE-1:0] Wgt_0_489;input [WEIGHT_SIZE-1:0] Wgt_0_490;input [WEIGHT_SIZE-1:0] Wgt_0_491;input [WEIGHT_SIZE-1:0] Wgt_0_492;input [WEIGHT_SIZE-1:0] Wgt_0_493;input [WEIGHT_SIZE-1:0] Wgt_0_494;input [WEIGHT_SIZE-1:0] Wgt_0_495;input [WEIGHT_SIZE-1:0] Wgt_0_496;input [WEIGHT_SIZE-1:0] Wgt_0_497;input [WEIGHT_SIZE-1:0] Wgt_0_498;input [WEIGHT_SIZE-1:0] Wgt_0_499;input [WEIGHT_SIZE-1:0] Wgt_0_500;input [WEIGHT_SIZE-1:0] Wgt_0_501;input [WEIGHT_SIZE-1:0] Wgt_0_502;input [WEIGHT_SIZE-1:0] Wgt_0_503;input [WEIGHT_SIZE-1:0] Wgt_0_504;input [WEIGHT_SIZE-1:0] Wgt_0_505;input [WEIGHT_SIZE-1:0] Wgt_0_506;input [WEIGHT_SIZE-1:0] Wgt_0_507;input [WEIGHT_SIZE-1:0] Wgt_0_508;input [WEIGHT_SIZE-1:0] Wgt_0_509;input [WEIGHT_SIZE-1:0] Wgt_0_510;input [WEIGHT_SIZE-1:0] Wgt_0_511;input [WEIGHT_SIZE-1:0] Wgt_0_512;input [WEIGHT_SIZE-1:0] Wgt_0_513;input [WEIGHT_SIZE-1:0] Wgt_0_514;input [WEIGHT_SIZE-1:0] Wgt_0_515;input [WEIGHT_SIZE-1:0] Wgt_0_516;input [WEIGHT_SIZE-1:0] Wgt_0_517;input [WEIGHT_SIZE-1:0] Wgt_0_518;input [WEIGHT_SIZE-1:0] Wgt_0_519;input [WEIGHT_SIZE-1:0] Wgt_0_520;input [WEIGHT_SIZE-1:0] Wgt_0_521;input [WEIGHT_SIZE-1:0] Wgt_0_522;input [WEIGHT_SIZE-1:0] Wgt_0_523;input [WEIGHT_SIZE-1:0] Wgt_0_524;input [WEIGHT_SIZE-1:0] Wgt_0_525;input [WEIGHT_SIZE-1:0] Wgt_0_526;input [WEIGHT_SIZE-1:0] Wgt_0_527;input [WEIGHT_SIZE-1:0] Wgt_0_528;input [WEIGHT_SIZE-1:0] Wgt_0_529;input [WEIGHT_SIZE-1:0] Wgt_0_530;input [WEIGHT_SIZE-1:0] Wgt_0_531;input [WEIGHT_SIZE-1:0] Wgt_0_532;input [WEIGHT_SIZE-1:0] Wgt_0_533;input [WEIGHT_SIZE-1:0] Wgt_0_534;input [WEIGHT_SIZE-1:0] Wgt_0_535;input [WEIGHT_SIZE-1:0] Wgt_0_536;input [WEIGHT_SIZE-1:0] Wgt_0_537;input [WEIGHT_SIZE-1:0] Wgt_0_538;input [WEIGHT_SIZE-1:0] Wgt_0_539;input [WEIGHT_SIZE-1:0] Wgt_0_540;input [WEIGHT_SIZE-1:0] Wgt_0_541;input [WEIGHT_SIZE-1:0] Wgt_0_542;input [WEIGHT_SIZE-1:0] Wgt_0_543;input [WEIGHT_SIZE-1:0] Wgt_0_544;input [WEIGHT_SIZE-1:0] Wgt_0_545;input [WEIGHT_SIZE-1:0] Wgt_0_546;input [WEIGHT_SIZE-1:0] Wgt_0_547;input [WEIGHT_SIZE-1:0] Wgt_0_548;input [WEIGHT_SIZE-1:0] Wgt_0_549;input [WEIGHT_SIZE-1:0] Wgt_0_550;input [WEIGHT_SIZE-1:0] Wgt_0_551;input [WEIGHT_SIZE-1:0] Wgt_0_552;input [WEIGHT_SIZE-1:0] Wgt_0_553;input [WEIGHT_SIZE-1:0] Wgt_0_554;input [WEIGHT_SIZE-1:0] Wgt_0_555;input [WEIGHT_SIZE-1:0] Wgt_0_556;input [WEIGHT_SIZE-1:0] Wgt_0_557;input [WEIGHT_SIZE-1:0] Wgt_0_558;input [WEIGHT_SIZE-1:0] Wgt_0_559;input [WEIGHT_SIZE-1:0] Wgt_0_560;input [WEIGHT_SIZE-1:0] Wgt_0_561;input [WEIGHT_SIZE-1:0] Wgt_0_562;input [WEIGHT_SIZE-1:0] Wgt_0_563;input [WEIGHT_SIZE-1:0] Wgt_0_564;input [WEIGHT_SIZE-1:0] Wgt_0_565;input [WEIGHT_SIZE-1:0] Wgt_0_566;input [WEIGHT_SIZE-1:0] Wgt_0_567;input [WEIGHT_SIZE-1:0] Wgt_0_568;input [WEIGHT_SIZE-1:0] Wgt_0_569;input [WEIGHT_SIZE-1:0] Wgt_0_570;input [WEIGHT_SIZE-1:0] Wgt_0_571;input [WEIGHT_SIZE-1:0] Wgt_0_572;input [WEIGHT_SIZE-1:0] Wgt_0_573;input [WEIGHT_SIZE-1:0] Wgt_0_574;input [WEIGHT_SIZE-1:0] Wgt_0_575;input [WEIGHT_SIZE-1:0] Wgt_0_576;input [WEIGHT_SIZE-1:0] Wgt_0_577;input [WEIGHT_SIZE-1:0] Wgt_0_578;input [WEIGHT_SIZE-1:0] Wgt_0_579;input [WEIGHT_SIZE-1:0] Wgt_0_580;input [WEIGHT_SIZE-1:0] Wgt_0_581;input [WEIGHT_SIZE-1:0] Wgt_0_582;input [WEIGHT_SIZE-1:0] Wgt_0_583;input [WEIGHT_SIZE-1:0] Wgt_0_584;input [WEIGHT_SIZE-1:0] Wgt_0_585;input [WEIGHT_SIZE-1:0] Wgt_0_586;input [WEIGHT_SIZE-1:0] Wgt_0_587;input [WEIGHT_SIZE-1:0] Wgt_0_588;input [WEIGHT_SIZE-1:0] Wgt_0_589;input [WEIGHT_SIZE-1:0] Wgt_0_590;input [WEIGHT_SIZE-1:0] Wgt_0_591;input [WEIGHT_SIZE-1:0] Wgt_0_592;input [WEIGHT_SIZE-1:0] Wgt_0_593;input [WEIGHT_SIZE-1:0] Wgt_0_594;input [WEIGHT_SIZE-1:0] Wgt_0_595;input [WEIGHT_SIZE-1:0] Wgt_0_596;input [WEIGHT_SIZE-1:0] Wgt_0_597;input [WEIGHT_SIZE-1:0] Wgt_0_598;input [WEIGHT_SIZE-1:0] Wgt_0_599;input [WEIGHT_SIZE-1:0] Wgt_0_600;input [WEIGHT_SIZE-1:0] Wgt_0_601;input [WEIGHT_SIZE-1:0] Wgt_0_602;input [WEIGHT_SIZE-1:0] Wgt_0_603;input [WEIGHT_SIZE-1:0] Wgt_0_604;input [WEIGHT_SIZE-1:0] Wgt_0_605;input [WEIGHT_SIZE-1:0] Wgt_0_606;input [WEIGHT_SIZE-1:0] Wgt_0_607;input [WEIGHT_SIZE-1:0] Wgt_0_608;input [WEIGHT_SIZE-1:0] Wgt_0_609;input [WEIGHT_SIZE-1:0] Wgt_0_610;input [WEIGHT_SIZE-1:0] Wgt_0_611;input [WEIGHT_SIZE-1:0] Wgt_0_612;input [WEIGHT_SIZE-1:0] Wgt_0_613;input [WEIGHT_SIZE-1:0] Wgt_0_614;input [WEIGHT_SIZE-1:0] Wgt_0_615;input [WEIGHT_SIZE-1:0] Wgt_0_616;input [WEIGHT_SIZE-1:0] Wgt_0_617;input [WEIGHT_SIZE-1:0] Wgt_0_618;input [WEIGHT_SIZE-1:0] Wgt_0_619;input [WEIGHT_SIZE-1:0] Wgt_0_620;input [WEIGHT_SIZE-1:0] Wgt_0_621;input [WEIGHT_SIZE-1:0] Wgt_0_622;input [WEIGHT_SIZE-1:0] Wgt_0_623;input [WEIGHT_SIZE-1:0] Wgt_0_624;input [WEIGHT_SIZE-1:0] Wgt_0_625;input [WEIGHT_SIZE-1:0] Wgt_0_626;input [WEIGHT_SIZE-1:0] Wgt_0_627;input [WEIGHT_SIZE-1:0] Wgt_0_628;input [WEIGHT_SIZE-1:0] Wgt_0_629;input [WEIGHT_SIZE-1:0] Wgt_0_630;input [WEIGHT_SIZE-1:0] Wgt_0_631;input [WEIGHT_SIZE-1:0] Wgt_0_632;input [WEIGHT_SIZE-1:0] Wgt_0_633;input [WEIGHT_SIZE-1:0] Wgt_0_634;input [WEIGHT_SIZE-1:0] Wgt_0_635;input [WEIGHT_SIZE-1:0] Wgt_0_636;input [WEIGHT_SIZE-1:0] Wgt_0_637;input [WEIGHT_SIZE-1:0] Wgt_0_638;input [WEIGHT_SIZE-1:0] Wgt_0_639;input [WEIGHT_SIZE-1:0] Wgt_0_640;input [WEIGHT_SIZE-1:0] Wgt_0_641;input [WEIGHT_SIZE-1:0] Wgt_0_642;input [WEIGHT_SIZE-1:0] Wgt_0_643;input [WEIGHT_SIZE-1:0] Wgt_0_644;input [WEIGHT_SIZE-1:0] Wgt_0_645;input [WEIGHT_SIZE-1:0] Wgt_0_646;input [WEIGHT_SIZE-1:0] Wgt_0_647;input [WEIGHT_SIZE-1:0] Wgt_0_648;input [WEIGHT_SIZE-1:0] Wgt_0_649;input [WEIGHT_SIZE-1:0] Wgt_0_650;input [WEIGHT_SIZE-1:0] Wgt_0_651;input [WEIGHT_SIZE-1:0] Wgt_0_652;input [WEIGHT_SIZE-1:0] Wgt_0_653;input [WEIGHT_SIZE-1:0] Wgt_0_654;input [WEIGHT_SIZE-1:0] Wgt_0_655;input [WEIGHT_SIZE-1:0] Wgt_0_656;input [WEIGHT_SIZE-1:0] Wgt_0_657;input [WEIGHT_SIZE-1:0] Wgt_0_658;input [WEIGHT_SIZE-1:0] Wgt_0_659;input [WEIGHT_SIZE-1:0] Wgt_0_660;input [WEIGHT_SIZE-1:0] Wgt_0_661;input [WEIGHT_SIZE-1:0] Wgt_0_662;input [WEIGHT_SIZE-1:0] Wgt_0_663;input [WEIGHT_SIZE-1:0] Wgt_0_664;input [WEIGHT_SIZE-1:0] Wgt_0_665;input [WEIGHT_SIZE-1:0] Wgt_0_666;input [WEIGHT_SIZE-1:0] Wgt_0_667;input [WEIGHT_SIZE-1:0] Wgt_0_668;input [WEIGHT_SIZE-1:0] Wgt_0_669;input [WEIGHT_SIZE-1:0] Wgt_0_670;input [WEIGHT_SIZE-1:0] Wgt_0_671;input [WEIGHT_SIZE-1:0] Wgt_0_672;input [WEIGHT_SIZE-1:0] Wgt_0_673;input [WEIGHT_SIZE-1:0] Wgt_0_674;input [WEIGHT_SIZE-1:0] Wgt_0_675;input [WEIGHT_SIZE-1:0] Wgt_0_676;input [WEIGHT_SIZE-1:0] Wgt_0_677;input [WEIGHT_SIZE-1:0] Wgt_0_678;input [WEIGHT_SIZE-1:0] Wgt_0_679;input [WEIGHT_SIZE-1:0] Wgt_0_680;input [WEIGHT_SIZE-1:0] Wgt_0_681;input [WEIGHT_SIZE-1:0] Wgt_0_682;input [WEIGHT_SIZE-1:0] Wgt_0_683;input [WEIGHT_SIZE-1:0] Wgt_0_684;input [WEIGHT_SIZE-1:0] Wgt_0_685;input [WEIGHT_SIZE-1:0] Wgt_0_686;input [WEIGHT_SIZE-1:0] Wgt_0_687;input [WEIGHT_SIZE-1:0] Wgt_0_688;input [WEIGHT_SIZE-1:0] Wgt_0_689;input [WEIGHT_SIZE-1:0] Wgt_0_690;input [WEIGHT_SIZE-1:0] Wgt_0_691;input [WEIGHT_SIZE-1:0] Wgt_0_692;input [WEIGHT_SIZE-1:0] Wgt_0_693;input [WEIGHT_SIZE-1:0] Wgt_0_694;input [WEIGHT_SIZE-1:0] Wgt_0_695;input [WEIGHT_SIZE-1:0] Wgt_0_696;input [WEIGHT_SIZE-1:0] Wgt_0_697;input [WEIGHT_SIZE-1:0] Wgt_0_698;input [WEIGHT_SIZE-1:0] Wgt_0_699;input [WEIGHT_SIZE-1:0] Wgt_0_700;input [WEIGHT_SIZE-1:0] Wgt_0_701;input [WEIGHT_SIZE-1:0] Wgt_0_702;input [WEIGHT_SIZE-1:0] Wgt_0_703;input [WEIGHT_SIZE-1:0] Wgt_0_704;input [WEIGHT_SIZE-1:0] Wgt_0_705;input [WEIGHT_SIZE-1:0] Wgt_0_706;input [WEIGHT_SIZE-1:0] Wgt_0_707;input [WEIGHT_SIZE-1:0] Wgt_0_708;input [WEIGHT_SIZE-1:0] Wgt_0_709;input [WEIGHT_SIZE-1:0] Wgt_0_710;input [WEIGHT_SIZE-1:0] Wgt_0_711;input [WEIGHT_SIZE-1:0] Wgt_0_712;input [WEIGHT_SIZE-1:0] Wgt_0_713;input [WEIGHT_SIZE-1:0] Wgt_0_714;input [WEIGHT_SIZE-1:0] Wgt_0_715;input [WEIGHT_SIZE-1:0] Wgt_0_716;input [WEIGHT_SIZE-1:0] Wgt_0_717;input [WEIGHT_SIZE-1:0] Wgt_0_718;input [WEIGHT_SIZE-1:0] Wgt_0_719;input [WEIGHT_SIZE-1:0] Wgt_0_720;input [WEIGHT_SIZE-1:0] Wgt_0_721;input [WEIGHT_SIZE-1:0] Wgt_0_722;input [WEIGHT_SIZE-1:0] Wgt_0_723;input [WEIGHT_SIZE-1:0] Wgt_0_724;input [WEIGHT_SIZE-1:0] Wgt_0_725;input [WEIGHT_SIZE-1:0] Wgt_0_726;input [WEIGHT_SIZE-1:0] Wgt_0_727;input [WEIGHT_SIZE-1:0] Wgt_0_728;input [WEIGHT_SIZE-1:0] Wgt_0_729;input [WEIGHT_SIZE-1:0] Wgt_0_730;input [WEIGHT_SIZE-1:0] Wgt_0_731;input [WEIGHT_SIZE-1:0] Wgt_0_732;input [WEIGHT_SIZE-1:0] Wgt_0_733;input [WEIGHT_SIZE-1:0] Wgt_0_734;input [WEIGHT_SIZE-1:0] Wgt_0_735;input [WEIGHT_SIZE-1:0] Wgt_0_736;input [WEIGHT_SIZE-1:0] Wgt_0_737;input [WEIGHT_SIZE-1:0] Wgt_0_738;input [WEIGHT_SIZE-1:0] Wgt_0_739;input [WEIGHT_SIZE-1:0] Wgt_0_740;input [WEIGHT_SIZE-1:0] Wgt_0_741;input [WEIGHT_SIZE-1:0] Wgt_0_742;input [WEIGHT_SIZE-1:0] Wgt_0_743;input [WEIGHT_SIZE-1:0] Wgt_0_744;input [WEIGHT_SIZE-1:0] Wgt_0_745;input [WEIGHT_SIZE-1:0] Wgt_0_746;input [WEIGHT_SIZE-1:0] Wgt_0_747;input [WEIGHT_SIZE-1:0] Wgt_0_748;input [WEIGHT_SIZE-1:0] Wgt_0_749;input [WEIGHT_SIZE-1:0] Wgt_0_750;input [WEIGHT_SIZE-1:0] Wgt_0_751;input [WEIGHT_SIZE-1:0] Wgt_0_752;input [WEIGHT_SIZE-1:0] Wgt_0_753;input [WEIGHT_SIZE-1:0] Wgt_0_754;input [WEIGHT_SIZE-1:0] Wgt_0_755;input [WEIGHT_SIZE-1:0] Wgt_0_756;input [WEIGHT_SIZE-1:0] Wgt_0_757;input [WEIGHT_SIZE-1:0] Wgt_0_758;input [WEIGHT_SIZE-1:0] Wgt_0_759;input [WEIGHT_SIZE-1:0] Wgt_0_760;input [WEIGHT_SIZE-1:0] Wgt_0_761;input [WEIGHT_SIZE-1:0] Wgt_0_762;input [WEIGHT_SIZE-1:0] Wgt_0_763;input [WEIGHT_SIZE-1:0] Wgt_0_764;input [WEIGHT_SIZE-1:0] Wgt_0_765;input [WEIGHT_SIZE-1:0] Wgt_0_766;input [WEIGHT_SIZE-1:0] Wgt_0_767;input [WEIGHT_SIZE-1:0] Wgt_0_768;input [WEIGHT_SIZE-1:0] Wgt_0_769;input [WEIGHT_SIZE-1:0] Wgt_0_770;input [WEIGHT_SIZE-1:0] Wgt_0_771;input [WEIGHT_SIZE-1:0] Wgt_0_772;input [WEIGHT_SIZE-1:0] Wgt_0_773;input [WEIGHT_SIZE-1:0] Wgt_0_774;input [WEIGHT_SIZE-1:0] Wgt_0_775;input [WEIGHT_SIZE-1:0] Wgt_0_776;input [WEIGHT_SIZE-1:0] Wgt_0_777;input [WEIGHT_SIZE-1:0] Wgt_0_778;input [WEIGHT_SIZE-1:0] Wgt_0_779;input [WEIGHT_SIZE-1:0] Wgt_0_780;input [WEIGHT_SIZE-1:0] Wgt_0_781;input [WEIGHT_SIZE-1:0] Wgt_0_782;input [WEIGHT_SIZE-1:0] Wgt_0_783;input [WEIGHT_SIZE-1:0] Wgt_0_784;input [WEIGHT_SIZE-1:0] Wgt_1_0;input [WEIGHT_SIZE-1:0] Wgt_1_1;input [WEIGHT_SIZE-1:0] Wgt_1_2;input [WEIGHT_SIZE-1:0] Wgt_1_3;input [WEIGHT_SIZE-1:0] Wgt_1_4;input [WEIGHT_SIZE-1:0] Wgt_1_5;input [WEIGHT_SIZE-1:0] Wgt_1_6;input [WEIGHT_SIZE-1:0] Wgt_1_7;input [WEIGHT_SIZE-1:0] Wgt_1_8;input [WEIGHT_SIZE-1:0] Wgt_1_9;input [WEIGHT_SIZE-1:0] Wgt_1_10;input [WEIGHT_SIZE-1:0] Wgt_1_11;input [WEIGHT_SIZE-1:0] Wgt_1_12;input [WEIGHT_SIZE-1:0] Wgt_1_13;input [WEIGHT_SIZE-1:0] Wgt_1_14;input [WEIGHT_SIZE-1:0] Wgt_1_15;input [WEIGHT_SIZE-1:0] Wgt_1_16;input [WEIGHT_SIZE-1:0] Wgt_1_17;input [WEIGHT_SIZE-1:0] Wgt_1_18;input [WEIGHT_SIZE-1:0] Wgt_1_19;input [WEIGHT_SIZE-1:0] Wgt_1_20;input [WEIGHT_SIZE-1:0] Wgt_1_21;input [WEIGHT_SIZE-1:0] Wgt_1_22;input [WEIGHT_SIZE-1:0] Wgt_1_23;input [WEIGHT_SIZE-1:0] Wgt_1_24;input [WEIGHT_SIZE-1:0] Wgt_1_25;input [WEIGHT_SIZE-1:0] Wgt_1_26;input [WEIGHT_SIZE-1:0] Wgt_1_27;input [WEIGHT_SIZE-1:0] Wgt_1_28;input [WEIGHT_SIZE-1:0] Wgt_1_29;input [WEIGHT_SIZE-1:0] Wgt_1_30;input [WEIGHT_SIZE-1:0] Wgt_1_31;input [WEIGHT_SIZE-1:0] Wgt_1_32;input [WEIGHT_SIZE-1:0] Wgt_1_33;input [WEIGHT_SIZE-1:0] Wgt_1_34;input [WEIGHT_SIZE-1:0] Wgt_1_35;input [WEIGHT_SIZE-1:0] Wgt_1_36;input [WEIGHT_SIZE-1:0] Wgt_1_37;input [WEIGHT_SIZE-1:0] Wgt_1_38;input [WEIGHT_SIZE-1:0] Wgt_1_39;input [WEIGHT_SIZE-1:0] Wgt_1_40;input [WEIGHT_SIZE-1:0] Wgt_1_41;input [WEIGHT_SIZE-1:0] Wgt_1_42;input [WEIGHT_SIZE-1:0] Wgt_1_43;input [WEIGHT_SIZE-1:0] Wgt_1_44;input [WEIGHT_SIZE-1:0] Wgt_1_45;input [WEIGHT_SIZE-1:0] Wgt_1_46;input [WEIGHT_SIZE-1:0] Wgt_1_47;input [WEIGHT_SIZE-1:0] Wgt_1_48;input [WEIGHT_SIZE-1:0] Wgt_1_49;input [WEIGHT_SIZE-1:0] Wgt_1_50;input [WEIGHT_SIZE-1:0] Wgt_1_51;input [WEIGHT_SIZE-1:0] Wgt_1_52;input [WEIGHT_SIZE-1:0] Wgt_1_53;input [WEIGHT_SIZE-1:0] Wgt_1_54;input [WEIGHT_SIZE-1:0] Wgt_1_55;input [WEIGHT_SIZE-1:0] Wgt_1_56;input [WEIGHT_SIZE-1:0] Wgt_1_57;input [WEIGHT_SIZE-1:0] Wgt_1_58;input [WEIGHT_SIZE-1:0] Wgt_1_59;input [WEIGHT_SIZE-1:0] Wgt_1_60;input [WEIGHT_SIZE-1:0] Wgt_1_61;input [WEIGHT_SIZE-1:0] Wgt_1_62;input [WEIGHT_SIZE-1:0] Wgt_1_63;input [WEIGHT_SIZE-1:0] Wgt_1_64;input [WEIGHT_SIZE-1:0] Wgt_1_65;input [WEIGHT_SIZE-1:0] Wgt_1_66;input [WEIGHT_SIZE-1:0] Wgt_1_67;input [WEIGHT_SIZE-1:0] Wgt_1_68;input [WEIGHT_SIZE-1:0] Wgt_1_69;input [WEIGHT_SIZE-1:0] Wgt_1_70;input [WEIGHT_SIZE-1:0] Wgt_1_71;input [WEIGHT_SIZE-1:0] Wgt_1_72;input [WEIGHT_SIZE-1:0] Wgt_1_73;input [WEIGHT_SIZE-1:0] Wgt_1_74;input [WEIGHT_SIZE-1:0] Wgt_1_75;input [WEIGHT_SIZE-1:0] Wgt_1_76;input [WEIGHT_SIZE-1:0] Wgt_1_77;input [WEIGHT_SIZE-1:0] Wgt_1_78;input [WEIGHT_SIZE-1:0] Wgt_1_79;input [WEIGHT_SIZE-1:0] Wgt_1_80;input [WEIGHT_SIZE-1:0] Wgt_1_81;input [WEIGHT_SIZE-1:0] Wgt_1_82;input [WEIGHT_SIZE-1:0] Wgt_1_83;input [WEIGHT_SIZE-1:0] Wgt_1_84;input [WEIGHT_SIZE-1:0] Wgt_1_85;input [WEIGHT_SIZE-1:0] Wgt_1_86;input [WEIGHT_SIZE-1:0] Wgt_1_87;input [WEIGHT_SIZE-1:0] Wgt_1_88;input [WEIGHT_SIZE-1:0] Wgt_1_89;input [WEIGHT_SIZE-1:0] Wgt_1_90;input [WEIGHT_SIZE-1:0] Wgt_1_91;input [WEIGHT_SIZE-1:0] Wgt_1_92;input [WEIGHT_SIZE-1:0] Wgt_1_93;input [WEIGHT_SIZE-1:0] Wgt_1_94;input [WEIGHT_SIZE-1:0] Wgt_1_95;input [WEIGHT_SIZE-1:0] Wgt_1_96;input [WEIGHT_SIZE-1:0] Wgt_1_97;input [WEIGHT_SIZE-1:0] Wgt_1_98;input [WEIGHT_SIZE-1:0] Wgt_1_99;input [WEIGHT_SIZE-1:0] Wgt_1_100;input [WEIGHT_SIZE-1:0] Wgt_1_101;input [WEIGHT_SIZE-1:0] Wgt_1_102;input [WEIGHT_SIZE-1:0] Wgt_1_103;input [WEIGHT_SIZE-1:0] Wgt_1_104;input [WEIGHT_SIZE-1:0] Wgt_1_105;input [WEIGHT_SIZE-1:0] Wgt_1_106;input [WEIGHT_SIZE-1:0] Wgt_1_107;input [WEIGHT_SIZE-1:0] Wgt_1_108;input [WEIGHT_SIZE-1:0] Wgt_1_109;input [WEIGHT_SIZE-1:0] Wgt_1_110;input [WEIGHT_SIZE-1:0] Wgt_1_111;input [WEIGHT_SIZE-1:0] Wgt_1_112;input [WEIGHT_SIZE-1:0] Wgt_1_113;input [WEIGHT_SIZE-1:0] Wgt_1_114;input [WEIGHT_SIZE-1:0] Wgt_1_115;input [WEIGHT_SIZE-1:0] Wgt_1_116;input [WEIGHT_SIZE-1:0] Wgt_1_117;input [WEIGHT_SIZE-1:0] Wgt_1_118;input [WEIGHT_SIZE-1:0] Wgt_1_119;input [WEIGHT_SIZE-1:0] Wgt_1_120;input [WEIGHT_SIZE-1:0] Wgt_1_121;input [WEIGHT_SIZE-1:0] Wgt_1_122;input [WEIGHT_SIZE-1:0] Wgt_1_123;input [WEIGHT_SIZE-1:0] Wgt_1_124;input [WEIGHT_SIZE-1:0] Wgt_1_125;input [WEIGHT_SIZE-1:0] Wgt_1_126;input [WEIGHT_SIZE-1:0] Wgt_1_127;input [WEIGHT_SIZE-1:0] Wgt_1_128;input [WEIGHT_SIZE-1:0] Wgt_1_129;input [WEIGHT_SIZE-1:0] Wgt_1_130;input [WEIGHT_SIZE-1:0] Wgt_1_131;input [WEIGHT_SIZE-1:0] Wgt_1_132;input [WEIGHT_SIZE-1:0] Wgt_1_133;input [WEIGHT_SIZE-1:0] Wgt_1_134;input [WEIGHT_SIZE-1:0] Wgt_1_135;input [WEIGHT_SIZE-1:0] Wgt_1_136;input [WEIGHT_SIZE-1:0] Wgt_1_137;input [WEIGHT_SIZE-1:0] Wgt_1_138;input [WEIGHT_SIZE-1:0] Wgt_1_139;input [WEIGHT_SIZE-1:0] Wgt_1_140;input [WEIGHT_SIZE-1:0] Wgt_1_141;input [WEIGHT_SIZE-1:0] Wgt_1_142;input [WEIGHT_SIZE-1:0] Wgt_1_143;input [WEIGHT_SIZE-1:0] Wgt_1_144;input [WEIGHT_SIZE-1:0] Wgt_1_145;input [WEIGHT_SIZE-1:0] Wgt_1_146;input [WEIGHT_SIZE-1:0] Wgt_1_147;input [WEIGHT_SIZE-1:0] Wgt_1_148;input [WEIGHT_SIZE-1:0] Wgt_1_149;input [WEIGHT_SIZE-1:0] Wgt_1_150;input [WEIGHT_SIZE-1:0] Wgt_1_151;input [WEIGHT_SIZE-1:0] Wgt_1_152;input [WEIGHT_SIZE-1:0] Wgt_1_153;input [WEIGHT_SIZE-1:0] Wgt_1_154;input [WEIGHT_SIZE-1:0] Wgt_1_155;input [WEIGHT_SIZE-1:0] Wgt_1_156;input [WEIGHT_SIZE-1:0] Wgt_1_157;input [WEIGHT_SIZE-1:0] Wgt_1_158;input [WEIGHT_SIZE-1:0] Wgt_1_159;input [WEIGHT_SIZE-1:0] Wgt_1_160;input [WEIGHT_SIZE-1:0] Wgt_1_161;input [WEIGHT_SIZE-1:0] Wgt_1_162;input [WEIGHT_SIZE-1:0] Wgt_1_163;input [WEIGHT_SIZE-1:0] Wgt_1_164;input [WEIGHT_SIZE-1:0] Wgt_1_165;input [WEIGHT_SIZE-1:0] Wgt_1_166;input [WEIGHT_SIZE-1:0] Wgt_1_167;input [WEIGHT_SIZE-1:0] Wgt_1_168;input [WEIGHT_SIZE-1:0] Wgt_1_169;input [WEIGHT_SIZE-1:0] Wgt_1_170;input [WEIGHT_SIZE-1:0] Wgt_1_171;input [WEIGHT_SIZE-1:0] Wgt_1_172;input [WEIGHT_SIZE-1:0] Wgt_1_173;input [WEIGHT_SIZE-1:0] Wgt_1_174;input [WEIGHT_SIZE-1:0] Wgt_1_175;input [WEIGHT_SIZE-1:0] Wgt_1_176;input [WEIGHT_SIZE-1:0] Wgt_1_177;input [WEIGHT_SIZE-1:0] Wgt_1_178;input [WEIGHT_SIZE-1:0] Wgt_1_179;input [WEIGHT_SIZE-1:0] Wgt_1_180;input [WEIGHT_SIZE-1:0] Wgt_1_181;input [WEIGHT_SIZE-1:0] Wgt_1_182;input [WEIGHT_SIZE-1:0] Wgt_1_183;input [WEIGHT_SIZE-1:0] Wgt_1_184;input [WEIGHT_SIZE-1:0] Wgt_1_185;input [WEIGHT_SIZE-1:0] Wgt_1_186;input [WEIGHT_SIZE-1:0] Wgt_1_187;input [WEIGHT_SIZE-1:0] Wgt_1_188;input [WEIGHT_SIZE-1:0] Wgt_1_189;input [WEIGHT_SIZE-1:0] Wgt_1_190;input [WEIGHT_SIZE-1:0] Wgt_1_191;input [WEIGHT_SIZE-1:0] Wgt_1_192;input [WEIGHT_SIZE-1:0] Wgt_1_193;input [WEIGHT_SIZE-1:0] Wgt_1_194;input [WEIGHT_SIZE-1:0] Wgt_1_195;input [WEIGHT_SIZE-1:0] Wgt_1_196;input [WEIGHT_SIZE-1:0] Wgt_1_197;input [WEIGHT_SIZE-1:0] Wgt_1_198;input [WEIGHT_SIZE-1:0] Wgt_1_199;input [WEIGHT_SIZE-1:0] Wgt_1_200;input [WEIGHT_SIZE-1:0] Wgt_1_201;input [WEIGHT_SIZE-1:0] Wgt_1_202;input [WEIGHT_SIZE-1:0] Wgt_1_203;input [WEIGHT_SIZE-1:0] Wgt_1_204;input [WEIGHT_SIZE-1:0] Wgt_1_205;input [WEIGHT_SIZE-1:0] Wgt_1_206;input [WEIGHT_SIZE-1:0] Wgt_1_207;input [WEIGHT_SIZE-1:0] Wgt_1_208;input [WEIGHT_SIZE-1:0] Wgt_1_209;input [WEIGHT_SIZE-1:0] Wgt_1_210;input [WEIGHT_SIZE-1:0] Wgt_1_211;input [WEIGHT_SIZE-1:0] Wgt_1_212;input [WEIGHT_SIZE-1:0] Wgt_1_213;input [WEIGHT_SIZE-1:0] Wgt_1_214;input [WEIGHT_SIZE-1:0] Wgt_1_215;input [WEIGHT_SIZE-1:0] Wgt_1_216;input [WEIGHT_SIZE-1:0] Wgt_1_217;input [WEIGHT_SIZE-1:0] Wgt_1_218;input [WEIGHT_SIZE-1:0] Wgt_1_219;input [WEIGHT_SIZE-1:0] Wgt_1_220;input [WEIGHT_SIZE-1:0] Wgt_1_221;input [WEIGHT_SIZE-1:0] Wgt_1_222;input [WEIGHT_SIZE-1:0] Wgt_1_223;input [WEIGHT_SIZE-1:0] Wgt_1_224;input [WEIGHT_SIZE-1:0] Wgt_1_225;input [WEIGHT_SIZE-1:0] Wgt_1_226;input [WEIGHT_SIZE-1:0] Wgt_1_227;input [WEIGHT_SIZE-1:0] Wgt_1_228;input [WEIGHT_SIZE-1:0] Wgt_1_229;input [WEIGHT_SIZE-1:0] Wgt_1_230;input [WEIGHT_SIZE-1:0] Wgt_1_231;input [WEIGHT_SIZE-1:0] Wgt_1_232;input [WEIGHT_SIZE-1:0] Wgt_1_233;input [WEIGHT_SIZE-1:0] Wgt_1_234;input [WEIGHT_SIZE-1:0] Wgt_1_235;input [WEIGHT_SIZE-1:0] Wgt_1_236;input [WEIGHT_SIZE-1:0] Wgt_1_237;input [WEIGHT_SIZE-1:0] Wgt_1_238;input [WEIGHT_SIZE-1:0] Wgt_1_239;input [WEIGHT_SIZE-1:0] Wgt_1_240;input [WEIGHT_SIZE-1:0] Wgt_1_241;input [WEIGHT_SIZE-1:0] Wgt_1_242;input [WEIGHT_SIZE-1:0] Wgt_1_243;input [WEIGHT_SIZE-1:0] Wgt_1_244;input [WEIGHT_SIZE-1:0] Wgt_1_245;input [WEIGHT_SIZE-1:0] Wgt_1_246;input [WEIGHT_SIZE-1:0] Wgt_1_247;input [WEIGHT_SIZE-1:0] Wgt_1_248;input [WEIGHT_SIZE-1:0] Wgt_1_249;input [WEIGHT_SIZE-1:0] Wgt_1_250;input [WEIGHT_SIZE-1:0] Wgt_1_251;input [WEIGHT_SIZE-1:0] Wgt_1_252;input [WEIGHT_SIZE-1:0] Wgt_1_253;input [WEIGHT_SIZE-1:0] Wgt_1_254;input [WEIGHT_SIZE-1:0] Wgt_1_255;input [WEIGHT_SIZE-1:0] Wgt_1_256;input [WEIGHT_SIZE-1:0] Wgt_1_257;input [WEIGHT_SIZE-1:0] Wgt_1_258;input [WEIGHT_SIZE-1:0] Wgt_1_259;input [WEIGHT_SIZE-1:0] Wgt_1_260;input [WEIGHT_SIZE-1:0] Wgt_1_261;input [WEIGHT_SIZE-1:0] Wgt_1_262;input [WEIGHT_SIZE-1:0] Wgt_1_263;input [WEIGHT_SIZE-1:0] Wgt_1_264;input [WEIGHT_SIZE-1:0] Wgt_1_265;input [WEIGHT_SIZE-1:0] Wgt_1_266;input [WEIGHT_SIZE-1:0] Wgt_1_267;input [WEIGHT_SIZE-1:0] Wgt_1_268;input [WEIGHT_SIZE-1:0] Wgt_1_269;input [WEIGHT_SIZE-1:0] Wgt_1_270;input [WEIGHT_SIZE-1:0] Wgt_1_271;input [WEIGHT_SIZE-1:0] Wgt_1_272;input [WEIGHT_SIZE-1:0] Wgt_1_273;input [WEIGHT_SIZE-1:0] Wgt_1_274;input [WEIGHT_SIZE-1:0] Wgt_1_275;input [WEIGHT_SIZE-1:0] Wgt_1_276;input [WEIGHT_SIZE-1:0] Wgt_1_277;input [WEIGHT_SIZE-1:0] Wgt_1_278;input [WEIGHT_SIZE-1:0] Wgt_1_279;input [WEIGHT_SIZE-1:0] Wgt_1_280;input [WEIGHT_SIZE-1:0] Wgt_1_281;input [WEIGHT_SIZE-1:0] Wgt_1_282;input [WEIGHT_SIZE-1:0] Wgt_1_283;input [WEIGHT_SIZE-1:0] Wgt_1_284;input [WEIGHT_SIZE-1:0] Wgt_1_285;input [WEIGHT_SIZE-1:0] Wgt_1_286;input [WEIGHT_SIZE-1:0] Wgt_1_287;input [WEIGHT_SIZE-1:0] Wgt_1_288;input [WEIGHT_SIZE-1:0] Wgt_1_289;input [WEIGHT_SIZE-1:0] Wgt_1_290;input [WEIGHT_SIZE-1:0] Wgt_1_291;input [WEIGHT_SIZE-1:0] Wgt_1_292;input [WEIGHT_SIZE-1:0] Wgt_1_293;input [WEIGHT_SIZE-1:0] Wgt_1_294;input [WEIGHT_SIZE-1:0] Wgt_1_295;input [WEIGHT_SIZE-1:0] Wgt_1_296;input [WEIGHT_SIZE-1:0] Wgt_1_297;input [WEIGHT_SIZE-1:0] Wgt_1_298;input [WEIGHT_SIZE-1:0] Wgt_1_299;input [WEIGHT_SIZE-1:0] Wgt_1_300;input [WEIGHT_SIZE-1:0] Wgt_1_301;input [WEIGHT_SIZE-1:0] Wgt_1_302;input [WEIGHT_SIZE-1:0] Wgt_1_303;input [WEIGHT_SIZE-1:0] Wgt_1_304;input [WEIGHT_SIZE-1:0] Wgt_1_305;input [WEIGHT_SIZE-1:0] Wgt_1_306;input [WEIGHT_SIZE-1:0] Wgt_1_307;input [WEIGHT_SIZE-1:0] Wgt_1_308;input [WEIGHT_SIZE-1:0] Wgt_1_309;input [WEIGHT_SIZE-1:0] Wgt_1_310;input [WEIGHT_SIZE-1:0] Wgt_1_311;input [WEIGHT_SIZE-1:0] Wgt_1_312;input [WEIGHT_SIZE-1:0] Wgt_1_313;input [WEIGHT_SIZE-1:0] Wgt_1_314;input [WEIGHT_SIZE-1:0] Wgt_1_315;input [WEIGHT_SIZE-1:0] Wgt_1_316;input [WEIGHT_SIZE-1:0] Wgt_1_317;input [WEIGHT_SIZE-1:0] Wgt_1_318;input [WEIGHT_SIZE-1:0] Wgt_1_319;input [WEIGHT_SIZE-1:0] Wgt_1_320;input [WEIGHT_SIZE-1:0] Wgt_1_321;input [WEIGHT_SIZE-1:0] Wgt_1_322;input [WEIGHT_SIZE-1:0] Wgt_1_323;input [WEIGHT_SIZE-1:0] Wgt_1_324;input [WEIGHT_SIZE-1:0] Wgt_1_325;input [WEIGHT_SIZE-1:0] Wgt_1_326;input [WEIGHT_SIZE-1:0] Wgt_1_327;input [WEIGHT_SIZE-1:0] Wgt_1_328;input [WEIGHT_SIZE-1:0] Wgt_1_329;input [WEIGHT_SIZE-1:0] Wgt_1_330;input [WEIGHT_SIZE-1:0] Wgt_1_331;input [WEIGHT_SIZE-1:0] Wgt_1_332;input [WEIGHT_SIZE-1:0] Wgt_1_333;input [WEIGHT_SIZE-1:0] Wgt_1_334;input [WEIGHT_SIZE-1:0] Wgt_1_335;input [WEIGHT_SIZE-1:0] Wgt_1_336;input [WEIGHT_SIZE-1:0] Wgt_1_337;input [WEIGHT_SIZE-1:0] Wgt_1_338;input [WEIGHT_SIZE-1:0] Wgt_1_339;input [WEIGHT_SIZE-1:0] Wgt_1_340;input [WEIGHT_SIZE-1:0] Wgt_1_341;input [WEIGHT_SIZE-1:0] Wgt_1_342;input [WEIGHT_SIZE-1:0] Wgt_1_343;input [WEIGHT_SIZE-1:0] Wgt_1_344;input [WEIGHT_SIZE-1:0] Wgt_1_345;input [WEIGHT_SIZE-1:0] Wgt_1_346;input [WEIGHT_SIZE-1:0] Wgt_1_347;input [WEIGHT_SIZE-1:0] Wgt_1_348;input [WEIGHT_SIZE-1:0] Wgt_1_349;input [WEIGHT_SIZE-1:0] Wgt_1_350;input [WEIGHT_SIZE-1:0] Wgt_1_351;input [WEIGHT_SIZE-1:0] Wgt_1_352;input [WEIGHT_SIZE-1:0] Wgt_1_353;input [WEIGHT_SIZE-1:0] Wgt_1_354;input [WEIGHT_SIZE-1:0] Wgt_1_355;input [WEIGHT_SIZE-1:0] Wgt_1_356;input [WEIGHT_SIZE-1:0] Wgt_1_357;input [WEIGHT_SIZE-1:0] Wgt_1_358;input [WEIGHT_SIZE-1:0] Wgt_1_359;input [WEIGHT_SIZE-1:0] Wgt_1_360;input [WEIGHT_SIZE-1:0] Wgt_1_361;input [WEIGHT_SIZE-1:0] Wgt_1_362;input [WEIGHT_SIZE-1:0] Wgt_1_363;input [WEIGHT_SIZE-1:0] Wgt_1_364;input [WEIGHT_SIZE-1:0] Wgt_1_365;input [WEIGHT_SIZE-1:0] Wgt_1_366;input [WEIGHT_SIZE-1:0] Wgt_1_367;input [WEIGHT_SIZE-1:0] Wgt_1_368;input [WEIGHT_SIZE-1:0] Wgt_1_369;input [WEIGHT_SIZE-1:0] Wgt_1_370;input [WEIGHT_SIZE-1:0] Wgt_1_371;input [WEIGHT_SIZE-1:0] Wgt_1_372;input [WEIGHT_SIZE-1:0] Wgt_1_373;input [WEIGHT_SIZE-1:0] Wgt_1_374;input [WEIGHT_SIZE-1:0] Wgt_1_375;input [WEIGHT_SIZE-1:0] Wgt_1_376;input [WEIGHT_SIZE-1:0] Wgt_1_377;input [WEIGHT_SIZE-1:0] Wgt_1_378;input [WEIGHT_SIZE-1:0] Wgt_1_379;input [WEIGHT_SIZE-1:0] Wgt_1_380;input [WEIGHT_SIZE-1:0] Wgt_1_381;input [WEIGHT_SIZE-1:0] Wgt_1_382;input [WEIGHT_SIZE-1:0] Wgt_1_383;input [WEIGHT_SIZE-1:0] Wgt_1_384;input [WEIGHT_SIZE-1:0] Wgt_1_385;input [WEIGHT_SIZE-1:0] Wgt_1_386;input [WEIGHT_SIZE-1:0] Wgt_1_387;input [WEIGHT_SIZE-1:0] Wgt_1_388;input [WEIGHT_SIZE-1:0] Wgt_1_389;input [WEIGHT_SIZE-1:0] Wgt_1_390;input [WEIGHT_SIZE-1:0] Wgt_1_391;input [WEIGHT_SIZE-1:0] Wgt_1_392;input [WEIGHT_SIZE-1:0] Wgt_1_393;input [WEIGHT_SIZE-1:0] Wgt_1_394;input [WEIGHT_SIZE-1:0] Wgt_1_395;input [WEIGHT_SIZE-1:0] Wgt_1_396;input [WEIGHT_SIZE-1:0] Wgt_1_397;input [WEIGHT_SIZE-1:0] Wgt_1_398;input [WEIGHT_SIZE-1:0] Wgt_1_399;input [WEIGHT_SIZE-1:0] Wgt_1_400;input [WEIGHT_SIZE-1:0] Wgt_1_401;input [WEIGHT_SIZE-1:0] Wgt_1_402;input [WEIGHT_SIZE-1:0] Wgt_1_403;input [WEIGHT_SIZE-1:0] Wgt_1_404;input [WEIGHT_SIZE-1:0] Wgt_1_405;input [WEIGHT_SIZE-1:0] Wgt_1_406;input [WEIGHT_SIZE-1:0] Wgt_1_407;input [WEIGHT_SIZE-1:0] Wgt_1_408;input [WEIGHT_SIZE-1:0] Wgt_1_409;input [WEIGHT_SIZE-1:0] Wgt_1_410;input [WEIGHT_SIZE-1:0] Wgt_1_411;input [WEIGHT_SIZE-1:0] Wgt_1_412;input [WEIGHT_SIZE-1:0] Wgt_1_413;input [WEIGHT_SIZE-1:0] Wgt_1_414;input [WEIGHT_SIZE-1:0] Wgt_1_415;input [WEIGHT_SIZE-1:0] Wgt_1_416;input [WEIGHT_SIZE-1:0] Wgt_1_417;input [WEIGHT_SIZE-1:0] Wgt_1_418;input [WEIGHT_SIZE-1:0] Wgt_1_419;input [WEIGHT_SIZE-1:0] Wgt_1_420;input [WEIGHT_SIZE-1:0] Wgt_1_421;input [WEIGHT_SIZE-1:0] Wgt_1_422;input [WEIGHT_SIZE-1:0] Wgt_1_423;input [WEIGHT_SIZE-1:0] Wgt_1_424;input [WEIGHT_SIZE-1:0] Wgt_1_425;input [WEIGHT_SIZE-1:0] Wgt_1_426;input [WEIGHT_SIZE-1:0] Wgt_1_427;input [WEIGHT_SIZE-1:0] Wgt_1_428;input [WEIGHT_SIZE-1:0] Wgt_1_429;input [WEIGHT_SIZE-1:0] Wgt_1_430;input [WEIGHT_SIZE-1:0] Wgt_1_431;input [WEIGHT_SIZE-1:0] Wgt_1_432;input [WEIGHT_SIZE-1:0] Wgt_1_433;input [WEIGHT_SIZE-1:0] Wgt_1_434;input [WEIGHT_SIZE-1:0] Wgt_1_435;input [WEIGHT_SIZE-1:0] Wgt_1_436;input [WEIGHT_SIZE-1:0] Wgt_1_437;input [WEIGHT_SIZE-1:0] Wgt_1_438;input [WEIGHT_SIZE-1:0] Wgt_1_439;input [WEIGHT_SIZE-1:0] Wgt_1_440;input [WEIGHT_SIZE-1:0] Wgt_1_441;input [WEIGHT_SIZE-1:0] Wgt_1_442;input [WEIGHT_SIZE-1:0] Wgt_1_443;input [WEIGHT_SIZE-1:0] Wgt_1_444;input [WEIGHT_SIZE-1:0] Wgt_1_445;input [WEIGHT_SIZE-1:0] Wgt_1_446;input [WEIGHT_SIZE-1:0] Wgt_1_447;input [WEIGHT_SIZE-1:0] Wgt_1_448;input [WEIGHT_SIZE-1:0] Wgt_1_449;input [WEIGHT_SIZE-1:0] Wgt_1_450;input [WEIGHT_SIZE-1:0] Wgt_1_451;input [WEIGHT_SIZE-1:0] Wgt_1_452;input [WEIGHT_SIZE-1:0] Wgt_1_453;input [WEIGHT_SIZE-1:0] Wgt_1_454;input [WEIGHT_SIZE-1:0] Wgt_1_455;input [WEIGHT_SIZE-1:0] Wgt_1_456;input [WEIGHT_SIZE-1:0] Wgt_1_457;input [WEIGHT_SIZE-1:0] Wgt_1_458;input [WEIGHT_SIZE-1:0] Wgt_1_459;input [WEIGHT_SIZE-1:0] Wgt_1_460;input [WEIGHT_SIZE-1:0] Wgt_1_461;input [WEIGHT_SIZE-1:0] Wgt_1_462;input [WEIGHT_SIZE-1:0] Wgt_1_463;input [WEIGHT_SIZE-1:0] Wgt_1_464;input [WEIGHT_SIZE-1:0] Wgt_1_465;input [WEIGHT_SIZE-1:0] Wgt_1_466;input [WEIGHT_SIZE-1:0] Wgt_1_467;input [WEIGHT_SIZE-1:0] Wgt_1_468;input [WEIGHT_SIZE-1:0] Wgt_1_469;input [WEIGHT_SIZE-1:0] Wgt_1_470;input [WEIGHT_SIZE-1:0] Wgt_1_471;input [WEIGHT_SIZE-1:0] Wgt_1_472;input [WEIGHT_SIZE-1:0] Wgt_1_473;input [WEIGHT_SIZE-1:0] Wgt_1_474;input [WEIGHT_SIZE-1:0] Wgt_1_475;input [WEIGHT_SIZE-1:0] Wgt_1_476;input [WEIGHT_SIZE-1:0] Wgt_1_477;input [WEIGHT_SIZE-1:0] Wgt_1_478;input [WEIGHT_SIZE-1:0] Wgt_1_479;input [WEIGHT_SIZE-1:0] Wgt_1_480;input [WEIGHT_SIZE-1:0] Wgt_1_481;input [WEIGHT_SIZE-1:0] Wgt_1_482;input [WEIGHT_SIZE-1:0] Wgt_1_483;input [WEIGHT_SIZE-1:0] Wgt_1_484;input [WEIGHT_SIZE-1:0] Wgt_1_485;input [WEIGHT_SIZE-1:0] Wgt_1_486;input [WEIGHT_SIZE-1:0] Wgt_1_487;input [WEIGHT_SIZE-1:0] Wgt_1_488;input [WEIGHT_SIZE-1:0] Wgt_1_489;input [WEIGHT_SIZE-1:0] Wgt_1_490;input [WEIGHT_SIZE-1:0] Wgt_1_491;input [WEIGHT_SIZE-1:0] Wgt_1_492;input [WEIGHT_SIZE-1:0] Wgt_1_493;input [WEIGHT_SIZE-1:0] Wgt_1_494;input [WEIGHT_SIZE-1:0] Wgt_1_495;input [WEIGHT_SIZE-1:0] Wgt_1_496;input [WEIGHT_SIZE-1:0] Wgt_1_497;input [WEIGHT_SIZE-1:0] Wgt_1_498;input [WEIGHT_SIZE-1:0] Wgt_1_499;input [WEIGHT_SIZE-1:0] Wgt_1_500;input [WEIGHT_SIZE-1:0] Wgt_1_501;input [WEIGHT_SIZE-1:0] Wgt_1_502;input [WEIGHT_SIZE-1:0] Wgt_1_503;input [WEIGHT_SIZE-1:0] Wgt_1_504;input [WEIGHT_SIZE-1:0] Wgt_1_505;input [WEIGHT_SIZE-1:0] Wgt_1_506;input [WEIGHT_SIZE-1:0] Wgt_1_507;input [WEIGHT_SIZE-1:0] Wgt_1_508;input [WEIGHT_SIZE-1:0] Wgt_1_509;input [WEIGHT_SIZE-1:0] Wgt_1_510;input [WEIGHT_SIZE-1:0] Wgt_1_511;input [WEIGHT_SIZE-1:0] Wgt_1_512;input [WEIGHT_SIZE-1:0] Wgt_1_513;input [WEIGHT_SIZE-1:0] Wgt_1_514;input [WEIGHT_SIZE-1:0] Wgt_1_515;input [WEIGHT_SIZE-1:0] Wgt_1_516;input [WEIGHT_SIZE-1:0] Wgt_1_517;input [WEIGHT_SIZE-1:0] Wgt_1_518;input [WEIGHT_SIZE-1:0] Wgt_1_519;input [WEIGHT_SIZE-1:0] Wgt_1_520;input [WEIGHT_SIZE-1:0] Wgt_1_521;input [WEIGHT_SIZE-1:0] Wgt_1_522;input [WEIGHT_SIZE-1:0] Wgt_1_523;input [WEIGHT_SIZE-1:0] Wgt_1_524;input [WEIGHT_SIZE-1:0] Wgt_1_525;input [WEIGHT_SIZE-1:0] Wgt_1_526;input [WEIGHT_SIZE-1:0] Wgt_1_527;input [WEIGHT_SIZE-1:0] Wgt_1_528;input [WEIGHT_SIZE-1:0] Wgt_1_529;input [WEIGHT_SIZE-1:0] Wgt_1_530;input [WEIGHT_SIZE-1:0] Wgt_1_531;input [WEIGHT_SIZE-1:0] Wgt_1_532;input [WEIGHT_SIZE-1:0] Wgt_1_533;input [WEIGHT_SIZE-1:0] Wgt_1_534;input [WEIGHT_SIZE-1:0] Wgt_1_535;input [WEIGHT_SIZE-1:0] Wgt_1_536;input [WEIGHT_SIZE-1:0] Wgt_1_537;input [WEIGHT_SIZE-1:0] Wgt_1_538;input [WEIGHT_SIZE-1:0] Wgt_1_539;input [WEIGHT_SIZE-1:0] Wgt_1_540;input [WEIGHT_SIZE-1:0] Wgt_1_541;input [WEIGHT_SIZE-1:0] Wgt_1_542;input [WEIGHT_SIZE-1:0] Wgt_1_543;input [WEIGHT_SIZE-1:0] Wgt_1_544;input [WEIGHT_SIZE-1:0] Wgt_1_545;input [WEIGHT_SIZE-1:0] Wgt_1_546;input [WEIGHT_SIZE-1:0] Wgt_1_547;input [WEIGHT_SIZE-1:0] Wgt_1_548;input [WEIGHT_SIZE-1:0] Wgt_1_549;input [WEIGHT_SIZE-1:0] Wgt_1_550;input [WEIGHT_SIZE-1:0] Wgt_1_551;input [WEIGHT_SIZE-1:0] Wgt_1_552;input [WEIGHT_SIZE-1:0] Wgt_1_553;input [WEIGHT_SIZE-1:0] Wgt_1_554;input [WEIGHT_SIZE-1:0] Wgt_1_555;input [WEIGHT_SIZE-1:0] Wgt_1_556;input [WEIGHT_SIZE-1:0] Wgt_1_557;input [WEIGHT_SIZE-1:0] Wgt_1_558;input [WEIGHT_SIZE-1:0] Wgt_1_559;input [WEIGHT_SIZE-1:0] Wgt_1_560;input [WEIGHT_SIZE-1:0] Wgt_1_561;input [WEIGHT_SIZE-1:0] Wgt_1_562;input [WEIGHT_SIZE-1:0] Wgt_1_563;input [WEIGHT_SIZE-1:0] Wgt_1_564;input [WEIGHT_SIZE-1:0] Wgt_1_565;input [WEIGHT_SIZE-1:0] Wgt_1_566;input [WEIGHT_SIZE-1:0] Wgt_1_567;input [WEIGHT_SIZE-1:0] Wgt_1_568;input [WEIGHT_SIZE-1:0] Wgt_1_569;input [WEIGHT_SIZE-1:0] Wgt_1_570;input [WEIGHT_SIZE-1:0] Wgt_1_571;input [WEIGHT_SIZE-1:0] Wgt_1_572;input [WEIGHT_SIZE-1:0] Wgt_1_573;input [WEIGHT_SIZE-1:0] Wgt_1_574;input [WEIGHT_SIZE-1:0] Wgt_1_575;input [WEIGHT_SIZE-1:0] Wgt_1_576;input [WEIGHT_SIZE-1:0] Wgt_1_577;input [WEIGHT_SIZE-1:0] Wgt_1_578;input [WEIGHT_SIZE-1:0] Wgt_1_579;input [WEIGHT_SIZE-1:0] Wgt_1_580;input [WEIGHT_SIZE-1:0] Wgt_1_581;input [WEIGHT_SIZE-1:0] Wgt_1_582;input [WEIGHT_SIZE-1:0] Wgt_1_583;input [WEIGHT_SIZE-1:0] Wgt_1_584;input [WEIGHT_SIZE-1:0] Wgt_1_585;input [WEIGHT_SIZE-1:0] Wgt_1_586;input [WEIGHT_SIZE-1:0] Wgt_1_587;input [WEIGHT_SIZE-1:0] Wgt_1_588;input [WEIGHT_SIZE-1:0] Wgt_1_589;input [WEIGHT_SIZE-1:0] Wgt_1_590;input [WEIGHT_SIZE-1:0] Wgt_1_591;input [WEIGHT_SIZE-1:0] Wgt_1_592;input [WEIGHT_SIZE-1:0] Wgt_1_593;input [WEIGHT_SIZE-1:0] Wgt_1_594;input [WEIGHT_SIZE-1:0] Wgt_1_595;input [WEIGHT_SIZE-1:0] Wgt_1_596;input [WEIGHT_SIZE-1:0] Wgt_1_597;input [WEIGHT_SIZE-1:0] Wgt_1_598;input [WEIGHT_SIZE-1:0] Wgt_1_599;input [WEIGHT_SIZE-1:0] Wgt_1_600;input [WEIGHT_SIZE-1:0] Wgt_1_601;input [WEIGHT_SIZE-1:0] Wgt_1_602;input [WEIGHT_SIZE-1:0] Wgt_1_603;input [WEIGHT_SIZE-1:0] Wgt_1_604;input [WEIGHT_SIZE-1:0] Wgt_1_605;input [WEIGHT_SIZE-1:0] Wgt_1_606;input [WEIGHT_SIZE-1:0] Wgt_1_607;input [WEIGHT_SIZE-1:0] Wgt_1_608;input [WEIGHT_SIZE-1:0] Wgt_1_609;input [WEIGHT_SIZE-1:0] Wgt_1_610;input [WEIGHT_SIZE-1:0] Wgt_1_611;input [WEIGHT_SIZE-1:0] Wgt_1_612;input [WEIGHT_SIZE-1:0] Wgt_1_613;input [WEIGHT_SIZE-1:0] Wgt_1_614;input [WEIGHT_SIZE-1:0] Wgt_1_615;input [WEIGHT_SIZE-1:0] Wgt_1_616;input [WEIGHT_SIZE-1:0] Wgt_1_617;input [WEIGHT_SIZE-1:0] Wgt_1_618;input [WEIGHT_SIZE-1:0] Wgt_1_619;input [WEIGHT_SIZE-1:0] Wgt_1_620;input [WEIGHT_SIZE-1:0] Wgt_1_621;input [WEIGHT_SIZE-1:0] Wgt_1_622;input [WEIGHT_SIZE-1:0] Wgt_1_623;input [WEIGHT_SIZE-1:0] Wgt_1_624;input [WEIGHT_SIZE-1:0] Wgt_1_625;input [WEIGHT_SIZE-1:0] Wgt_1_626;input [WEIGHT_SIZE-1:0] Wgt_1_627;input [WEIGHT_SIZE-1:0] Wgt_1_628;input [WEIGHT_SIZE-1:0] Wgt_1_629;input [WEIGHT_SIZE-1:0] Wgt_1_630;input [WEIGHT_SIZE-1:0] Wgt_1_631;input [WEIGHT_SIZE-1:0] Wgt_1_632;input [WEIGHT_SIZE-1:0] Wgt_1_633;input [WEIGHT_SIZE-1:0] Wgt_1_634;input [WEIGHT_SIZE-1:0] Wgt_1_635;input [WEIGHT_SIZE-1:0] Wgt_1_636;input [WEIGHT_SIZE-1:0] Wgt_1_637;input [WEIGHT_SIZE-1:0] Wgt_1_638;input [WEIGHT_SIZE-1:0] Wgt_1_639;input [WEIGHT_SIZE-1:0] Wgt_1_640;input [WEIGHT_SIZE-1:0] Wgt_1_641;input [WEIGHT_SIZE-1:0] Wgt_1_642;input [WEIGHT_SIZE-1:0] Wgt_1_643;input [WEIGHT_SIZE-1:0] Wgt_1_644;input [WEIGHT_SIZE-1:0] Wgt_1_645;input [WEIGHT_SIZE-1:0] Wgt_1_646;input [WEIGHT_SIZE-1:0] Wgt_1_647;input [WEIGHT_SIZE-1:0] Wgt_1_648;input [WEIGHT_SIZE-1:0] Wgt_1_649;input [WEIGHT_SIZE-1:0] Wgt_1_650;input [WEIGHT_SIZE-1:0] Wgt_1_651;input [WEIGHT_SIZE-1:0] Wgt_1_652;input [WEIGHT_SIZE-1:0] Wgt_1_653;input [WEIGHT_SIZE-1:0] Wgt_1_654;input [WEIGHT_SIZE-1:0] Wgt_1_655;input [WEIGHT_SIZE-1:0] Wgt_1_656;input [WEIGHT_SIZE-1:0] Wgt_1_657;input [WEIGHT_SIZE-1:0] Wgt_1_658;input [WEIGHT_SIZE-1:0] Wgt_1_659;input [WEIGHT_SIZE-1:0] Wgt_1_660;input [WEIGHT_SIZE-1:0] Wgt_1_661;input [WEIGHT_SIZE-1:0] Wgt_1_662;input [WEIGHT_SIZE-1:0] Wgt_1_663;input [WEIGHT_SIZE-1:0] Wgt_1_664;input [WEIGHT_SIZE-1:0] Wgt_1_665;input [WEIGHT_SIZE-1:0] Wgt_1_666;input [WEIGHT_SIZE-1:0] Wgt_1_667;input [WEIGHT_SIZE-1:0] Wgt_1_668;input [WEIGHT_SIZE-1:0] Wgt_1_669;input [WEIGHT_SIZE-1:0] Wgt_1_670;input [WEIGHT_SIZE-1:0] Wgt_1_671;input [WEIGHT_SIZE-1:0] Wgt_1_672;input [WEIGHT_SIZE-1:0] Wgt_1_673;input [WEIGHT_SIZE-1:0] Wgt_1_674;input [WEIGHT_SIZE-1:0] Wgt_1_675;input [WEIGHT_SIZE-1:0] Wgt_1_676;input [WEIGHT_SIZE-1:0] Wgt_1_677;input [WEIGHT_SIZE-1:0] Wgt_1_678;input [WEIGHT_SIZE-1:0] Wgt_1_679;input [WEIGHT_SIZE-1:0] Wgt_1_680;input [WEIGHT_SIZE-1:0] Wgt_1_681;input [WEIGHT_SIZE-1:0] Wgt_1_682;input [WEIGHT_SIZE-1:0] Wgt_1_683;input [WEIGHT_SIZE-1:0] Wgt_1_684;input [WEIGHT_SIZE-1:0] Wgt_1_685;input [WEIGHT_SIZE-1:0] Wgt_1_686;input [WEIGHT_SIZE-1:0] Wgt_1_687;input [WEIGHT_SIZE-1:0] Wgt_1_688;input [WEIGHT_SIZE-1:0] Wgt_1_689;input [WEIGHT_SIZE-1:0] Wgt_1_690;input [WEIGHT_SIZE-1:0] Wgt_1_691;input [WEIGHT_SIZE-1:0] Wgt_1_692;input [WEIGHT_SIZE-1:0] Wgt_1_693;input [WEIGHT_SIZE-1:0] Wgt_1_694;input [WEIGHT_SIZE-1:0] Wgt_1_695;input [WEIGHT_SIZE-1:0] Wgt_1_696;input [WEIGHT_SIZE-1:0] Wgt_1_697;input [WEIGHT_SIZE-1:0] Wgt_1_698;input [WEIGHT_SIZE-1:0] Wgt_1_699;input [WEIGHT_SIZE-1:0] Wgt_1_700;input [WEIGHT_SIZE-1:0] Wgt_1_701;input [WEIGHT_SIZE-1:0] Wgt_1_702;input [WEIGHT_SIZE-1:0] Wgt_1_703;input [WEIGHT_SIZE-1:0] Wgt_1_704;input [WEIGHT_SIZE-1:0] Wgt_1_705;input [WEIGHT_SIZE-1:0] Wgt_1_706;input [WEIGHT_SIZE-1:0] Wgt_1_707;input [WEIGHT_SIZE-1:0] Wgt_1_708;input [WEIGHT_SIZE-1:0] Wgt_1_709;input [WEIGHT_SIZE-1:0] Wgt_1_710;input [WEIGHT_SIZE-1:0] Wgt_1_711;input [WEIGHT_SIZE-1:0] Wgt_1_712;input [WEIGHT_SIZE-1:0] Wgt_1_713;input [WEIGHT_SIZE-1:0] Wgt_1_714;input [WEIGHT_SIZE-1:0] Wgt_1_715;input [WEIGHT_SIZE-1:0] Wgt_1_716;input [WEIGHT_SIZE-1:0] Wgt_1_717;input [WEIGHT_SIZE-1:0] Wgt_1_718;input [WEIGHT_SIZE-1:0] Wgt_1_719;input [WEIGHT_SIZE-1:0] Wgt_1_720;input [WEIGHT_SIZE-1:0] Wgt_1_721;input [WEIGHT_SIZE-1:0] Wgt_1_722;input [WEIGHT_SIZE-1:0] Wgt_1_723;input [WEIGHT_SIZE-1:0] Wgt_1_724;input [WEIGHT_SIZE-1:0] Wgt_1_725;input [WEIGHT_SIZE-1:0] Wgt_1_726;input [WEIGHT_SIZE-1:0] Wgt_1_727;input [WEIGHT_SIZE-1:0] Wgt_1_728;input [WEIGHT_SIZE-1:0] Wgt_1_729;input [WEIGHT_SIZE-1:0] Wgt_1_730;input [WEIGHT_SIZE-1:0] Wgt_1_731;input [WEIGHT_SIZE-1:0] Wgt_1_732;input [WEIGHT_SIZE-1:0] Wgt_1_733;input [WEIGHT_SIZE-1:0] Wgt_1_734;input [WEIGHT_SIZE-1:0] Wgt_1_735;input [WEIGHT_SIZE-1:0] Wgt_1_736;input [WEIGHT_SIZE-1:0] Wgt_1_737;input [WEIGHT_SIZE-1:0] Wgt_1_738;input [WEIGHT_SIZE-1:0] Wgt_1_739;input [WEIGHT_SIZE-1:0] Wgt_1_740;input [WEIGHT_SIZE-1:0] Wgt_1_741;input [WEIGHT_SIZE-1:0] Wgt_1_742;input [WEIGHT_SIZE-1:0] Wgt_1_743;input [WEIGHT_SIZE-1:0] Wgt_1_744;input [WEIGHT_SIZE-1:0] Wgt_1_745;input [WEIGHT_SIZE-1:0] Wgt_1_746;input [WEIGHT_SIZE-1:0] Wgt_1_747;input [WEIGHT_SIZE-1:0] Wgt_1_748;input [WEIGHT_SIZE-1:0] Wgt_1_749;input [WEIGHT_SIZE-1:0] Wgt_1_750;input [WEIGHT_SIZE-1:0] Wgt_1_751;input [WEIGHT_SIZE-1:0] Wgt_1_752;input [WEIGHT_SIZE-1:0] Wgt_1_753;input [WEIGHT_SIZE-1:0] Wgt_1_754;input [WEIGHT_SIZE-1:0] Wgt_1_755;input [WEIGHT_SIZE-1:0] Wgt_1_756;input [WEIGHT_SIZE-1:0] Wgt_1_757;input [WEIGHT_SIZE-1:0] Wgt_1_758;input [WEIGHT_SIZE-1:0] Wgt_1_759;input [WEIGHT_SIZE-1:0] Wgt_1_760;input [WEIGHT_SIZE-1:0] Wgt_1_761;input [WEIGHT_SIZE-1:0] Wgt_1_762;input [WEIGHT_SIZE-1:0] Wgt_1_763;input [WEIGHT_SIZE-1:0] Wgt_1_764;input [WEIGHT_SIZE-1:0] Wgt_1_765;input [WEIGHT_SIZE-1:0] Wgt_1_766;input [WEIGHT_SIZE-1:0] Wgt_1_767;input [WEIGHT_SIZE-1:0] Wgt_1_768;input [WEIGHT_SIZE-1:0] Wgt_1_769;input [WEIGHT_SIZE-1:0] Wgt_1_770;input [WEIGHT_SIZE-1:0] Wgt_1_771;input [WEIGHT_SIZE-1:0] Wgt_1_772;input [WEIGHT_SIZE-1:0] Wgt_1_773;input [WEIGHT_SIZE-1:0] Wgt_1_774;input [WEIGHT_SIZE-1:0] Wgt_1_775;input [WEIGHT_SIZE-1:0] Wgt_1_776;input [WEIGHT_SIZE-1:0] Wgt_1_777;input [WEIGHT_SIZE-1:0] Wgt_1_778;input [WEIGHT_SIZE-1:0] Wgt_1_779;input [WEIGHT_SIZE-1:0] Wgt_1_780;input [WEIGHT_SIZE-1:0] Wgt_1_781;input [WEIGHT_SIZE-1:0] Wgt_1_782;input [WEIGHT_SIZE-1:0] Wgt_1_783;input [WEIGHT_SIZE-1:0] Wgt_1_784;input [WEIGHT_SIZE-1:0] Wgt_2_0;input [WEIGHT_SIZE-1:0] Wgt_2_1;input [WEIGHT_SIZE-1:0] Wgt_2_2;input [WEIGHT_SIZE-1:0] Wgt_2_3;input [WEIGHT_SIZE-1:0] Wgt_2_4;input [WEIGHT_SIZE-1:0] Wgt_2_5;input [WEIGHT_SIZE-1:0] Wgt_2_6;input [WEIGHT_SIZE-1:0] Wgt_2_7;input [WEIGHT_SIZE-1:0] Wgt_2_8;input [WEIGHT_SIZE-1:0] Wgt_2_9;input [WEIGHT_SIZE-1:0] Wgt_2_10;input [WEIGHT_SIZE-1:0] Wgt_2_11;input [WEIGHT_SIZE-1:0] Wgt_2_12;input [WEIGHT_SIZE-1:0] Wgt_2_13;input [WEIGHT_SIZE-1:0] Wgt_2_14;input [WEIGHT_SIZE-1:0] Wgt_2_15;input [WEIGHT_SIZE-1:0] Wgt_2_16;input [WEIGHT_SIZE-1:0] Wgt_2_17;input [WEIGHT_SIZE-1:0] Wgt_2_18;input [WEIGHT_SIZE-1:0] Wgt_2_19;input [WEIGHT_SIZE-1:0] Wgt_2_20;input [WEIGHT_SIZE-1:0] Wgt_2_21;input [WEIGHT_SIZE-1:0] Wgt_2_22;input [WEIGHT_SIZE-1:0] Wgt_2_23;input [WEIGHT_SIZE-1:0] Wgt_2_24;input [WEIGHT_SIZE-1:0] Wgt_2_25;input [WEIGHT_SIZE-1:0] Wgt_2_26;input [WEIGHT_SIZE-1:0] Wgt_2_27;input [WEIGHT_SIZE-1:0] Wgt_2_28;input [WEIGHT_SIZE-1:0] Wgt_2_29;input [WEIGHT_SIZE-1:0] Wgt_2_30;input [WEIGHT_SIZE-1:0] Wgt_2_31;input [WEIGHT_SIZE-1:0] Wgt_2_32;input [WEIGHT_SIZE-1:0] Wgt_2_33;input [WEIGHT_SIZE-1:0] Wgt_2_34;input [WEIGHT_SIZE-1:0] Wgt_2_35;input [WEIGHT_SIZE-1:0] Wgt_2_36;input [WEIGHT_SIZE-1:0] Wgt_2_37;input [WEIGHT_SIZE-1:0] Wgt_2_38;input [WEIGHT_SIZE-1:0] Wgt_2_39;input [WEIGHT_SIZE-1:0] Wgt_2_40;input [WEIGHT_SIZE-1:0] Wgt_2_41;input [WEIGHT_SIZE-1:0] Wgt_2_42;input [WEIGHT_SIZE-1:0] Wgt_2_43;input [WEIGHT_SIZE-1:0] Wgt_2_44;input [WEIGHT_SIZE-1:0] Wgt_2_45;input [WEIGHT_SIZE-1:0] Wgt_2_46;input [WEIGHT_SIZE-1:0] Wgt_2_47;input [WEIGHT_SIZE-1:0] Wgt_2_48;input [WEIGHT_SIZE-1:0] Wgt_2_49;input [WEIGHT_SIZE-1:0] Wgt_2_50;input [WEIGHT_SIZE-1:0] Wgt_2_51;input [WEIGHT_SIZE-1:0] Wgt_2_52;input [WEIGHT_SIZE-1:0] Wgt_2_53;input [WEIGHT_SIZE-1:0] Wgt_2_54;input [WEIGHT_SIZE-1:0] Wgt_2_55;input [WEIGHT_SIZE-1:0] Wgt_2_56;input [WEIGHT_SIZE-1:0] Wgt_2_57;input [WEIGHT_SIZE-1:0] Wgt_2_58;input [WEIGHT_SIZE-1:0] Wgt_2_59;input [WEIGHT_SIZE-1:0] Wgt_2_60;input [WEIGHT_SIZE-1:0] Wgt_2_61;input [WEIGHT_SIZE-1:0] Wgt_2_62;input [WEIGHT_SIZE-1:0] Wgt_2_63;input [WEIGHT_SIZE-1:0] Wgt_2_64;input [WEIGHT_SIZE-1:0] Wgt_2_65;input [WEIGHT_SIZE-1:0] Wgt_2_66;input [WEIGHT_SIZE-1:0] Wgt_2_67;input [WEIGHT_SIZE-1:0] Wgt_2_68;input [WEIGHT_SIZE-1:0] Wgt_2_69;input [WEIGHT_SIZE-1:0] Wgt_2_70;input [WEIGHT_SIZE-1:0] Wgt_2_71;input [WEIGHT_SIZE-1:0] Wgt_2_72;input [WEIGHT_SIZE-1:0] Wgt_2_73;input [WEIGHT_SIZE-1:0] Wgt_2_74;input [WEIGHT_SIZE-1:0] Wgt_2_75;input [WEIGHT_SIZE-1:0] Wgt_2_76;input [WEIGHT_SIZE-1:0] Wgt_2_77;input [WEIGHT_SIZE-1:0] Wgt_2_78;input [WEIGHT_SIZE-1:0] Wgt_2_79;input [WEIGHT_SIZE-1:0] Wgt_2_80;input [WEIGHT_SIZE-1:0] Wgt_2_81;input [WEIGHT_SIZE-1:0] Wgt_2_82;input [WEIGHT_SIZE-1:0] Wgt_2_83;input [WEIGHT_SIZE-1:0] Wgt_2_84;input [WEIGHT_SIZE-1:0] Wgt_2_85;input [WEIGHT_SIZE-1:0] Wgt_2_86;input [WEIGHT_SIZE-1:0] Wgt_2_87;input [WEIGHT_SIZE-1:0] Wgt_2_88;input [WEIGHT_SIZE-1:0] Wgt_2_89;input [WEIGHT_SIZE-1:0] Wgt_2_90;input [WEIGHT_SIZE-1:0] Wgt_2_91;input [WEIGHT_SIZE-1:0] Wgt_2_92;input [WEIGHT_SIZE-1:0] Wgt_2_93;input [WEIGHT_SIZE-1:0] Wgt_2_94;input [WEIGHT_SIZE-1:0] Wgt_2_95;input [WEIGHT_SIZE-1:0] Wgt_2_96;input [WEIGHT_SIZE-1:0] Wgt_2_97;input [WEIGHT_SIZE-1:0] Wgt_2_98;input [WEIGHT_SIZE-1:0] Wgt_2_99;input [WEIGHT_SIZE-1:0] Wgt_2_100;input [WEIGHT_SIZE-1:0] Wgt_2_101;input [WEIGHT_SIZE-1:0] Wgt_2_102;input [WEIGHT_SIZE-1:0] Wgt_2_103;input [WEIGHT_SIZE-1:0] Wgt_2_104;input [WEIGHT_SIZE-1:0] Wgt_2_105;input [WEIGHT_SIZE-1:0] Wgt_2_106;input [WEIGHT_SIZE-1:0] Wgt_2_107;input [WEIGHT_SIZE-1:0] Wgt_2_108;input [WEIGHT_SIZE-1:0] Wgt_2_109;input [WEIGHT_SIZE-1:0] Wgt_2_110;input [WEIGHT_SIZE-1:0] Wgt_2_111;input [WEIGHT_SIZE-1:0] Wgt_2_112;input [WEIGHT_SIZE-1:0] Wgt_2_113;input [WEIGHT_SIZE-1:0] Wgt_2_114;input [WEIGHT_SIZE-1:0] Wgt_2_115;input [WEIGHT_SIZE-1:0] Wgt_2_116;input [WEIGHT_SIZE-1:0] Wgt_2_117;input [WEIGHT_SIZE-1:0] Wgt_2_118;input [WEIGHT_SIZE-1:0] Wgt_2_119;input [WEIGHT_SIZE-1:0] Wgt_2_120;input [WEIGHT_SIZE-1:0] Wgt_2_121;input [WEIGHT_SIZE-1:0] Wgt_2_122;input [WEIGHT_SIZE-1:0] Wgt_2_123;input [WEIGHT_SIZE-1:0] Wgt_2_124;input [WEIGHT_SIZE-1:0] Wgt_2_125;input [WEIGHT_SIZE-1:0] Wgt_2_126;input [WEIGHT_SIZE-1:0] Wgt_2_127;input [WEIGHT_SIZE-1:0] Wgt_2_128;input [WEIGHT_SIZE-1:0] Wgt_2_129;input [WEIGHT_SIZE-1:0] Wgt_2_130;input [WEIGHT_SIZE-1:0] Wgt_2_131;input [WEIGHT_SIZE-1:0] Wgt_2_132;input [WEIGHT_SIZE-1:0] Wgt_2_133;input [WEIGHT_SIZE-1:0] Wgt_2_134;input [WEIGHT_SIZE-1:0] Wgt_2_135;input [WEIGHT_SIZE-1:0] Wgt_2_136;input [WEIGHT_SIZE-1:0] Wgt_2_137;input [WEIGHT_SIZE-1:0] Wgt_2_138;input [WEIGHT_SIZE-1:0] Wgt_2_139;input [WEIGHT_SIZE-1:0] Wgt_2_140;input [WEIGHT_SIZE-1:0] Wgt_2_141;input [WEIGHT_SIZE-1:0] Wgt_2_142;input [WEIGHT_SIZE-1:0] Wgt_2_143;input [WEIGHT_SIZE-1:0] Wgt_2_144;input [WEIGHT_SIZE-1:0] Wgt_2_145;input [WEIGHT_SIZE-1:0] Wgt_2_146;input [WEIGHT_SIZE-1:0] Wgt_2_147;input [WEIGHT_SIZE-1:0] Wgt_2_148;input [WEIGHT_SIZE-1:0] Wgt_2_149;input [WEIGHT_SIZE-1:0] Wgt_2_150;input [WEIGHT_SIZE-1:0] Wgt_2_151;input [WEIGHT_SIZE-1:0] Wgt_2_152;input [WEIGHT_SIZE-1:0] Wgt_2_153;input [WEIGHT_SIZE-1:0] Wgt_2_154;input [WEIGHT_SIZE-1:0] Wgt_2_155;input [WEIGHT_SIZE-1:0] Wgt_2_156;input [WEIGHT_SIZE-1:0] Wgt_2_157;input [WEIGHT_SIZE-1:0] Wgt_2_158;input [WEIGHT_SIZE-1:0] Wgt_2_159;input [WEIGHT_SIZE-1:0] Wgt_2_160;input [WEIGHT_SIZE-1:0] Wgt_2_161;input [WEIGHT_SIZE-1:0] Wgt_2_162;input [WEIGHT_SIZE-1:0] Wgt_2_163;input [WEIGHT_SIZE-1:0] Wgt_2_164;input [WEIGHT_SIZE-1:0] Wgt_2_165;input [WEIGHT_SIZE-1:0] Wgt_2_166;input [WEIGHT_SIZE-1:0] Wgt_2_167;input [WEIGHT_SIZE-1:0] Wgt_2_168;input [WEIGHT_SIZE-1:0] Wgt_2_169;input [WEIGHT_SIZE-1:0] Wgt_2_170;input [WEIGHT_SIZE-1:0] Wgt_2_171;input [WEIGHT_SIZE-1:0] Wgt_2_172;input [WEIGHT_SIZE-1:0] Wgt_2_173;input [WEIGHT_SIZE-1:0] Wgt_2_174;input [WEIGHT_SIZE-1:0] Wgt_2_175;input [WEIGHT_SIZE-1:0] Wgt_2_176;input [WEIGHT_SIZE-1:0] Wgt_2_177;input [WEIGHT_SIZE-1:0] Wgt_2_178;input [WEIGHT_SIZE-1:0] Wgt_2_179;input [WEIGHT_SIZE-1:0] Wgt_2_180;input [WEIGHT_SIZE-1:0] Wgt_2_181;input [WEIGHT_SIZE-1:0] Wgt_2_182;input [WEIGHT_SIZE-1:0] Wgt_2_183;input [WEIGHT_SIZE-1:0] Wgt_2_184;input [WEIGHT_SIZE-1:0] Wgt_2_185;input [WEIGHT_SIZE-1:0] Wgt_2_186;input [WEIGHT_SIZE-1:0] Wgt_2_187;input [WEIGHT_SIZE-1:0] Wgt_2_188;input [WEIGHT_SIZE-1:0] Wgt_2_189;input [WEIGHT_SIZE-1:0] Wgt_2_190;input [WEIGHT_SIZE-1:0] Wgt_2_191;input [WEIGHT_SIZE-1:0] Wgt_2_192;input [WEIGHT_SIZE-1:0] Wgt_2_193;input [WEIGHT_SIZE-1:0] Wgt_2_194;input [WEIGHT_SIZE-1:0] Wgt_2_195;input [WEIGHT_SIZE-1:0] Wgt_2_196;input [WEIGHT_SIZE-1:0] Wgt_2_197;input [WEIGHT_SIZE-1:0] Wgt_2_198;input [WEIGHT_SIZE-1:0] Wgt_2_199;input [WEIGHT_SIZE-1:0] Wgt_2_200;input [WEIGHT_SIZE-1:0] Wgt_2_201;input [WEIGHT_SIZE-1:0] Wgt_2_202;input [WEIGHT_SIZE-1:0] Wgt_2_203;input [WEIGHT_SIZE-1:0] Wgt_2_204;input [WEIGHT_SIZE-1:0] Wgt_2_205;input [WEIGHT_SIZE-1:0] Wgt_2_206;input [WEIGHT_SIZE-1:0] Wgt_2_207;input [WEIGHT_SIZE-1:0] Wgt_2_208;input [WEIGHT_SIZE-1:0] Wgt_2_209;input [WEIGHT_SIZE-1:0] Wgt_2_210;input [WEIGHT_SIZE-1:0] Wgt_2_211;input [WEIGHT_SIZE-1:0] Wgt_2_212;input [WEIGHT_SIZE-1:0] Wgt_2_213;input [WEIGHT_SIZE-1:0] Wgt_2_214;input [WEIGHT_SIZE-1:0] Wgt_2_215;input [WEIGHT_SIZE-1:0] Wgt_2_216;input [WEIGHT_SIZE-1:0] Wgt_2_217;input [WEIGHT_SIZE-1:0] Wgt_2_218;input [WEIGHT_SIZE-1:0] Wgt_2_219;input [WEIGHT_SIZE-1:0] Wgt_2_220;input [WEIGHT_SIZE-1:0] Wgt_2_221;input [WEIGHT_SIZE-1:0] Wgt_2_222;input [WEIGHT_SIZE-1:0] Wgt_2_223;input [WEIGHT_SIZE-1:0] Wgt_2_224;input [WEIGHT_SIZE-1:0] Wgt_2_225;input [WEIGHT_SIZE-1:0] Wgt_2_226;input [WEIGHT_SIZE-1:0] Wgt_2_227;input [WEIGHT_SIZE-1:0] Wgt_2_228;input [WEIGHT_SIZE-1:0] Wgt_2_229;input [WEIGHT_SIZE-1:0] Wgt_2_230;input [WEIGHT_SIZE-1:0] Wgt_2_231;input [WEIGHT_SIZE-1:0] Wgt_2_232;input [WEIGHT_SIZE-1:0] Wgt_2_233;input [WEIGHT_SIZE-1:0] Wgt_2_234;input [WEIGHT_SIZE-1:0] Wgt_2_235;input [WEIGHT_SIZE-1:0] Wgt_2_236;input [WEIGHT_SIZE-1:0] Wgt_2_237;input [WEIGHT_SIZE-1:0] Wgt_2_238;input [WEIGHT_SIZE-1:0] Wgt_2_239;input [WEIGHT_SIZE-1:0] Wgt_2_240;input [WEIGHT_SIZE-1:0] Wgt_2_241;input [WEIGHT_SIZE-1:0] Wgt_2_242;input [WEIGHT_SIZE-1:0] Wgt_2_243;input [WEIGHT_SIZE-1:0] Wgt_2_244;input [WEIGHT_SIZE-1:0] Wgt_2_245;input [WEIGHT_SIZE-1:0] Wgt_2_246;input [WEIGHT_SIZE-1:0] Wgt_2_247;input [WEIGHT_SIZE-1:0] Wgt_2_248;input [WEIGHT_SIZE-1:0] Wgt_2_249;input [WEIGHT_SIZE-1:0] Wgt_2_250;input [WEIGHT_SIZE-1:0] Wgt_2_251;input [WEIGHT_SIZE-1:0] Wgt_2_252;input [WEIGHT_SIZE-1:0] Wgt_2_253;input [WEIGHT_SIZE-1:0] Wgt_2_254;input [WEIGHT_SIZE-1:0] Wgt_2_255;input [WEIGHT_SIZE-1:0] Wgt_2_256;input [WEIGHT_SIZE-1:0] Wgt_2_257;input [WEIGHT_SIZE-1:0] Wgt_2_258;input [WEIGHT_SIZE-1:0] Wgt_2_259;input [WEIGHT_SIZE-1:0] Wgt_2_260;input [WEIGHT_SIZE-1:0] Wgt_2_261;input [WEIGHT_SIZE-1:0] Wgt_2_262;input [WEIGHT_SIZE-1:0] Wgt_2_263;input [WEIGHT_SIZE-1:0] Wgt_2_264;input [WEIGHT_SIZE-1:0] Wgt_2_265;input [WEIGHT_SIZE-1:0] Wgt_2_266;input [WEIGHT_SIZE-1:0] Wgt_2_267;input [WEIGHT_SIZE-1:0] Wgt_2_268;input [WEIGHT_SIZE-1:0] Wgt_2_269;input [WEIGHT_SIZE-1:0] Wgt_2_270;input [WEIGHT_SIZE-1:0] Wgt_2_271;input [WEIGHT_SIZE-1:0] Wgt_2_272;input [WEIGHT_SIZE-1:0] Wgt_2_273;input [WEIGHT_SIZE-1:0] Wgt_2_274;input [WEIGHT_SIZE-1:0] Wgt_2_275;input [WEIGHT_SIZE-1:0] Wgt_2_276;input [WEIGHT_SIZE-1:0] Wgt_2_277;input [WEIGHT_SIZE-1:0] Wgt_2_278;input [WEIGHT_SIZE-1:0] Wgt_2_279;input [WEIGHT_SIZE-1:0] Wgt_2_280;input [WEIGHT_SIZE-1:0] Wgt_2_281;input [WEIGHT_SIZE-1:0] Wgt_2_282;input [WEIGHT_SIZE-1:0] Wgt_2_283;input [WEIGHT_SIZE-1:0] Wgt_2_284;input [WEIGHT_SIZE-1:0] Wgt_2_285;input [WEIGHT_SIZE-1:0] Wgt_2_286;input [WEIGHT_SIZE-1:0] Wgt_2_287;input [WEIGHT_SIZE-1:0] Wgt_2_288;input [WEIGHT_SIZE-1:0] Wgt_2_289;input [WEIGHT_SIZE-1:0] Wgt_2_290;input [WEIGHT_SIZE-1:0] Wgt_2_291;input [WEIGHT_SIZE-1:0] Wgt_2_292;input [WEIGHT_SIZE-1:0] Wgt_2_293;input [WEIGHT_SIZE-1:0] Wgt_2_294;input [WEIGHT_SIZE-1:0] Wgt_2_295;input [WEIGHT_SIZE-1:0] Wgt_2_296;input [WEIGHT_SIZE-1:0] Wgt_2_297;input [WEIGHT_SIZE-1:0] Wgt_2_298;input [WEIGHT_SIZE-1:0] Wgt_2_299;input [WEIGHT_SIZE-1:0] Wgt_2_300;input [WEIGHT_SIZE-1:0] Wgt_2_301;input [WEIGHT_SIZE-1:0] Wgt_2_302;input [WEIGHT_SIZE-1:0] Wgt_2_303;input [WEIGHT_SIZE-1:0] Wgt_2_304;input [WEIGHT_SIZE-1:0] Wgt_2_305;input [WEIGHT_SIZE-1:0] Wgt_2_306;input [WEIGHT_SIZE-1:0] Wgt_2_307;input [WEIGHT_SIZE-1:0] Wgt_2_308;input [WEIGHT_SIZE-1:0] Wgt_2_309;input [WEIGHT_SIZE-1:0] Wgt_2_310;input [WEIGHT_SIZE-1:0] Wgt_2_311;input [WEIGHT_SIZE-1:0] Wgt_2_312;input [WEIGHT_SIZE-1:0] Wgt_2_313;input [WEIGHT_SIZE-1:0] Wgt_2_314;input [WEIGHT_SIZE-1:0] Wgt_2_315;input [WEIGHT_SIZE-1:0] Wgt_2_316;input [WEIGHT_SIZE-1:0] Wgt_2_317;input [WEIGHT_SIZE-1:0] Wgt_2_318;input [WEIGHT_SIZE-1:0] Wgt_2_319;input [WEIGHT_SIZE-1:0] Wgt_2_320;input [WEIGHT_SIZE-1:0] Wgt_2_321;input [WEIGHT_SIZE-1:0] Wgt_2_322;input [WEIGHT_SIZE-1:0] Wgt_2_323;input [WEIGHT_SIZE-1:0] Wgt_2_324;input [WEIGHT_SIZE-1:0] Wgt_2_325;input [WEIGHT_SIZE-1:0] Wgt_2_326;input [WEIGHT_SIZE-1:0] Wgt_2_327;input [WEIGHT_SIZE-1:0] Wgt_2_328;input [WEIGHT_SIZE-1:0] Wgt_2_329;input [WEIGHT_SIZE-1:0] Wgt_2_330;input [WEIGHT_SIZE-1:0] Wgt_2_331;input [WEIGHT_SIZE-1:0] Wgt_2_332;input [WEIGHT_SIZE-1:0] Wgt_2_333;input [WEIGHT_SIZE-1:0] Wgt_2_334;input [WEIGHT_SIZE-1:0] Wgt_2_335;input [WEIGHT_SIZE-1:0] Wgt_2_336;input [WEIGHT_SIZE-1:0] Wgt_2_337;input [WEIGHT_SIZE-1:0] Wgt_2_338;input [WEIGHT_SIZE-1:0] Wgt_2_339;input [WEIGHT_SIZE-1:0] Wgt_2_340;input [WEIGHT_SIZE-1:0] Wgt_2_341;input [WEIGHT_SIZE-1:0] Wgt_2_342;input [WEIGHT_SIZE-1:0] Wgt_2_343;input [WEIGHT_SIZE-1:0] Wgt_2_344;input [WEIGHT_SIZE-1:0] Wgt_2_345;input [WEIGHT_SIZE-1:0] Wgt_2_346;input [WEIGHT_SIZE-1:0] Wgt_2_347;input [WEIGHT_SIZE-1:0] Wgt_2_348;input [WEIGHT_SIZE-1:0] Wgt_2_349;input [WEIGHT_SIZE-1:0] Wgt_2_350;input [WEIGHT_SIZE-1:0] Wgt_2_351;input [WEIGHT_SIZE-1:0] Wgt_2_352;input [WEIGHT_SIZE-1:0] Wgt_2_353;input [WEIGHT_SIZE-1:0] Wgt_2_354;input [WEIGHT_SIZE-1:0] Wgt_2_355;input [WEIGHT_SIZE-1:0] Wgt_2_356;input [WEIGHT_SIZE-1:0] Wgt_2_357;input [WEIGHT_SIZE-1:0] Wgt_2_358;input [WEIGHT_SIZE-1:0] Wgt_2_359;input [WEIGHT_SIZE-1:0] Wgt_2_360;input [WEIGHT_SIZE-1:0] Wgt_2_361;input [WEIGHT_SIZE-1:0] Wgt_2_362;input [WEIGHT_SIZE-1:0] Wgt_2_363;input [WEIGHT_SIZE-1:0] Wgt_2_364;input [WEIGHT_SIZE-1:0] Wgt_2_365;input [WEIGHT_SIZE-1:0] Wgt_2_366;input [WEIGHT_SIZE-1:0] Wgt_2_367;input [WEIGHT_SIZE-1:0] Wgt_2_368;input [WEIGHT_SIZE-1:0] Wgt_2_369;input [WEIGHT_SIZE-1:0] Wgt_2_370;input [WEIGHT_SIZE-1:0] Wgt_2_371;input [WEIGHT_SIZE-1:0] Wgt_2_372;input [WEIGHT_SIZE-1:0] Wgt_2_373;input [WEIGHT_SIZE-1:0] Wgt_2_374;input [WEIGHT_SIZE-1:0] Wgt_2_375;input [WEIGHT_SIZE-1:0] Wgt_2_376;input [WEIGHT_SIZE-1:0] Wgt_2_377;input [WEIGHT_SIZE-1:0] Wgt_2_378;input [WEIGHT_SIZE-1:0] Wgt_2_379;input [WEIGHT_SIZE-1:0] Wgt_2_380;input [WEIGHT_SIZE-1:0] Wgt_2_381;input [WEIGHT_SIZE-1:0] Wgt_2_382;input [WEIGHT_SIZE-1:0] Wgt_2_383;input [WEIGHT_SIZE-1:0] Wgt_2_384;input [WEIGHT_SIZE-1:0] Wgt_2_385;input [WEIGHT_SIZE-1:0] Wgt_2_386;input [WEIGHT_SIZE-1:0] Wgt_2_387;input [WEIGHT_SIZE-1:0] Wgt_2_388;input [WEIGHT_SIZE-1:0] Wgt_2_389;input [WEIGHT_SIZE-1:0] Wgt_2_390;input [WEIGHT_SIZE-1:0] Wgt_2_391;input [WEIGHT_SIZE-1:0] Wgt_2_392;input [WEIGHT_SIZE-1:0] Wgt_2_393;input [WEIGHT_SIZE-1:0] Wgt_2_394;input [WEIGHT_SIZE-1:0] Wgt_2_395;input [WEIGHT_SIZE-1:0] Wgt_2_396;input [WEIGHT_SIZE-1:0] Wgt_2_397;input [WEIGHT_SIZE-1:0] Wgt_2_398;input [WEIGHT_SIZE-1:0] Wgt_2_399;input [WEIGHT_SIZE-1:0] Wgt_2_400;input [WEIGHT_SIZE-1:0] Wgt_2_401;input [WEIGHT_SIZE-1:0] Wgt_2_402;input [WEIGHT_SIZE-1:0] Wgt_2_403;input [WEIGHT_SIZE-1:0] Wgt_2_404;input [WEIGHT_SIZE-1:0] Wgt_2_405;input [WEIGHT_SIZE-1:0] Wgt_2_406;input [WEIGHT_SIZE-1:0] Wgt_2_407;input [WEIGHT_SIZE-1:0] Wgt_2_408;input [WEIGHT_SIZE-1:0] Wgt_2_409;input [WEIGHT_SIZE-1:0] Wgt_2_410;input [WEIGHT_SIZE-1:0] Wgt_2_411;input [WEIGHT_SIZE-1:0] Wgt_2_412;input [WEIGHT_SIZE-1:0] Wgt_2_413;input [WEIGHT_SIZE-1:0] Wgt_2_414;input [WEIGHT_SIZE-1:0] Wgt_2_415;input [WEIGHT_SIZE-1:0] Wgt_2_416;input [WEIGHT_SIZE-1:0] Wgt_2_417;input [WEIGHT_SIZE-1:0] Wgt_2_418;input [WEIGHT_SIZE-1:0] Wgt_2_419;input [WEIGHT_SIZE-1:0] Wgt_2_420;input [WEIGHT_SIZE-1:0] Wgt_2_421;input [WEIGHT_SIZE-1:0] Wgt_2_422;input [WEIGHT_SIZE-1:0] Wgt_2_423;input [WEIGHT_SIZE-1:0] Wgt_2_424;input [WEIGHT_SIZE-1:0] Wgt_2_425;input [WEIGHT_SIZE-1:0] Wgt_2_426;input [WEIGHT_SIZE-1:0] Wgt_2_427;input [WEIGHT_SIZE-1:0] Wgt_2_428;input [WEIGHT_SIZE-1:0] Wgt_2_429;input [WEIGHT_SIZE-1:0] Wgt_2_430;input [WEIGHT_SIZE-1:0] Wgt_2_431;input [WEIGHT_SIZE-1:0] Wgt_2_432;input [WEIGHT_SIZE-1:0] Wgt_2_433;input [WEIGHT_SIZE-1:0] Wgt_2_434;input [WEIGHT_SIZE-1:0] Wgt_2_435;input [WEIGHT_SIZE-1:0] Wgt_2_436;input [WEIGHT_SIZE-1:0] Wgt_2_437;input [WEIGHT_SIZE-1:0] Wgt_2_438;input [WEIGHT_SIZE-1:0] Wgt_2_439;input [WEIGHT_SIZE-1:0] Wgt_2_440;input [WEIGHT_SIZE-1:0] Wgt_2_441;input [WEIGHT_SIZE-1:0] Wgt_2_442;input [WEIGHT_SIZE-1:0] Wgt_2_443;input [WEIGHT_SIZE-1:0] Wgt_2_444;input [WEIGHT_SIZE-1:0] Wgt_2_445;input [WEIGHT_SIZE-1:0] Wgt_2_446;input [WEIGHT_SIZE-1:0] Wgt_2_447;input [WEIGHT_SIZE-1:0] Wgt_2_448;input [WEIGHT_SIZE-1:0] Wgt_2_449;input [WEIGHT_SIZE-1:0] Wgt_2_450;input [WEIGHT_SIZE-1:0] Wgt_2_451;input [WEIGHT_SIZE-1:0] Wgt_2_452;input [WEIGHT_SIZE-1:0] Wgt_2_453;input [WEIGHT_SIZE-1:0] Wgt_2_454;input [WEIGHT_SIZE-1:0] Wgt_2_455;input [WEIGHT_SIZE-1:0] Wgt_2_456;input [WEIGHT_SIZE-1:0] Wgt_2_457;input [WEIGHT_SIZE-1:0] Wgt_2_458;input [WEIGHT_SIZE-1:0] Wgt_2_459;input [WEIGHT_SIZE-1:0] Wgt_2_460;input [WEIGHT_SIZE-1:0] Wgt_2_461;input [WEIGHT_SIZE-1:0] Wgt_2_462;input [WEIGHT_SIZE-1:0] Wgt_2_463;input [WEIGHT_SIZE-1:0] Wgt_2_464;input [WEIGHT_SIZE-1:0] Wgt_2_465;input [WEIGHT_SIZE-1:0] Wgt_2_466;input [WEIGHT_SIZE-1:0] Wgt_2_467;input [WEIGHT_SIZE-1:0] Wgt_2_468;input [WEIGHT_SIZE-1:0] Wgt_2_469;input [WEIGHT_SIZE-1:0] Wgt_2_470;input [WEIGHT_SIZE-1:0] Wgt_2_471;input [WEIGHT_SIZE-1:0] Wgt_2_472;input [WEIGHT_SIZE-1:0] Wgt_2_473;input [WEIGHT_SIZE-1:0] Wgt_2_474;input [WEIGHT_SIZE-1:0] Wgt_2_475;input [WEIGHT_SIZE-1:0] Wgt_2_476;input [WEIGHT_SIZE-1:0] Wgt_2_477;input [WEIGHT_SIZE-1:0] Wgt_2_478;input [WEIGHT_SIZE-1:0] Wgt_2_479;input [WEIGHT_SIZE-1:0] Wgt_2_480;input [WEIGHT_SIZE-1:0] Wgt_2_481;input [WEIGHT_SIZE-1:0] Wgt_2_482;input [WEIGHT_SIZE-1:0] Wgt_2_483;input [WEIGHT_SIZE-1:0] Wgt_2_484;input [WEIGHT_SIZE-1:0] Wgt_2_485;input [WEIGHT_SIZE-1:0] Wgt_2_486;input [WEIGHT_SIZE-1:0] Wgt_2_487;input [WEIGHT_SIZE-1:0] Wgt_2_488;input [WEIGHT_SIZE-1:0] Wgt_2_489;input [WEIGHT_SIZE-1:0] Wgt_2_490;input [WEIGHT_SIZE-1:0] Wgt_2_491;input [WEIGHT_SIZE-1:0] Wgt_2_492;input [WEIGHT_SIZE-1:0] Wgt_2_493;input [WEIGHT_SIZE-1:0] Wgt_2_494;input [WEIGHT_SIZE-1:0] Wgt_2_495;input [WEIGHT_SIZE-1:0] Wgt_2_496;input [WEIGHT_SIZE-1:0] Wgt_2_497;input [WEIGHT_SIZE-1:0] Wgt_2_498;input [WEIGHT_SIZE-1:0] Wgt_2_499;input [WEIGHT_SIZE-1:0] Wgt_2_500;input [WEIGHT_SIZE-1:0] Wgt_2_501;input [WEIGHT_SIZE-1:0] Wgt_2_502;input [WEIGHT_SIZE-1:0] Wgt_2_503;input [WEIGHT_SIZE-1:0] Wgt_2_504;input [WEIGHT_SIZE-1:0] Wgt_2_505;input [WEIGHT_SIZE-1:0] Wgt_2_506;input [WEIGHT_SIZE-1:0] Wgt_2_507;input [WEIGHT_SIZE-1:0] Wgt_2_508;input [WEIGHT_SIZE-1:0] Wgt_2_509;input [WEIGHT_SIZE-1:0] Wgt_2_510;input [WEIGHT_SIZE-1:0] Wgt_2_511;input [WEIGHT_SIZE-1:0] Wgt_2_512;input [WEIGHT_SIZE-1:0] Wgt_2_513;input [WEIGHT_SIZE-1:0] Wgt_2_514;input [WEIGHT_SIZE-1:0] Wgt_2_515;input [WEIGHT_SIZE-1:0] Wgt_2_516;input [WEIGHT_SIZE-1:0] Wgt_2_517;input [WEIGHT_SIZE-1:0] Wgt_2_518;input [WEIGHT_SIZE-1:0] Wgt_2_519;input [WEIGHT_SIZE-1:0] Wgt_2_520;input [WEIGHT_SIZE-1:0] Wgt_2_521;input [WEIGHT_SIZE-1:0] Wgt_2_522;input [WEIGHT_SIZE-1:0] Wgt_2_523;input [WEIGHT_SIZE-1:0] Wgt_2_524;input [WEIGHT_SIZE-1:0] Wgt_2_525;input [WEIGHT_SIZE-1:0] Wgt_2_526;input [WEIGHT_SIZE-1:0] Wgt_2_527;input [WEIGHT_SIZE-1:0] Wgt_2_528;input [WEIGHT_SIZE-1:0] Wgt_2_529;input [WEIGHT_SIZE-1:0] Wgt_2_530;input [WEIGHT_SIZE-1:0] Wgt_2_531;input [WEIGHT_SIZE-1:0] Wgt_2_532;input [WEIGHT_SIZE-1:0] Wgt_2_533;input [WEIGHT_SIZE-1:0] Wgt_2_534;input [WEIGHT_SIZE-1:0] Wgt_2_535;input [WEIGHT_SIZE-1:0] Wgt_2_536;input [WEIGHT_SIZE-1:0] Wgt_2_537;input [WEIGHT_SIZE-1:0] Wgt_2_538;input [WEIGHT_SIZE-1:0] Wgt_2_539;input [WEIGHT_SIZE-1:0] Wgt_2_540;input [WEIGHT_SIZE-1:0] Wgt_2_541;input [WEIGHT_SIZE-1:0] Wgt_2_542;input [WEIGHT_SIZE-1:0] Wgt_2_543;input [WEIGHT_SIZE-1:0] Wgt_2_544;input [WEIGHT_SIZE-1:0] Wgt_2_545;input [WEIGHT_SIZE-1:0] Wgt_2_546;input [WEIGHT_SIZE-1:0] Wgt_2_547;input [WEIGHT_SIZE-1:0] Wgt_2_548;input [WEIGHT_SIZE-1:0] Wgt_2_549;input [WEIGHT_SIZE-1:0] Wgt_2_550;input [WEIGHT_SIZE-1:0] Wgt_2_551;input [WEIGHT_SIZE-1:0] Wgt_2_552;input [WEIGHT_SIZE-1:0] Wgt_2_553;input [WEIGHT_SIZE-1:0] Wgt_2_554;input [WEIGHT_SIZE-1:0] Wgt_2_555;input [WEIGHT_SIZE-1:0] Wgt_2_556;input [WEIGHT_SIZE-1:0] Wgt_2_557;input [WEIGHT_SIZE-1:0] Wgt_2_558;input [WEIGHT_SIZE-1:0] Wgt_2_559;input [WEIGHT_SIZE-1:0] Wgt_2_560;input [WEIGHT_SIZE-1:0] Wgt_2_561;input [WEIGHT_SIZE-1:0] Wgt_2_562;input [WEIGHT_SIZE-1:0] Wgt_2_563;input [WEIGHT_SIZE-1:0] Wgt_2_564;input [WEIGHT_SIZE-1:0] Wgt_2_565;input [WEIGHT_SIZE-1:0] Wgt_2_566;input [WEIGHT_SIZE-1:0] Wgt_2_567;input [WEIGHT_SIZE-1:0] Wgt_2_568;input [WEIGHT_SIZE-1:0] Wgt_2_569;input [WEIGHT_SIZE-1:0] Wgt_2_570;input [WEIGHT_SIZE-1:0] Wgt_2_571;input [WEIGHT_SIZE-1:0] Wgt_2_572;input [WEIGHT_SIZE-1:0] Wgt_2_573;input [WEIGHT_SIZE-1:0] Wgt_2_574;input [WEIGHT_SIZE-1:0] Wgt_2_575;input [WEIGHT_SIZE-1:0] Wgt_2_576;input [WEIGHT_SIZE-1:0] Wgt_2_577;input [WEIGHT_SIZE-1:0] Wgt_2_578;input [WEIGHT_SIZE-1:0] Wgt_2_579;input [WEIGHT_SIZE-1:0] Wgt_2_580;input [WEIGHT_SIZE-1:0] Wgt_2_581;input [WEIGHT_SIZE-1:0] Wgt_2_582;input [WEIGHT_SIZE-1:0] Wgt_2_583;input [WEIGHT_SIZE-1:0] Wgt_2_584;input [WEIGHT_SIZE-1:0] Wgt_2_585;input [WEIGHT_SIZE-1:0] Wgt_2_586;input [WEIGHT_SIZE-1:0] Wgt_2_587;input [WEIGHT_SIZE-1:0] Wgt_2_588;input [WEIGHT_SIZE-1:0] Wgt_2_589;input [WEIGHT_SIZE-1:0] Wgt_2_590;input [WEIGHT_SIZE-1:0] Wgt_2_591;input [WEIGHT_SIZE-1:0] Wgt_2_592;input [WEIGHT_SIZE-1:0] Wgt_2_593;input [WEIGHT_SIZE-1:0] Wgt_2_594;input [WEIGHT_SIZE-1:0] Wgt_2_595;input [WEIGHT_SIZE-1:0] Wgt_2_596;input [WEIGHT_SIZE-1:0] Wgt_2_597;input [WEIGHT_SIZE-1:0] Wgt_2_598;input [WEIGHT_SIZE-1:0] Wgt_2_599;input [WEIGHT_SIZE-1:0] Wgt_2_600;input [WEIGHT_SIZE-1:0] Wgt_2_601;input [WEIGHT_SIZE-1:0] Wgt_2_602;input [WEIGHT_SIZE-1:0] Wgt_2_603;input [WEIGHT_SIZE-1:0] Wgt_2_604;input [WEIGHT_SIZE-1:0] Wgt_2_605;input [WEIGHT_SIZE-1:0] Wgt_2_606;input [WEIGHT_SIZE-1:0] Wgt_2_607;input [WEIGHT_SIZE-1:0] Wgt_2_608;input [WEIGHT_SIZE-1:0] Wgt_2_609;input [WEIGHT_SIZE-1:0] Wgt_2_610;input [WEIGHT_SIZE-1:0] Wgt_2_611;input [WEIGHT_SIZE-1:0] Wgt_2_612;input [WEIGHT_SIZE-1:0] Wgt_2_613;input [WEIGHT_SIZE-1:0] Wgt_2_614;input [WEIGHT_SIZE-1:0] Wgt_2_615;input [WEIGHT_SIZE-1:0] Wgt_2_616;input [WEIGHT_SIZE-1:0] Wgt_2_617;input [WEIGHT_SIZE-1:0] Wgt_2_618;input [WEIGHT_SIZE-1:0] Wgt_2_619;input [WEIGHT_SIZE-1:0] Wgt_2_620;input [WEIGHT_SIZE-1:0] Wgt_2_621;input [WEIGHT_SIZE-1:0] Wgt_2_622;input [WEIGHT_SIZE-1:0] Wgt_2_623;input [WEIGHT_SIZE-1:0] Wgt_2_624;input [WEIGHT_SIZE-1:0] Wgt_2_625;input [WEIGHT_SIZE-1:0] Wgt_2_626;input [WEIGHT_SIZE-1:0] Wgt_2_627;input [WEIGHT_SIZE-1:0] Wgt_2_628;input [WEIGHT_SIZE-1:0] Wgt_2_629;input [WEIGHT_SIZE-1:0] Wgt_2_630;input [WEIGHT_SIZE-1:0] Wgt_2_631;input [WEIGHT_SIZE-1:0] Wgt_2_632;input [WEIGHT_SIZE-1:0] Wgt_2_633;input [WEIGHT_SIZE-1:0] Wgt_2_634;input [WEIGHT_SIZE-1:0] Wgt_2_635;input [WEIGHT_SIZE-1:0] Wgt_2_636;input [WEIGHT_SIZE-1:0] Wgt_2_637;input [WEIGHT_SIZE-1:0] Wgt_2_638;input [WEIGHT_SIZE-1:0] Wgt_2_639;input [WEIGHT_SIZE-1:0] Wgt_2_640;input [WEIGHT_SIZE-1:0] Wgt_2_641;input [WEIGHT_SIZE-1:0] Wgt_2_642;input [WEIGHT_SIZE-1:0] Wgt_2_643;input [WEIGHT_SIZE-1:0] Wgt_2_644;input [WEIGHT_SIZE-1:0] Wgt_2_645;input [WEIGHT_SIZE-1:0] Wgt_2_646;input [WEIGHT_SIZE-1:0] Wgt_2_647;input [WEIGHT_SIZE-1:0] Wgt_2_648;input [WEIGHT_SIZE-1:0] Wgt_2_649;input [WEIGHT_SIZE-1:0] Wgt_2_650;input [WEIGHT_SIZE-1:0] Wgt_2_651;input [WEIGHT_SIZE-1:0] Wgt_2_652;input [WEIGHT_SIZE-1:0] Wgt_2_653;input [WEIGHT_SIZE-1:0] Wgt_2_654;input [WEIGHT_SIZE-1:0] Wgt_2_655;input [WEIGHT_SIZE-1:0] Wgt_2_656;input [WEIGHT_SIZE-1:0] Wgt_2_657;input [WEIGHT_SIZE-1:0] Wgt_2_658;input [WEIGHT_SIZE-1:0] Wgt_2_659;input [WEIGHT_SIZE-1:0] Wgt_2_660;input [WEIGHT_SIZE-1:0] Wgt_2_661;input [WEIGHT_SIZE-1:0] Wgt_2_662;input [WEIGHT_SIZE-1:0] Wgt_2_663;input [WEIGHT_SIZE-1:0] Wgt_2_664;input [WEIGHT_SIZE-1:0] Wgt_2_665;input [WEIGHT_SIZE-1:0] Wgt_2_666;input [WEIGHT_SIZE-1:0] Wgt_2_667;input [WEIGHT_SIZE-1:0] Wgt_2_668;input [WEIGHT_SIZE-1:0] Wgt_2_669;input [WEIGHT_SIZE-1:0] Wgt_2_670;input [WEIGHT_SIZE-1:0] Wgt_2_671;input [WEIGHT_SIZE-1:0] Wgt_2_672;input [WEIGHT_SIZE-1:0] Wgt_2_673;input [WEIGHT_SIZE-1:0] Wgt_2_674;input [WEIGHT_SIZE-1:0] Wgt_2_675;input [WEIGHT_SIZE-1:0] Wgt_2_676;input [WEIGHT_SIZE-1:0] Wgt_2_677;input [WEIGHT_SIZE-1:0] Wgt_2_678;input [WEIGHT_SIZE-1:0] Wgt_2_679;input [WEIGHT_SIZE-1:0] Wgt_2_680;input [WEIGHT_SIZE-1:0] Wgt_2_681;input [WEIGHT_SIZE-1:0] Wgt_2_682;input [WEIGHT_SIZE-1:0] Wgt_2_683;input [WEIGHT_SIZE-1:0] Wgt_2_684;input [WEIGHT_SIZE-1:0] Wgt_2_685;input [WEIGHT_SIZE-1:0] Wgt_2_686;input [WEIGHT_SIZE-1:0] Wgt_2_687;input [WEIGHT_SIZE-1:0] Wgt_2_688;input [WEIGHT_SIZE-1:0] Wgt_2_689;input [WEIGHT_SIZE-1:0] Wgt_2_690;input [WEIGHT_SIZE-1:0] Wgt_2_691;input [WEIGHT_SIZE-1:0] Wgt_2_692;input [WEIGHT_SIZE-1:0] Wgt_2_693;input [WEIGHT_SIZE-1:0] Wgt_2_694;input [WEIGHT_SIZE-1:0] Wgt_2_695;input [WEIGHT_SIZE-1:0] Wgt_2_696;input [WEIGHT_SIZE-1:0] Wgt_2_697;input [WEIGHT_SIZE-1:0] Wgt_2_698;input [WEIGHT_SIZE-1:0] Wgt_2_699;input [WEIGHT_SIZE-1:0] Wgt_2_700;input [WEIGHT_SIZE-1:0] Wgt_2_701;input [WEIGHT_SIZE-1:0] Wgt_2_702;input [WEIGHT_SIZE-1:0] Wgt_2_703;input [WEIGHT_SIZE-1:0] Wgt_2_704;input [WEIGHT_SIZE-1:0] Wgt_2_705;input [WEIGHT_SIZE-1:0] Wgt_2_706;input [WEIGHT_SIZE-1:0] Wgt_2_707;input [WEIGHT_SIZE-1:0] Wgt_2_708;input [WEIGHT_SIZE-1:0] Wgt_2_709;input [WEIGHT_SIZE-1:0] Wgt_2_710;input [WEIGHT_SIZE-1:0] Wgt_2_711;input [WEIGHT_SIZE-1:0] Wgt_2_712;input [WEIGHT_SIZE-1:0] Wgt_2_713;input [WEIGHT_SIZE-1:0] Wgt_2_714;input [WEIGHT_SIZE-1:0] Wgt_2_715;input [WEIGHT_SIZE-1:0] Wgt_2_716;input [WEIGHT_SIZE-1:0] Wgt_2_717;input [WEIGHT_SIZE-1:0] Wgt_2_718;input [WEIGHT_SIZE-1:0] Wgt_2_719;input [WEIGHT_SIZE-1:0] Wgt_2_720;input [WEIGHT_SIZE-1:0] Wgt_2_721;input [WEIGHT_SIZE-1:0] Wgt_2_722;input [WEIGHT_SIZE-1:0] Wgt_2_723;input [WEIGHT_SIZE-1:0] Wgt_2_724;input [WEIGHT_SIZE-1:0] Wgt_2_725;input [WEIGHT_SIZE-1:0] Wgt_2_726;input [WEIGHT_SIZE-1:0] Wgt_2_727;input [WEIGHT_SIZE-1:0] Wgt_2_728;input [WEIGHT_SIZE-1:0] Wgt_2_729;input [WEIGHT_SIZE-1:0] Wgt_2_730;input [WEIGHT_SIZE-1:0] Wgt_2_731;input [WEIGHT_SIZE-1:0] Wgt_2_732;input [WEIGHT_SIZE-1:0] Wgt_2_733;input [WEIGHT_SIZE-1:0] Wgt_2_734;input [WEIGHT_SIZE-1:0] Wgt_2_735;input [WEIGHT_SIZE-1:0] Wgt_2_736;input [WEIGHT_SIZE-1:0] Wgt_2_737;input [WEIGHT_SIZE-1:0] Wgt_2_738;input [WEIGHT_SIZE-1:0] Wgt_2_739;input [WEIGHT_SIZE-1:0] Wgt_2_740;input [WEIGHT_SIZE-1:0] Wgt_2_741;input [WEIGHT_SIZE-1:0] Wgt_2_742;input [WEIGHT_SIZE-1:0] Wgt_2_743;input [WEIGHT_SIZE-1:0] Wgt_2_744;input [WEIGHT_SIZE-1:0] Wgt_2_745;input [WEIGHT_SIZE-1:0] Wgt_2_746;input [WEIGHT_SIZE-1:0] Wgt_2_747;input [WEIGHT_SIZE-1:0] Wgt_2_748;input [WEIGHT_SIZE-1:0] Wgt_2_749;input [WEIGHT_SIZE-1:0] Wgt_2_750;input [WEIGHT_SIZE-1:0] Wgt_2_751;input [WEIGHT_SIZE-1:0] Wgt_2_752;input [WEIGHT_SIZE-1:0] Wgt_2_753;input [WEIGHT_SIZE-1:0] Wgt_2_754;input [WEIGHT_SIZE-1:0] Wgt_2_755;input [WEIGHT_SIZE-1:0] Wgt_2_756;input [WEIGHT_SIZE-1:0] Wgt_2_757;input [WEIGHT_SIZE-1:0] Wgt_2_758;input [WEIGHT_SIZE-1:0] Wgt_2_759;input [WEIGHT_SIZE-1:0] Wgt_2_760;input [WEIGHT_SIZE-1:0] Wgt_2_761;input [WEIGHT_SIZE-1:0] Wgt_2_762;input [WEIGHT_SIZE-1:0] Wgt_2_763;input [WEIGHT_SIZE-1:0] Wgt_2_764;input [WEIGHT_SIZE-1:0] Wgt_2_765;input [WEIGHT_SIZE-1:0] Wgt_2_766;input [WEIGHT_SIZE-1:0] Wgt_2_767;input [WEIGHT_SIZE-1:0] Wgt_2_768;input [WEIGHT_SIZE-1:0] Wgt_2_769;input [WEIGHT_SIZE-1:0] Wgt_2_770;input [WEIGHT_SIZE-1:0] Wgt_2_771;input [WEIGHT_SIZE-1:0] Wgt_2_772;input [WEIGHT_SIZE-1:0] Wgt_2_773;input [WEIGHT_SIZE-1:0] Wgt_2_774;input [WEIGHT_SIZE-1:0] Wgt_2_775;input [WEIGHT_SIZE-1:0] Wgt_2_776;input [WEIGHT_SIZE-1:0] Wgt_2_777;input [WEIGHT_SIZE-1:0] Wgt_2_778;input [WEIGHT_SIZE-1:0] Wgt_2_779;input [WEIGHT_SIZE-1:0] Wgt_2_780;input [WEIGHT_SIZE-1:0] Wgt_2_781;input [WEIGHT_SIZE-1:0] Wgt_2_782;input [WEIGHT_SIZE-1:0] Wgt_2_783;input [WEIGHT_SIZE-1:0] Wgt_2_784;input [WEIGHT_SIZE-1:0] Wgt_3_0;input [WEIGHT_SIZE-1:0] Wgt_3_1;input [WEIGHT_SIZE-1:0] Wgt_3_2;input [WEIGHT_SIZE-1:0] Wgt_3_3;input [WEIGHT_SIZE-1:0] Wgt_3_4;input [WEIGHT_SIZE-1:0] Wgt_3_5;input [WEIGHT_SIZE-1:0] Wgt_3_6;input [WEIGHT_SIZE-1:0] Wgt_3_7;input [WEIGHT_SIZE-1:0] Wgt_3_8;input [WEIGHT_SIZE-1:0] Wgt_3_9;input [WEIGHT_SIZE-1:0] Wgt_3_10;input [WEIGHT_SIZE-1:0] Wgt_3_11;input [WEIGHT_SIZE-1:0] Wgt_3_12;input [WEIGHT_SIZE-1:0] Wgt_3_13;input [WEIGHT_SIZE-1:0] Wgt_3_14;input [WEIGHT_SIZE-1:0] Wgt_3_15;input [WEIGHT_SIZE-1:0] Wgt_3_16;input [WEIGHT_SIZE-1:0] Wgt_3_17;input [WEIGHT_SIZE-1:0] Wgt_3_18;input [WEIGHT_SIZE-1:0] Wgt_3_19;input [WEIGHT_SIZE-1:0] Wgt_3_20;input [WEIGHT_SIZE-1:0] Wgt_3_21;input [WEIGHT_SIZE-1:0] Wgt_3_22;input [WEIGHT_SIZE-1:0] Wgt_3_23;input [WEIGHT_SIZE-1:0] Wgt_3_24;input [WEIGHT_SIZE-1:0] Wgt_3_25;input [WEIGHT_SIZE-1:0] Wgt_3_26;input [WEIGHT_SIZE-1:0] Wgt_3_27;input [WEIGHT_SIZE-1:0] Wgt_3_28;input [WEIGHT_SIZE-1:0] Wgt_3_29;input [WEIGHT_SIZE-1:0] Wgt_3_30;input [WEIGHT_SIZE-1:0] Wgt_3_31;input [WEIGHT_SIZE-1:0] Wgt_3_32;input [WEIGHT_SIZE-1:0] Wgt_3_33;input [WEIGHT_SIZE-1:0] Wgt_3_34;input [WEIGHT_SIZE-1:0] Wgt_3_35;input [WEIGHT_SIZE-1:0] Wgt_3_36;input [WEIGHT_SIZE-1:0] Wgt_3_37;input [WEIGHT_SIZE-1:0] Wgt_3_38;input [WEIGHT_SIZE-1:0] Wgt_3_39;input [WEIGHT_SIZE-1:0] Wgt_3_40;input [WEIGHT_SIZE-1:0] Wgt_3_41;input [WEIGHT_SIZE-1:0] Wgt_3_42;input [WEIGHT_SIZE-1:0] Wgt_3_43;input [WEIGHT_SIZE-1:0] Wgt_3_44;input [WEIGHT_SIZE-1:0] Wgt_3_45;input [WEIGHT_SIZE-1:0] Wgt_3_46;input [WEIGHT_SIZE-1:0] Wgt_3_47;input [WEIGHT_SIZE-1:0] Wgt_3_48;input [WEIGHT_SIZE-1:0] Wgt_3_49;input [WEIGHT_SIZE-1:0] Wgt_3_50;input [WEIGHT_SIZE-1:0] Wgt_3_51;input [WEIGHT_SIZE-1:0] Wgt_3_52;input [WEIGHT_SIZE-1:0] Wgt_3_53;input [WEIGHT_SIZE-1:0] Wgt_3_54;input [WEIGHT_SIZE-1:0] Wgt_3_55;input [WEIGHT_SIZE-1:0] Wgt_3_56;input [WEIGHT_SIZE-1:0] Wgt_3_57;input [WEIGHT_SIZE-1:0] Wgt_3_58;input [WEIGHT_SIZE-1:0] Wgt_3_59;input [WEIGHT_SIZE-1:0] Wgt_3_60;input [WEIGHT_SIZE-1:0] Wgt_3_61;input [WEIGHT_SIZE-1:0] Wgt_3_62;input [WEIGHT_SIZE-1:0] Wgt_3_63;input [WEIGHT_SIZE-1:0] Wgt_3_64;input [WEIGHT_SIZE-1:0] Wgt_3_65;input [WEIGHT_SIZE-1:0] Wgt_3_66;input [WEIGHT_SIZE-1:0] Wgt_3_67;input [WEIGHT_SIZE-1:0] Wgt_3_68;input [WEIGHT_SIZE-1:0] Wgt_3_69;input [WEIGHT_SIZE-1:0] Wgt_3_70;input [WEIGHT_SIZE-1:0] Wgt_3_71;input [WEIGHT_SIZE-1:0] Wgt_3_72;input [WEIGHT_SIZE-1:0] Wgt_3_73;input [WEIGHT_SIZE-1:0] Wgt_3_74;input [WEIGHT_SIZE-1:0] Wgt_3_75;input [WEIGHT_SIZE-1:0] Wgt_3_76;input [WEIGHT_SIZE-1:0] Wgt_3_77;input [WEIGHT_SIZE-1:0] Wgt_3_78;input [WEIGHT_SIZE-1:0] Wgt_3_79;input [WEIGHT_SIZE-1:0] Wgt_3_80;input [WEIGHT_SIZE-1:0] Wgt_3_81;input [WEIGHT_SIZE-1:0] Wgt_3_82;input [WEIGHT_SIZE-1:0] Wgt_3_83;input [WEIGHT_SIZE-1:0] Wgt_3_84;input [WEIGHT_SIZE-1:0] Wgt_3_85;input [WEIGHT_SIZE-1:0] Wgt_3_86;input [WEIGHT_SIZE-1:0] Wgt_3_87;input [WEIGHT_SIZE-1:0] Wgt_3_88;input [WEIGHT_SIZE-1:0] Wgt_3_89;input [WEIGHT_SIZE-1:0] Wgt_3_90;input [WEIGHT_SIZE-1:0] Wgt_3_91;input [WEIGHT_SIZE-1:0] Wgt_3_92;input [WEIGHT_SIZE-1:0] Wgt_3_93;input [WEIGHT_SIZE-1:0] Wgt_3_94;input [WEIGHT_SIZE-1:0] Wgt_3_95;input [WEIGHT_SIZE-1:0] Wgt_3_96;input [WEIGHT_SIZE-1:0] Wgt_3_97;input [WEIGHT_SIZE-1:0] Wgt_3_98;input [WEIGHT_SIZE-1:0] Wgt_3_99;input [WEIGHT_SIZE-1:0] Wgt_3_100;input [WEIGHT_SIZE-1:0] Wgt_3_101;input [WEIGHT_SIZE-1:0] Wgt_3_102;input [WEIGHT_SIZE-1:0] Wgt_3_103;input [WEIGHT_SIZE-1:0] Wgt_3_104;input [WEIGHT_SIZE-1:0] Wgt_3_105;input [WEIGHT_SIZE-1:0] Wgt_3_106;input [WEIGHT_SIZE-1:0] Wgt_3_107;input [WEIGHT_SIZE-1:0] Wgt_3_108;input [WEIGHT_SIZE-1:0] Wgt_3_109;input [WEIGHT_SIZE-1:0] Wgt_3_110;input [WEIGHT_SIZE-1:0] Wgt_3_111;input [WEIGHT_SIZE-1:0] Wgt_3_112;input [WEIGHT_SIZE-1:0] Wgt_3_113;input [WEIGHT_SIZE-1:0] Wgt_3_114;input [WEIGHT_SIZE-1:0] Wgt_3_115;input [WEIGHT_SIZE-1:0] Wgt_3_116;input [WEIGHT_SIZE-1:0] Wgt_3_117;input [WEIGHT_SIZE-1:0] Wgt_3_118;input [WEIGHT_SIZE-1:0] Wgt_3_119;input [WEIGHT_SIZE-1:0] Wgt_3_120;input [WEIGHT_SIZE-1:0] Wgt_3_121;input [WEIGHT_SIZE-1:0] Wgt_3_122;input [WEIGHT_SIZE-1:0] Wgt_3_123;input [WEIGHT_SIZE-1:0] Wgt_3_124;input [WEIGHT_SIZE-1:0] Wgt_3_125;input [WEIGHT_SIZE-1:0] Wgt_3_126;input [WEIGHT_SIZE-1:0] Wgt_3_127;input [WEIGHT_SIZE-1:0] Wgt_3_128;input [WEIGHT_SIZE-1:0] Wgt_3_129;input [WEIGHT_SIZE-1:0] Wgt_3_130;input [WEIGHT_SIZE-1:0] Wgt_3_131;input [WEIGHT_SIZE-1:0] Wgt_3_132;input [WEIGHT_SIZE-1:0] Wgt_3_133;input [WEIGHT_SIZE-1:0] Wgt_3_134;input [WEIGHT_SIZE-1:0] Wgt_3_135;input [WEIGHT_SIZE-1:0] Wgt_3_136;input [WEIGHT_SIZE-1:0] Wgt_3_137;input [WEIGHT_SIZE-1:0] Wgt_3_138;input [WEIGHT_SIZE-1:0] Wgt_3_139;input [WEIGHT_SIZE-1:0] Wgt_3_140;input [WEIGHT_SIZE-1:0] Wgt_3_141;input [WEIGHT_SIZE-1:0] Wgt_3_142;input [WEIGHT_SIZE-1:0] Wgt_3_143;input [WEIGHT_SIZE-1:0] Wgt_3_144;input [WEIGHT_SIZE-1:0] Wgt_3_145;input [WEIGHT_SIZE-1:0] Wgt_3_146;input [WEIGHT_SIZE-1:0] Wgt_3_147;input [WEIGHT_SIZE-1:0] Wgt_3_148;input [WEIGHT_SIZE-1:0] Wgt_3_149;input [WEIGHT_SIZE-1:0] Wgt_3_150;input [WEIGHT_SIZE-1:0] Wgt_3_151;input [WEIGHT_SIZE-1:0] Wgt_3_152;input [WEIGHT_SIZE-1:0] Wgt_3_153;input [WEIGHT_SIZE-1:0] Wgt_3_154;input [WEIGHT_SIZE-1:0] Wgt_3_155;input [WEIGHT_SIZE-1:0] Wgt_3_156;input [WEIGHT_SIZE-1:0] Wgt_3_157;input [WEIGHT_SIZE-1:0] Wgt_3_158;input [WEIGHT_SIZE-1:0] Wgt_3_159;input [WEIGHT_SIZE-1:0] Wgt_3_160;input [WEIGHT_SIZE-1:0] Wgt_3_161;input [WEIGHT_SIZE-1:0] Wgt_3_162;input [WEIGHT_SIZE-1:0] Wgt_3_163;input [WEIGHT_SIZE-1:0] Wgt_3_164;input [WEIGHT_SIZE-1:0] Wgt_3_165;input [WEIGHT_SIZE-1:0] Wgt_3_166;input [WEIGHT_SIZE-1:0] Wgt_3_167;input [WEIGHT_SIZE-1:0] Wgt_3_168;input [WEIGHT_SIZE-1:0] Wgt_3_169;input [WEIGHT_SIZE-1:0] Wgt_3_170;input [WEIGHT_SIZE-1:0] Wgt_3_171;input [WEIGHT_SIZE-1:0] Wgt_3_172;input [WEIGHT_SIZE-1:0] Wgt_3_173;input [WEIGHT_SIZE-1:0] Wgt_3_174;input [WEIGHT_SIZE-1:0] Wgt_3_175;input [WEIGHT_SIZE-1:0] Wgt_3_176;input [WEIGHT_SIZE-1:0] Wgt_3_177;input [WEIGHT_SIZE-1:0] Wgt_3_178;input [WEIGHT_SIZE-1:0] Wgt_3_179;input [WEIGHT_SIZE-1:0] Wgt_3_180;input [WEIGHT_SIZE-1:0] Wgt_3_181;input [WEIGHT_SIZE-1:0] Wgt_3_182;input [WEIGHT_SIZE-1:0] Wgt_3_183;input [WEIGHT_SIZE-1:0] Wgt_3_184;input [WEIGHT_SIZE-1:0] Wgt_3_185;input [WEIGHT_SIZE-1:0] Wgt_3_186;input [WEIGHT_SIZE-1:0] Wgt_3_187;input [WEIGHT_SIZE-1:0] Wgt_3_188;input [WEIGHT_SIZE-1:0] Wgt_3_189;input [WEIGHT_SIZE-1:0] Wgt_3_190;input [WEIGHT_SIZE-1:0] Wgt_3_191;input [WEIGHT_SIZE-1:0] Wgt_3_192;input [WEIGHT_SIZE-1:0] Wgt_3_193;input [WEIGHT_SIZE-1:0] Wgt_3_194;input [WEIGHT_SIZE-1:0] Wgt_3_195;input [WEIGHT_SIZE-1:0] Wgt_3_196;input [WEIGHT_SIZE-1:0] Wgt_3_197;input [WEIGHT_SIZE-1:0] Wgt_3_198;input [WEIGHT_SIZE-1:0] Wgt_3_199;input [WEIGHT_SIZE-1:0] Wgt_3_200;input [WEIGHT_SIZE-1:0] Wgt_3_201;input [WEIGHT_SIZE-1:0] Wgt_3_202;input [WEIGHT_SIZE-1:0] Wgt_3_203;input [WEIGHT_SIZE-1:0] Wgt_3_204;input [WEIGHT_SIZE-1:0] Wgt_3_205;input [WEIGHT_SIZE-1:0] Wgt_3_206;input [WEIGHT_SIZE-1:0] Wgt_3_207;input [WEIGHT_SIZE-1:0] Wgt_3_208;input [WEIGHT_SIZE-1:0] Wgt_3_209;input [WEIGHT_SIZE-1:0] Wgt_3_210;input [WEIGHT_SIZE-1:0] Wgt_3_211;input [WEIGHT_SIZE-1:0] Wgt_3_212;input [WEIGHT_SIZE-1:0] Wgt_3_213;input [WEIGHT_SIZE-1:0] Wgt_3_214;input [WEIGHT_SIZE-1:0] Wgt_3_215;input [WEIGHT_SIZE-1:0] Wgt_3_216;input [WEIGHT_SIZE-1:0] Wgt_3_217;input [WEIGHT_SIZE-1:0] Wgt_3_218;input [WEIGHT_SIZE-1:0] Wgt_3_219;input [WEIGHT_SIZE-1:0] Wgt_3_220;input [WEIGHT_SIZE-1:0] Wgt_3_221;input [WEIGHT_SIZE-1:0] Wgt_3_222;input [WEIGHT_SIZE-1:0] Wgt_3_223;input [WEIGHT_SIZE-1:0] Wgt_3_224;input [WEIGHT_SIZE-1:0] Wgt_3_225;input [WEIGHT_SIZE-1:0] Wgt_3_226;input [WEIGHT_SIZE-1:0] Wgt_3_227;input [WEIGHT_SIZE-1:0] Wgt_3_228;input [WEIGHT_SIZE-1:0] Wgt_3_229;input [WEIGHT_SIZE-1:0] Wgt_3_230;input [WEIGHT_SIZE-1:0] Wgt_3_231;input [WEIGHT_SIZE-1:0] Wgt_3_232;input [WEIGHT_SIZE-1:0] Wgt_3_233;input [WEIGHT_SIZE-1:0] Wgt_3_234;input [WEIGHT_SIZE-1:0] Wgt_3_235;input [WEIGHT_SIZE-1:0] Wgt_3_236;input [WEIGHT_SIZE-1:0] Wgt_3_237;input [WEIGHT_SIZE-1:0] Wgt_3_238;input [WEIGHT_SIZE-1:0] Wgt_3_239;input [WEIGHT_SIZE-1:0] Wgt_3_240;input [WEIGHT_SIZE-1:0] Wgt_3_241;input [WEIGHT_SIZE-1:0] Wgt_3_242;input [WEIGHT_SIZE-1:0] Wgt_3_243;input [WEIGHT_SIZE-1:0] Wgt_3_244;input [WEIGHT_SIZE-1:0] Wgt_3_245;input [WEIGHT_SIZE-1:0] Wgt_3_246;input [WEIGHT_SIZE-1:0] Wgt_3_247;input [WEIGHT_SIZE-1:0] Wgt_3_248;input [WEIGHT_SIZE-1:0] Wgt_3_249;input [WEIGHT_SIZE-1:0] Wgt_3_250;input [WEIGHT_SIZE-1:0] Wgt_3_251;input [WEIGHT_SIZE-1:0] Wgt_3_252;input [WEIGHT_SIZE-1:0] Wgt_3_253;input [WEIGHT_SIZE-1:0] Wgt_3_254;input [WEIGHT_SIZE-1:0] Wgt_3_255;input [WEIGHT_SIZE-1:0] Wgt_3_256;input [WEIGHT_SIZE-1:0] Wgt_3_257;input [WEIGHT_SIZE-1:0] Wgt_3_258;input [WEIGHT_SIZE-1:0] Wgt_3_259;input [WEIGHT_SIZE-1:0] Wgt_3_260;input [WEIGHT_SIZE-1:0] Wgt_3_261;input [WEIGHT_SIZE-1:0] Wgt_3_262;input [WEIGHT_SIZE-1:0] Wgt_3_263;input [WEIGHT_SIZE-1:0] Wgt_3_264;input [WEIGHT_SIZE-1:0] Wgt_3_265;input [WEIGHT_SIZE-1:0] Wgt_3_266;input [WEIGHT_SIZE-1:0] Wgt_3_267;input [WEIGHT_SIZE-1:0] Wgt_3_268;input [WEIGHT_SIZE-1:0] Wgt_3_269;input [WEIGHT_SIZE-1:0] Wgt_3_270;input [WEIGHT_SIZE-1:0] Wgt_3_271;input [WEIGHT_SIZE-1:0] Wgt_3_272;input [WEIGHT_SIZE-1:0] Wgt_3_273;input [WEIGHT_SIZE-1:0] Wgt_3_274;input [WEIGHT_SIZE-1:0] Wgt_3_275;input [WEIGHT_SIZE-1:0] Wgt_3_276;input [WEIGHT_SIZE-1:0] Wgt_3_277;input [WEIGHT_SIZE-1:0] Wgt_3_278;input [WEIGHT_SIZE-1:0] Wgt_3_279;input [WEIGHT_SIZE-1:0] Wgt_3_280;input [WEIGHT_SIZE-1:0] Wgt_3_281;input [WEIGHT_SIZE-1:0] Wgt_3_282;input [WEIGHT_SIZE-1:0] Wgt_3_283;input [WEIGHT_SIZE-1:0] Wgt_3_284;input [WEIGHT_SIZE-1:0] Wgt_3_285;input [WEIGHT_SIZE-1:0] Wgt_3_286;input [WEIGHT_SIZE-1:0] Wgt_3_287;input [WEIGHT_SIZE-1:0] Wgt_3_288;input [WEIGHT_SIZE-1:0] Wgt_3_289;input [WEIGHT_SIZE-1:0] Wgt_3_290;input [WEIGHT_SIZE-1:0] Wgt_3_291;input [WEIGHT_SIZE-1:0] Wgt_3_292;input [WEIGHT_SIZE-1:0] Wgt_3_293;input [WEIGHT_SIZE-1:0] Wgt_3_294;input [WEIGHT_SIZE-1:0] Wgt_3_295;input [WEIGHT_SIZE-1:0] Wgt_3_296;input [WEIGHT_SIZE-1:0] Wgt_3_297;input [WEIGHT_SIZE-1:0] Wgt_3_298;input [WEIGHT_SIZE-1:0] Wgt_3_299;input [WEIGHT_SIZE-1:0] Wgt_3_300;input [WEIGHT_SIZE-1:0] Wgt_3_301;input [WEIGHT_SIZE-1:0] Wgt_3_302;input [WEIGHT_SIZE-1:0] Wgt_3_303;input [WEIGHT_SIZE-1:0] Wgt_3_304;input [WEIGHT_SIZE-1:0] Wgt_3_305;input [WEIGHT_SIZE-1:0] Wgt_3_306;input [WEIGHT_SIZE-1:0] Wgt_3_307;input [WEIGHT_SIZE-1:0] Wgt_3_308;input [WEIGHT_SIZE-1:0] Wgt_3_309;input [WEIGHT_SIZE-1:0] Wgt_3_310;input [WEIGHT_SIZE-1:0] Wgt_3_311;input [WEIGHT_SIZE-1:0] Wgt_3_312;input [WEIGHT_SIZE-1:0] Wgt_3_313;input [WEIGHT_SIZE-1:0] Wgt_3_314;input [WEIGHT_SIZE-1:0] Wgt_3_315;input [WEIGHT_SIZE-1:0] Wgt_3_316;input [WEIGHT_SIZE-1:0] Wgt_3_317;input [WEIGHT_SIZE-1:0] Wgt_3_318;input [WEIGHT_SIZE-1:0] Wgt_3_319;input [WEIGHT_SIZE-1:0] Wgt_3_320;input [WEIGHT_SIZE-1:0] Wgt_3_321;input [WEIGHT_SIZE-1:0] Wgt_3_322;input [WEIGHT_SIZE-1:0] Wgt_3_323;input [WEIGHT_SIZE-1:0] Wgt_3_324;input [WEIGHT_SIZE-1:0] Wgt_3_325;input [WEIGHT_SIZE-1:0] Wgt_3_326;input [WEIGHT_SIZE-1:0] Wgt_3_327;input [WEIGHT_SIZE-1:0] Wgt_3_328;input [WEIGHT_SIZE-1:0] Wgt_3_329;input [WEIGHT_SIZE-1:0] Wgt_3_330;input [WEIGHT_SIZE-1:0] Wgt_3_331;input [WEIGHT_SIZE-1:0] Wgt_3_332;input [WEIGHT_SIZE-1:0] Wgt_3_333;input [WEIGHT_SIZE-1:0] Wgt_3_334;input [WEIGHT_SIZE-1:0] Wgt_3_335;input [WEIGHT_SIZE-1:0] Wgt_3_336;input [WEIGHT_SIZE-1:0] Wgt_3_337;input [WEIGHT_SIZE-1:0] Wgt_3_338;input [WEIGHT_SIZE-1:0] Wgt_3_339;input [WEIGHT_SIZE-1:0] Wgt_3_340;input [WEIGHT_SIZE-1:0] Wgt_3_341;input [WEIGHT_SIZE-1:0] Wgt_3_342;input [WEIGHT_SIZE-1:0] Wgt_3_343;input [WEIGHT_SIZE-1:0] Wgt_3_344;input [WEIGHT_SIZE-1:0] Wgt_3_345;input [WEIGHT_SIZE-1:0] Wgt_3_346;input [WEIGHT_SIZE-1:0] Wgt_3_347;input [WEIGHT_SIZE-1:0] Wgt_3_348;input [WEIGHT_SIZE-1:0] Wgt_3_349;input [WEIGHT_SIZE-1:0] Wgt_3_350;input [WEIGHT_SIZE-1:0] Wgt_3_351;input [WEIGHT_SIZE-1:0] Wgt_3_352;input [WEIGHT_SIZE-1:0] Wgt_3_353;input [WEIGHT_SIZE-1:0] Wgt_3_354;input [WEIGHT_SIZE-1:0] Wgt_3_355;input [WEIGHT_SIZE-1:0] Wgt_3_356;input [WEIGHT_SIZE-1:0] Wgt_3_357;input [WEIGHT_SIZE-1:0] Wgt_3_358;input [WEIGHT_SIZE-1:0] Wgt_3_359;input [WEIGHT_SIZE-1:0] Wgt_3_360;input [WEIGHT_SIZE-1:0] Wgt_3_361;input [WEIGHT_SIZE-1:0] Wgt_3_362;input [WEIGHT_SIZE-1:0] Wgt_3_363;input [WEIGHT_SIZE-1:0] Wgt_3_364;input [WEIGHT_SIZE-1:0] Wgt_3_365;input [WEIGHT_SIZE-1:0] Wgt_3_366;input [WEIGHT_SIZE-1:0] Wgt_3_367;input [WEIGHT_SIZE-1:0] Wgt_3_368;input [WEIGHT_SIZE-1:0] Wgt_3_369;input [WEIGHT_SIZE-1:0] Wgt_3_370;input [WEIGHT_SIZE-1:0] Wgt_3_371;input [WEIGHT_SIZE-1:0] Wgt_3_372;input [WEIGHT_SIZE-1:0] Wgt_3_373;input [WEIGHT_SIZE-1:0] Wgt_3_374;input [WEIGHT_SIZE-1:0] Wgt_3_375;input [WEIGHT_SIZE-1:0] Wgt_3_376;input [WEIGHT_SIZE-1:0] Wgt_3_377;input [WEIGHT_SIZE-1:0] Wgt_3_378;input [WEIGHT_SIZE-1:0] Wgt_3_379;input [WEIGHT_SIZE-1:0] Wgt_3_380;input [WEIGHT_SIZE-1:0] Wgt_3_381;input [WEIGHT_SIZE-1:0] Wgt_3_382;input [WEIGHT_SIZE-1:0] Wgt_3_383;input [WEIGHT_SIZE-1:0] Wgt_3_384;input [WEIGHT_SIZE-1:0] Wgt_3_385;input [WEIGHT_SIZE-1:0] Wgt_3_386;input [WEIGHT_SIZE-1:0] Wgt_3_387;input [WEIGHT_SIZE-1:0] Wgt_3_388;input [WEIGHT_SIZE-1:0] Wgt_3_389;input [WEIGHT_SIZE-1:0] Wgt_3_390;input [WEIGHT_SIZE-1:0] Wgt_3_391;input [WEIGHT_SIZE-1:0] Wgt_3_392;input [WEIGHT_SIZE-1:0] Wgt_3_393;input [WEIGHT_SIZE-1:0] Wgt_3_394;input [WEIGHT_SIZE-1:0] Wgt_3_395;input [WEIGHT_SIZE-1:0] Wgt_3_396;input [WEIGHT_SIZE-1:0] Wgt_3_397;input [WEIGHT_SIZE-1:0] Wgt_3_398;input [WEIGHT_SIZE-1:0] Wgt_3_399;input [WEIGHT_SIZE-1:0] Wgt_3_400;input [WEIGHT_SIZE-1:0] Wgt_3_401;input [WEIGHT_SIZE-1:0] Wgt_3_402;input [WEIGHT_SIZE-1:0] Wgt_3_403;input [WEIGHT_SIZE-1:0] Wgt_3_404;input [WEIGHT_SIZE-1:0] Wgt_3_405;input [WEIGHT_SIZE-1:0] Wgt_3_406;input [WEIGHT_SIZE-1:0] Wgt_3_407;input [WEIGHT_SIZE-1:0] Wgt_3_408;input [WEIGHT_SIZE-1:0] Wgt_3_409;input [WEIGHT_SIZE-1:0] Wgt_3_410;input [WEIGHT_SIZE-1:0] Wgt_3_411;input [WEIGHT_SIZE-1:0] Wgt_3_412;input [WEIGHT_SIZE-1:0] Wgt_3_413;input [WEIGHT_SIZE-1:0] Wgt_3_414;input [WEIGHT_SIZE-1:0] Wgt_3_415;input [WEIGHT_SIZE-1:0] Wgt_3_416;input [WEIGHT_SIZE-1:0] Wgt_3_417;input [WEIGHT_SIZE-1:0] Wgt_3_418;input [WEIGHT_SIZE-1:0] Wgt_3_419;input [WEIGHT_SIZE-1:0] Wgt_3_420;input [WEIGHT_SIZE-1:0] Wgt_3_421;input [WEIGHT_SIZE-1:0] Wgt_3_422;input [WEIGHT_SIZE-1:0] Wgt_3_423;input [WEIGHT_SIZE-1:0] Wgt_3_424;input [WEIGHT_SIZE-1:0] Wgt_3_425;input [WEIGHT_SIZE-1:0] Wgt_3_426;input [WEIGHT_SIZE-1:0] Wgt_3_427;input [WEIGHT_SIZE-1:0] Wgt_3_428;input [WEIGHT_SIZE-1:0] Wgt_3_429;input [WEIGHT_SIZE-1:0] Wgt_3_430;input [WEIGHT_SIZE-1:0] Wgt_3_431;input [WEIGHT_SIZE-1:0] Wgt_3_432;input [WEIGHT_SIZE-1:0] Wgt_3_433;input [WEIGHT_SIZE-1:0] Wgt_3_434;input [WEIGHT_SIZE-1:0] Wgt_3_435;input [WEIGHT_SIZE-1:0] Wgt_3_436;input [WEIGHT_SIZE-1:0] Wgt_3_437;input [WEIGHT_SIZE-1:0] Wgt_3_438;input [WEIGHT_SIZE-1:0] Wgt_3_439;input [WEIGHT_SIZE-1:0] Wgt_3_440;input [WEIGHT_SIZE-1:0] Wgt_3_441;input [WEIGHT_SIZE-1:0] Wgt_3_442;input [WEIGHT_SIZE-1:0] Wgt_3_443;input [WEIGHT_SIZE-1:0] Wgt_3_444;input [WEIGHT_SIZE-1:0] Wgt_3_445;input [WEIGHT_SIZE-1:0] Wgt_3_446;input [WEIGHT_SIZE-1:0] Wgt_3_447;input [WEIGHT_SIZE-1:0] Wgt_3_448;input [WEIGHT_SIZE-1:0] Wgt_3_449;input [WEIGHT_SIZE-1:0] Wgt_3_450;input [WEIGHT_SIZE-1:0] Wgt_3_451;input [WEIGHT_SIZE-1:0] Wgt_3_452;input [WEIGHT_SIZE-1:0] Wgt_3_453;input [WEIGHT_SIZE-1:0] Wgt_3_454;input [WEIGHT_SIZE-1:0] Wgt_3_455;input [WEIGHT_SIZE-1:0] Wgt_3_456;input [WEIGHT_SIZE-1:0] Wgt_3_457;input [WEIGHT_SIZE-1:0] Wgt_3_458;input [WEIGHT_SIZE-1:0] Wgt_3_459;input [WEIGHT_SIZE-1:0] Wgt_3_460;input [WEIGHT_SIZE-1:0] Wgt_3_461;input [WEIGHT_SIZE-1:0] Wgt_3_462;input [WEIGHT_SIZE-1:0] Wgt_3_463;input [WEIGHT_SIZE-1:0] Wgt_3_464;input [WEIGHT_SIZE-1:0] Wgt_3_465;input [WEIGHT_SIZE-1:0] Wgt_3_466;input [WEIGHT_SIZE-1:0] Wgt_3_467;input [WEIGHT_SIZE-1:0] Wgt_3_468;input [WEIGHT_SIZE-1:0] Wgt_3_469;input [WEIGHT_SIZE-1:0] Wgt_3_470;input [WEIGHT_SIZE-1:0] Wgt_3_471;input [WEIGHT_SIZE-1:0] Wgt_3_472;input [WEIGHT_SIZE-1:0] Wgt_3_473;input [WEIGHT_SIZE-1:0] Wgt_3_474;input [WEIGHT_SIZE-1:0] Wgt_3_475;input [WEIGHT_SIZE-1:0] Wgt_3_476;input [WEIGHT_SIZE-1:0] Wgt_3_477;input [WEIGHT_SIZE-1:0] Wgt_3_478;input [WEIGHT_SIZE-1:0] Wgt_3_479;input [WEIGHT_SIZE-1:0] Wgt_3_480;input [WEIGHT_SIZE-1:0] Wgt_3_481;input [WEIGHT_SIZE-1:0] Wgt_3_482;input [WEIGHT_SIZE-1:0] Wgt_3_483;input [WEIGHT_SIZE-1:0] Wgt_3_484;input [WEIGHT_SIZE-1:0] Wgt_3_485;input [WEIGHT_SIZE-1:0] Wgt_3_486;input [WEIGHT_SIZE-1:0] Wgt_3_487;input [WEIGHT_SIZE-1:0] Wgt_3_488;input [WEIGHT_SIZE-1:0] Wgt_3_489;input [WEIGHT_SIZE-1:0] Wgt_3_490;input [WEIGHT_SIZE-1:0] Wgt_3_491;input [WEIGHT_SIZE-1:0] Wgt_3_492;input [WEIGHT_SIZE-1:0] Wgt_3_493;input [WEIGHT_SIZE-1:0] Wgt_3_494;input [WEIGHT_SIZE-1:0] Wgt_3_495;input [WEIGHT_SIZE-1:0] Wgt_3_496;input [WEIGHT_SIZE-1:0] Wgt_3_497;input [WEIGHT_SIZE-1:0] Wgt_3_498;input [WEIGHT_SIZE-1:0] Wgt_3_499;input [WEIGHT_SIZE-1:0] Wgt_3_500;input [WEIGHT_SIZE-1:0] Wgt_3_501;input [WEIGHT_SIZE-1:0] Wgt_3_502;input [WEIGHT_SIZE-1:0] Wgt_3_503;input [WEIGHT_SIZE-1:0] Wgt_3_504;input [WEIGHT_SIZE-1:0] Wgt_3_505;input [WEIGHT_SIZE-1:0] Wgt_3_506;input [WEIGHT_SIZE-1:0] Wgt_3_507;input [WEIGHT_SIZE-1:0] Wgt_3_508;input [WEIGHT_SIZE-1:0] Wgt_3_509;input [WEIGHT_SIZE-1:0] Wgt_3_510;input [WEIGHT_SIZE-1:0] Wgt_3_511;input [WEIGHT_SIZE-1:0] Wgt_3_512;input [WEIGHT_SIZE-1:0] Wgt_3_513;input [WEIGHT_SIZE-1:0] Wgt_3_514;input [WEIGHT_SIZE-1:0] Wgt_3_515;input [WEIGHT_SIZE-1:0] Wgt_3_516;input [WEIGHT_SIZE-1:0] Wgt_3_517;input [WEIGHT_SIZE-1:0] Wgt_3_518;input [WEIGHT_SIZE-1:0] Wgt_3_519;input [WEIGHT_SIZE-1:0] Wgt_3_520;input [WEIGHT_SIZE-1:0] Wgt_3_521;input [WEIGHT_SIZE-1:0] Wgt_3_522;input [WEIGHT_SIZE-1:0] Wgt_3_523;input [WEIGHT_SIZE-1:0] Wgt_3_524;input [WEIGHT_SIZE-1:0] Wgt_3_525;input [WEIGHT_SIZE-1:0] Wgt_3_526;input [WEIGHT_SIZE-1:0] Wgt_3_527;input [WEIGHT_SIZE-1:0] Wgt_3_528;input [WEIGHT_SIZE-1:0] Wgt_3_529;input [WEIGHT_SIZE-1:0] Wgt_3_530;input [WEIGHT_SIZE-1:0] Wgt_3_531;input [WEIGHT_SIZE-1:0] Wgt_3_532;input [WEIGHT_SIZE-1:0] Wgt_3_533;input [WEIGHT_SIZE-1:0] Wgt_3_534;input [WEIGHT_SIZE-1:0] Wgt_3_535;input [WEIGHT_SIZE-1:0] Wgt_3_536;input [WEIGHT_SIZE-1:0] Wgt_3_537;input [WEIGHT_SIZE-1:0] Wgt_3_538;input [WEIGHT_SIZE-1:0] Wgt_3_539;input [WEIGHT_SIZE-1:0] Wgt_3_540;input [WEIGHT_SIZE-1:0] Wgt_3_541;input [WEIGHT_SIZE-1:0] Wgt_3_542;input [WEIGHT_SIZE-1:0] Wgt_3_543;input [WEIGHT_SIZE-1:0] Wgt_3_544;input [WEIGHT_SIZE-1:0] Wgt_3_545;input [WEIGHT_SIZE-1:0] Wgt_3_546;input [WEIGHT_SIZE-1:0] Wgt_3_547;input [WEIGHT_SIZE-1:0] Wgt_3_548;input [WEIGHT_SIZE-1:0] Wgt_3_549;input [WEIGHT_SIZE-1:0] Wgt_3_550;input [WEIGHT_SIZE-1:0] Wgt_3_551;input [WEIGHT_SIZE-1:0] Wgt_3_552;input [WEIGHT_SIZE-1:0] Wgt_3_553;input [WEIGHT_SIZE-1:0] Wgt_3_554;input [WEIGHT_SIZE-1:0] Wgt_3_555;input [WEIGHT_SIZE-1:0] Wgt_3_556;input [WEIGHT_SIZE-1:0] Wgt_3_557;input [WEIGHT_SIZE-1:0] Wgt_3_558;input [WEIGHT_SIZE-1:0] Wgt_3_559;input [WEIGHT_SIZE-1:0] Wgt_3_560;input [WEIGHT_SIZE-1:0] Wgt_3_561;input [WEIGHT_SIZE-1:0] Wgt_3_562;input [WEIGHT_SIZE-1:0] Wgt_3_563;input [WEIGHT_SIZE-1:0] Wgt_3_564;input [WEIGHT_SIZE-1:0] Wgt_3_565;input [WEIGHT_SIZE-1:0] Wgt_3_566;input [WEIGHT_SIZE-1:0] Wgt_3_567;input [WEIGHT_SIZE-1:0] Wgt_3_568;input [WEIGHT_SIZE-1:0] Wgt_3_569;input [WEIGHT_SIZE-1:0] Wgt_3_570;input [WEIGHT_SIZE-1:0] Wgt_3_571;input [WEIGHT_SIZE-1:0] Wgt_3_572;input [WEIGHT_SIZE-1:0] Wgt_3_573;input [WEIGHT_SIZE-1:0] Wgt_3_574;input [WEIGHT_SIZE-1:0] Wgt_3_575;input [WEIGHT_SIZE-1:0] Wgt_3_576;input [WEIGHT_SIZE-1:0] Wgt_3_577;input [WEIGHT_SIZE-1:0] Wgt_3_578;input [WEIGHT_SIZE-1:0] Wgt_3_579;input [WEIGHT_SIZE-1:0] Wgt_3_580;input [WEIGHT_SIZE-1:0] Wgt_3_581;input [WEIGHT_SIZE-1:0] Wgt_3_582;input [WEIGHT_SIZE-1:0] Wgt_3_583;input [WEIGHT_SIZE-1:0] Wgt_3_584;input [WEIGHT_SIZE-1:0] Wgt_3_585;input [WEIGHT_SIZE-1:0] Wgt_3_586;input [WEIGHT_SIZE-1:0] Wgt_3_587;input [WEIGHT_SIZE-1:0] Wgt_3_588;input [WEIGHT_SIZE-1:0] Wgt_3_589;input [WEIGHT_SIZE-1:0] Wgt_3_590;input [WEIGHT_SIZE-1:0] Wgt_3_591;input [WEIGHT_SIZE-1:0] Wgt_3_592;input [WEIGHT_SIZE-1:0] Wgt_3_593;input [WEIGHT_SIZE-1:0] Wgt_3_594;input [WEIGHT_SIZE-1:0] Wgt_3_595;input [WEIGHT_SIZE-1:0] Wgt_3_596;input [WEIGHT_SIZE-1:0] Wgt_3_597;input [WEIGHT_SIZE-1:0] Wgt_3_598;input [WEIGHT_SIZE-1:0] Wgt_3_599;input [WEIGHT_SIZE-1:0] Wgt_3_600;input [WEIGHT_SIZE-1:0] Wgt_3_601;input [WEIGHT_SIZE-1:0] Wgt_3_602;input [WEIGHT_SIZE-1:0] Wgt_3_603;input [WEIGHT_SIZE-1:0] Wgt_3_604;input [WEIGHT_SIZE-1:0] Wgt_3_605;input [WEIGHT_SIZE-1:0] Wgt_3_606;input [WEIGHT_SIZE-1:0] Wgt_3_607;input [WEIGHT_SIZE-1:0] Wgt_3_608;input [WEIGHT_SIZE-1:0] Wgt_3_609;input [WEIGHT_SIZE-1:0] Wgt_3_610;input [WEIGHT_SIZE-1:0] Wgt_3_611;input [WEIGHT_SIZE-1:0] Wgt_3_612;input [WEIGHT_SIZE-1:0] Wgt_3_613;input [WEIGHT_SIZE-1:0] Wgt_3_614;input [WEIGHT_SIZE-1:0] Wgt_3_615;input [WEIGHT_SIZE-1:0] Wgt_3_616;input [WEIGHT_SIZE-1:0] Wgt_3_617;input [WEIGHT_SIZE-1:0] Wgt_3_618;input [WEIGHT_SIZE-1:0] Wgt_3_619;input [WEIGHT_SIZE-1:0] Wgt_3_620;input [WEIGHT_SIZE-1:0] Wgt_3_621;input [WEIGHT_SIZE-1:0] Wgt_3_622;input [WEIGHT_SIZE-1:0] Wgt_3_623;input [WEIGHT_SIZE-1:0] Wgt_3_624;input [WEIGHT_SIZE-1:0] Wgt_3_625;input [WEIGHT_SIZE-1:0] Wgt_3_626;input [WEIGHT_SIZE-1:0] Wgt_3_627;input [WEIGHT_SIZE-1:0] Wgt_3_628;input [WEIGHT_SIZE-1:0] Wgt_3_629;input [WEIGHT_SIZE-1:0] Wgt_3_630;input [WEIGHT_SIZE-1:0] Wgt_3_631;input [WEIGHT_SIZE-1:0] Wgt_3_632;input [WEIGHT_SIZE-1:0] Wgt_3_633;input [WEIGHT_SIZE-1:0] Wgt_3_634;input [WEIGHT_SIZE-1:0] Wgt_3_635;input [WEIGHT_SIZE-1:0] Wgt_3_636;input [WEIGHT_SIZE-1:0] Wgt_3_637;input [WEIGHT_SIZE-1:0] Wgt_3_638;input [WEIGHT_SIZE-1:0] Wgt_3_639;input [WEIGHT_SIZE-1:0] Wgt_3_640;input [WEIGHT_SIZE-1:0] Wgt_3_641;input [WEIGHT_SIZE-1:0] Wgt_3_642;input [WEIGHT_SIZE-1:0] Wgt_3_643;input [WEIGHT_SIZE-1:0] Wgt_3_644;input [WEIGHT_SIZE-1:0] Wgt_3_645;input [WEIGHT_SIZE-1:0] Wgt_3_646;input [WEIGHT_SIZE-1:0] Wgt_3_647;input [WEIGHT_SIZE-1:0] Wgt_3_648;input [WEIGHT_SIZE-1:0] Wgt_3_649;input [WEIGHT_SIZE-1:0] Wgt_3_650;input [WEIGHT_SIZE-1:0] Wgt_3_651;input [WEIGHT_SIZE-1:0] Wgt_3_652;input [WEIGHT_SIZE-1:0] Wgt_3_653;input [WEIGHT_SIZE-1:0] Wgt_3_654;input [WEIGHT_SIZE-1:0] Wgt_3_655;input [WEIGHT_SIZE-1:0] Wgt_3_656;input [WEIGHT_SIZE-1:0] Wgt_3_657;input [WEIGHT_SIZE-1:0] Wgt_3_658;input [WEIGHT_SIZE-1:0] Wgt_3_659;input [WEIGHT_SIZE-1:0] Wgt_3_660;input [WEIGHT_SIZE-1:0] Wgt_3_661;input [WEIGHT_SIZE-1:0] Wgt_3_662;input [WEIGHT_SIZE-1:0] Wgt_3_663;input [WEIGHT_SIZE-1:0] Wgt_3_664;input [WEIGHT_SIZE-1:0] Wgt_3_665;input [WEIGHT_SIZE-1:0] Wgt_3_666;input [WEIGHT_SIZE-1:0] Wgt_3_667;input [WEIGHT_SIZE-1:0] Wgt_3_668;input [WEIGHT_SIZE-1:0] Wgt_3_669;input [WEIGHT_SIZE-1:0] Wgt_3_670;input [WEIGHT_SIZE-1:0] Wgt_3_671;input [WEIGHT_SIZE-1:0] Wgt_3_672;input [WEIGHT_SIZE-1:0] Wgt_3_673;input [WEIGHT_SIZE-1:0] Wgt_3_674;input [WEIGHT_SIZE-1:0] Wgt_3_675;input [WEIGHT_SIZE-1:0] Wgt_3_676;input [WEIGHT_SIZE-1:0] Wgt_3_677;input [WEIGHT_SIZE-1:0] Wgt_3_678;input [WEIGHT_SIZE-1:0] Wgt_3_679;input [WEIGHT_SIZE-1:0] Wgt_3_680;input [WEIGHT_SIZE-1:0] Wgt_3_681;input [WEIGHT_SIZE-1:0] Wgt_3_682;input [WEIGHT_SIZE-1:0] Wgt_3_683;input [WEIGHT_SIZE-1:0] Wgt_3_684;input [WEIGHT_SIZE-1:0] Wgt_3_685;input [WEIGHT_SIZE-1:0] Wgt_3_686;input [WEIGHT_SIZE-1:0] Wgt_3_687;input [WEIGHT_SIZE-1:0] Wgt_3_688;input [WEIGHT_SIZE-1:0] Wgt_3_689;input [WEIGHT_SIZE-1:0] Wgt_3_690;input [WEIGHT_SIZE-1:0] Wgt_3_691;input [WEIGHT_SIZE-1:0] Wgt_3_692;input [WEIGHT_SIZE-1:0] Wgt_3_693;input [WEIGHT_SIZE-1:0] Wgt_3_694;input [WEIGHT_SIZE-1:0] Wgt_3_695;input [WEIGHT_SIZE-1:0] Wgt_3_696;input [WEIGHT_SIZE-1:0] Wgt_3_697;input [WEIGHT_SIZE-1:0] Wgt_3_698;input [WEIGHT_SIZE-1:0] Wgt_3_699;input [WEIGHT_SIZE-1:0] Wgt_3_700;input [WEIGHT_SIZE-1:0] Wgt_3_701;input [WEIGHT_SIZE-1:0] Wgt_3_702;input [WEIGHT_SIZE-1:0] Wgt_3_703;input [WEIGHT_SIZE-1:0] Wgt_3_704;input [WEIGHT_SIZE-1:0] Wgt_3_705;input [WEIGHT_SIZE-1:0] Wgt_3_706;input [WEIGHT_SIZE-1:0] Wgt_3_707;input [WEIGHT_SIZE-1:0] Wgt_3_708;input [WEIGHT_SIZE-1:0] Wgt_3_709;input [WEIGHT_SIZE-1:0] Wgt_3_710;input [WEIGHT_SIZE-1:0] Wgt_3_711;input [WEIGHT_SIZE-1:0] Wgt_3_712;input [WEIGHT_SIZE-1:0] Wgt_3_713;input [WEIGHT_SIZE-1:0] Wgt_3_714;input [WEIGHT_SIZE-1:0] Wgt_3_715;input [WEIGHT_SIZE-1:0] Wgt_3_716;input [WEIGHT_SIZE-1:0] Wgt_3_717;input [WEIGHT_SIZE-1:0] Wgt_3_718;input [WEIGHT_SIZE-1:0] Wgt_3_719;input [WEIGHT_SIZE-1:0] Wgt_3_720;input [WEIGHT_SIZE-1:0] Wgt_3_721;input [WEIGHT_SIZE-1:0] Wgt_3_722;input [WEIGHT_SIZE-1:0] Wgt_3_723;input [WEIGHT_SIZE-1:0] Wgt_3_724;input [WEIGHT_SIZE-1:0] Wgt_3_725;input [WEIGHT_SIZE-1:0] Wgt_3_726;input [WEIGHT_SIZE-1:0] Wgt_3_727;input [WEIGHT_SIZE-1:0] Wgt_3_728;input [WEIGHT_SIZE-1:0] Wgt_3_729;input [WEIGHT_SIZE-1:0] Wgt_3_730;input [WEIGHT_SIZE-1:0] Wgt_3_731;input [WEIGHT_SIZE-1:0] Wgt_3_732;input [WEIGHT_SIZE-1:0] Wgt_3_733;input [WEIGHT_SIZE-1:0] Wgt_3_734;input [WEIGHT_SIZE-1:0] Wgt_3_735;input [WEIGHT_SIZE-1:0] Wgt_3_736;input [WEIGHT_SIZE-1:0] Wgt_3_737;input [WEIGHT_SIZE-1:0] Wgt_3_738;input [WEIGHT_SIZE-1:0] Wgt_3_739;input [WEIGHT_SIZE-1:0] Wgt_3_740;input [WEIGHT_SIZE-1:0] Wgt_3_741;input [WEIGHT_SIZE-1:0] Wgt_3_742;input [WEIGHT_SIZE-1:0] Wgt_3_743;input [WEIGHT_SIZE-1:0] Wgt_3_744;input [WEIGHT_SIZE-1:0] Wgt_3_745;input [WEIGHT_SIZE-1:0] Wgt_3_746;input [WEIGHT_SIZE-1:0] Wgt_3_747;input [WEIGHT_SIZE-1:0] Wgt_3_748;input [WEIGHT_SIZE-1:0] Wgt_3_749;input [WEIGHT_SIZE-1:0] Wgt_3_750;input [WEIGHT_SIZE-1:0] Wgt_3_751;input [WEIGHT_SIZE-1:0] Wgt_3_752;input [WEIGHT_SIZE-1:0] Wgt_3_753;input [WEIGHT_SIZE-1:0] Wgt_3_754;input [WEIGHT_SIZE-1:0] Wgt_3_755;input [WEIGHT_SIZE-1:0] Wgt_3_756;input [WEIGHT_SIZE-1:0] Wgt_3_757;input [WEIGHT_SIZE-1:0] Wgt_3_758;input [WEIGHT_SIZE-1:0] Wgt_3_759;input [WEIGHT_SIZE-1:0] Wgt_3_760;input [WEIGHT_SIZE-1:0] Wgt_3_761;input [WEIGHT_SIZE-1:0] Wgt_3_762;input [WEIGHT_SIZE-1:0] Wgt_3_763;input [WEIGHT_SIZE-1:0] Wgt_3_764;input [WEIGHT_SIZE-1:0] Wgt_3_765;input [WEIGHT_SIZE-1:0] Wgt_3_766;input [WEIGHT_SIZE-1:0] Wgt_3_767;input [WEIGHT_SIZE-1:0] Wgt_3_768;input [WEIGHT_SIZE-1:0] Wgt_3_769;input [WEIGHT_SIZE-1:0] Wgt_3_770;input [WEIGHT_SIZE-1:0] Wgt_3_771;input [WEIGHT_SIZE-1:0] Wgt_3_772;input [WEIGHT_SIZE-1:0] Wgt_3_773;input [WEIGHT_SIZE-1:0] Wgt_3_774;input [WEIGHT_SIZE-1:0] Wgt_3_775;input [WEIGHT_SIZE-1:0] Wgt_3_776;input [WEIGHT_SIZE-1:0] Wgt_3_777;input [WEIGHT_SIZE-1:0] Wgt_3_778;input [WEIGHT_SIZE-1:0] Wgt_3_779;input [WEIGHT_SIZE-1:0] Wgt_3_780;input [WEIGHT_SIZE-1:0] Wgt_3_781;input [WEIGHT_SIZE-1:0] Wgt_3_782;input [WEIGHT_SIZE-1:0] Wgt_3_783;input [WEIGHT_SIZE-1:0] Wgt_3_784;input [WEIGHT_SIZE-1:0] Wgt_4_0;input [WEIGHT_SIZE-1:0] Wgt_4_1;input [WEIGHT_SIZE-1:0] Wgt_4_2;input [WEIGHT_SIZE-1:0] Wgt_4_3;input [WEIGHT_SIZE-1:0] Wgt_4_4;input [WEIGHT_SIZE-1:0] Wgt_4_5;input [WEIGHT_SIZE-1:0] Wgt_4_6;input [WEIGHT_SIZE-1:0] Wgt_4_7;input [WEIGHT_SIZE-1:0] Wgt_4_8;input [WEIGHT_SIZE-1:0] Wgt_4_9;input [WEIGHT_SIZE-1:0] Wgt_4_10;input [WEIGHT_SIZE-1:0] Wgt_4_11;input [WEIGHT_SIZE-1:0] Wgt_4_12;input [WEIGHT_SIZE-1:0] Wgt_4_13;input [WEIGHT_SIZE-1:0] Wgt_4_14;input [WEIGHT_SIZE-1:0] Wgt_4_15;input [WEIGHT_SIZE-1:0] Wgt_4_16;input [WEIGHT_SIZE-1:0] Wgt_4_17;input [WEIGHT_SIZE-1:0] Wgt_4_18;input [WEIGHT_SIZE-1:0] Wgt_4_19;input [WEIGHT_SIZE-1:0] Wgt_4_20;input [WEIGHT_SIZE-1:0] Wgt_4_21;input [WEIGHT_SIZE-1:0] Wgt_4_22;input [WEIGHT_SIZE-1:0] Wgt_4_23;input [WEIGHT_SIZE-1:0] Wgt_4_24;input [WEIGHT_SIZE-1:0] Wgt_4_25;input [WEIGHT_SIZE-1:0] Wgt_4_26;input [WEIGHT_SIZE-1:0] Wgt_4_27;input [WEIGHT_SIZE-1:0] Wgt_4_28;input [WEIGHT_SIZE-1:0] Wgt_4_29;input [WEIGHT_SIZE-1:0] Wgt_4_30;input [WEIGHT_SIZE-1:0] Wgt_4_31;input [WEIGHT_SIZE-1:0] Wgt_4_32;input [WEIGHT_SIZE-1:0] Wgt_4_33;input [WEIGHT_SIZE-1:0] Wgt_4_34;input [WEIGHT_SIZE-1:0] Wgt_4_35;input [WEIGHT_SIZE-1:0] Wgt_4_36;input [WEIGHT_SIZE-1:0] Wgt_4_37;input [WEIGHT_SIZE-1:0] Wgt_4_38;input [WEIGHT_SIZE-1:0] Wgt_4_39;input [WEIGHT_SIZE-1:0] Wgt_4_40;input [WEIGHT_SIZE-1:0] Wgt_4_41;input [WEIGHT_SIZE-1:0] Wgt_4_42;input [WEIGHT_SIZE-1:0] Wgt_4_43;input [WEIGHT_SIZE-1:0] Wgt_4_44;input [WEIGHT_SIZE-1:0] Wgt_4_45;input [WEIGHT_SIZE-1:0] Wgt_4_46;input [WEIGHT_SIZE-1:0] Wgt_4_47;input [WEIGHT_SIZE-1:0] Wgt_4_48;input [WEIGHT_SIZE-1:0] Wgt_4_49;input [WEIGHT_SIZE-1:0] Wgt_4_50;input [WEIGHT_SIZE-1:0] Wgt_4_51;input [WEIGHT_SIZE-1:0] Wgt_4_52;input [WEIGHT_SIZE-1:0] Wgt_4_53;input [WEIGHT_SIZE-1:0] Wgt_4_54;input [WEIGHT_SIZE-1:0] Wgt_4_55;input [WEIGHT_SIZE-1:0] Wgt_4_56;input [WEIGHT_SIZE-1:0] Wgt_4_57;input [WEIGHT_SIZE-1:0] Wgt_4_58;input [WEIGHT_SIZE-1:0] Wgt_4_59;input [WEIGHT_SIZE-1:0] Wgt_4_60;input [WEIGHT_SIZE-1:0] Wgt_4_61;input [WEIGHT_SIZE-1:0] Wgt_4_62;input [WEIGHT_SIZE-1:0] Wgt_4_63;input [WEIGHT_SIZE-1:0] Wgt_4_64;input [WEIGHT_SIZE-1:0] Wgt_4_65;input [WEIGHT_SIZE-1:0] Wgt_4_66;input [WEIGHT_SIZE-1:0] Wgt_4_67;input [WEIGHT_SIZE-1:0] Wgt_4_68;input [WEIGHT_SIZE-1:0] Wgt_4_69;input [WEIGHT_SIZE-1:0] Wgt_4_70;input [WEIGHT_SIZE-1:0] Wgt_4_71;input [WEIGHT_SIZE-1:0] Wgt_4_72;input [WEIGHT_SIZE-1:0] Wgt_4_73;input [WEIGHT_SIZE-1:0] Wgt_4_74;input [WEIGHT_SIZE-1:0] Wgt_4_75;input [WEIGHT_SIZE-1:0] Wgt_4_76;input [WEIGHT_SIZE-1:0] Wgt_4_77;input [WEIGHT_SIZE-1:0] Wgt_4_78;input [WEIGHT_SIZE-1:0] Wgt_4_79;input [WEIGHT_SIZE-1:0] Wgt_4_80;input [WEIGHT_SIZE-1:0] Wgt_4_81;input [WEIGHT_SIZE-1:0] Wgt_4_82;input [WEIGHT_SIZE-1:0] Wgt_4_83;input [WEIGHT_SIZE-1:0] Wgt_4_84;input [WEIGHT_SIZE-1:0] Wgt_4_85;input [WEIGHT_SIZE-1:0] Wgt_4_86;input [WEIGHT_SIZE-1:0] Wgt_4_87;input [WEIGHT_SIZE-1:0] Wgt_4_88;input [WEIGHT_SIZE-1:0] Wgt_4_89;input [WEIGHT_SIZE-1:0] Wgt_4_90;input [WEIGHT_SIZE-1:0] Wgt_4_91;input [WEIGHT_SIZE-1:0] Wgt_4_92;input [WEIGHT_SIZE-1:0] Wgt_4_93;input [WEIGHT_SIZE-1:0] Wgt_4_94;input [WEIGHT_SIZE-1:0] Wgt_4_95;input [WEIGHT_SIZE-1:0] Wgt_4_96;input [WEIGHT_SIZE-1:0] Wgt_4_97;input [WEIGHT_SIZE-1:0] Wgt_4_98;input [WEIGHT_SIZE-1:0] Wgt_4_99;input [WEIGHT_SIZE-1:0] Wgt_4_100;input [WEIGHT_SIZE-1:0] Wgt_4_101;input [WEIGHT_SIZE-1:0] Wgt_4_102;input [WEIGHT_SIZE-1:0] Wgt_4_103;input [WEIGHT_SIZE-1:0] Wgt_4_104;input [WEIGHT_SIZE-1:0] Wgt_4_105;input [WEIGHT_SIZE-1:0] Wgt_4_106;input [WEIGHT_SIZE-1:0] Wgt_4_107;input [WEIGHT_SIZE-1:0] Wgt_4_108;input [WEIGHT_SIZE-1:0] Wgt_4_109;input [WEIGHT_SIZE-1:0] Wgt_4_110;input [WEIGHT_SIZE-1:0] Wgt_4_111;input [WEIGHT_SIZE-1:0] Wgt_4_112;input [WEIGHT_SIZE-1:0] Wgt_4_113;input [WEIGHT_SIZE-1:0] Wgt_4_114;input [WEIGHT_SIZE-1:0] Wgt_4_115;input [WEIGHT_SIZE-1:0] Wgt_4_116;input [WEIGHT_SIZE-1:0] Wgt_4_117;input [WEIGHT_SIZE-1:0] Wgt_4_118;input [WEIGHT_SIZE-1:0] Wgt_4_119;input [WEIGHT_SIZE-1:0] Wgt_4_120;input [WEIGHT_SIZE-1:0] Wgt_4_121;input [WEIGHT_SIZE-1:0] Wgt_4_122;input [WEIGHT_SIZE-1:0] Wgt_4_123;input [WEIGHT_SIZE-1:0] Wgt_4_124;input [WEIGHT_SIZE-1:0] Wgt_4_125;input [WEIGHT_SIZE-1:0] Wgt_4_126;input [WEIGHT_SIZE-1:0] Wgt_4_127;input [WEIGHT_SIZE-1:0] Wgt_4_128;input [WEIGHT_SIZE-1:0] Wgt_4_129;input [WEIGHT_SIZE-1:0] Wgt_4_130;input [WEIGHT_SIZE-1:0] Wgt_4_131;input [WEIGHT_SIZE-1:0] Wgt_4_132;input [WEIGHT_SIZE-1:0] Wgt_4_133;input [WEIGHT_SIZE-1:0] Wgt_4_134;input [WEIGHT_SIZE-1:0] Wgt_4_135;input [WEIGHT_SIZE-1:0] Wgt_4_136;input [WEIGHT_SIZE-1:0] Wgt_4_137;input [WEIGHT_SIZE-1:0] Wgt_4_138;input [WEIGHT_SIZE-1:0] Wgt_4_139;input [WEIGHT_SIZE-1:0] Wgt_4_140;input [WEIGHT_SIZE-1:0] Wgt_4_141;input [WEIGHT_SIZE-1:0] Wgt_4_142;input [WEIGHT_SIZE-1:0] Wgt_4_143;input [WEIGHT_SIZE-1:0] Wgt_4_144;input [WEIGHT_SIZE-1:0] Wgt_4_145;input [WEIGHT_SIZE-1:0] Wgt_4_146;input [WEIGHT_SIZE-1:0] Wgt_4_147;input [WEIGHT_SIZE-1:0] Wgt_4_148;input [WEIGHT_SIZE-1:0] Wgt_4_149;input [WEIGHT_SIZE-1:0] Wgt_4_150;input [WEIGHT_SIZE-1:0] Wgt_4_151;input [WEIGHT_SIZE-1:0] Wgt_4_152;input [WEIGHT_SIZE-1:0] Wgt_4_153;input [WEIGHT_SIZE-1:0] Wgt_4_154;input [WEIGHT_SIZE-1:0] Wgt_4_155;input [WEIGHT_SIZE-1:0] Wgt_4_156;input [WEIGHT_SIZE-1:0] Wgt_4_157;input [WEIGHT_SIZE-1:0] Wgt_4_158;input [WEIGHT_SIZE-1:0] Wgt_4_159;input [WEIGHT_SIZE-1:0] Wgt_4_160;input [WEIGHT_SIZE-1:0] Wgt_4_161;input [WEIGHT_SIZE-1:0] Wgt_4_162;input [WEIGHT_SIZE-1:0] Wgt_4_163;input [WEIGHT_SIZE-1:0] Wgt_4_164;input [WEIGHT_SIZE-1:0] Wgt_4_165;input [WEIGHT_SIZE-1:0] Wgt_4_166;input [WEIGHT_SIZE-1:0] Wgt_4_167;input [WEIGHT_SIZE-1:0] Wgt_4_168;input [WEIGHT_SIZE-1:0] Wgt_4_169;input [WEIGHT_SIZE-1:0] Wgt_4_170;input [WEIGHT_SIZE-1:0] Wgt_4_171;input [WEIGHT_SIZE-1:0] Wgt_4_172;input [WEIGHT_SIZE-1:0] Wgt_4_173;input [WEIGHT_SIZE-1:0] Wgt_4_174;input [WEIGHT_SIZE-1:0] Wgt_4_175;input [WEIGHT_SIZE-1:0] Wgt_4_176;input [WEIGHT_SIZE-1:0] Wgt_4_177;input [WEIGHT_SIZE-1:0] Wgt_4_178;input [WEIGHT_SIZE-1:0] Wgt_4_179;input [WEIGHT_SIZE-1:0] Wgt_4_180;input [WEIGHT_SIZE-1:0] Wgt_4_181;input [WEIGHT_SIZE-1:0] Wgt_4_182;input [WEIGHT_SIZE-1:0] Wgt_4_183;input [WEIGHT_SIZE-1:0] Wgt_4_184;input [WEIGHT_SIZE-1:0] Wgt_4_185;input [WEIGHT_SIZE-1:0] Wgt_4_186;input [WEIGHT_SIZE-1:0] Wgt_4_187;input [WEIGHT_SIZE-1:0] Wgt_4_188;input [WEIGHT_SIZE-1:0] Wgt_4_189;input [WEIGHT_SIZE-1:0] Wgt_4_190;input [WEIGHT_SIZE-1:0] Wgt_4_191;input [WEIGHT_SIZE-1:0] Wgt_4_192;input [WEIGHT_SIZE-1:0] Wgt_4_193;input [WEIGHT_SIZE-1:0] Wgt_4_194;input [WEIGHT_SIZE-1:0] Wgt_4_195;input [WEIGHT_SIZE-1:0] Wgt_4_196;input [WEIGHT_SIZE-1:0] Wgt_4_197;input [WEIGHT_SIZE-1:0] Wgt_4_198;input [WEIGHT_SIZE-1:0] Wgt_4_199;input [WEIGHT_SIZE-1:0] Wgt_4_200;input [WEIGHT_SIZE-1:0] Wgt_4_201;input [WEIGHT_SIZE-1:0] Wgt_4_202;input [WEIGHT_SIZE-1:0] Wgt_4_203;input [WEIGHT_SIZE-1:0] Wgt_4_204;input [WEIGHT_SIZE-1:0] Wgt_4_205;input [WEIGHT_SIZE-1:0] Wgt_4_206;input [WEIGHT_SIZE-1:0] Wgt_4_207;input [WEIGHT_SIZE-1:0] Wgt_4_208;input [WEIGHT_SIZE-1:0] Wgt_4_209;input [WEIGHT_SIZE-1:0] Wgt_4_210;input [WEIGHT_SIZE-1:0] Wgt_4_211;input [WEIGHT_SIZE-1:0] Wgt_4_212;input [WEIGHT_SIZE-1:0] Wgt_4_213;input [WEIGHT_SIZE-1:0] Wgt_4_214;input [WEIGHT_SIZE-1:0] Wgt_4_215;input [WEIGHT_SIZE-1:0] Wgt_4_216;input [WEIGHT_SIZE-1:0] Wgt_4_217;input [WEIGHT_SIZE-1:0] Wgt_4_218;input [WEIGHT_SIZE-1:0] Wgt_4_219;input [WEIGHT_SIZE-1:0] Wgt_4_220;input [WEIGHT_SIZE-1:0] Wgt_4_221;input [WEIGHT_SIZE-1:0] Wgt_4_222;input [WEIGHT_SIZE-1:0] Wgt_4_223;input [WEIGHT_SIZE-1:0] Wgt_4_224;input [WEIGHT_SIZE-1:0] Wgt_4_225;input [WEIGHT_SIZE-1:0] Wgt_4_226;input [WEIGHT_SIZE-1:0] Wgt_4_227;input [WEIGHT_SIZE-1:0] Wgt_4_228;input [WEIGHT_SIZE-1:0] Wgt_4_229;input [WEIGHT_SIZE-1:0] Wgt_4_230;input [WEIGHT_SIZE-1:0] Wgt_4_231;input [WEIGHT_SIZE-1:0] Wgt_4_232;input [WEIGHT_SIZE-1:0] Wgt_4_233;input [WEIGHT_SIZE-1:0] Wgt_4_234;input [WEIGHT_SIZE-1:0] Wgt_4_235;input [WEIGHT_SIZE-1:0] Wgt_4_236;input [WEIGHT_SIZE-1:0] Wgt_4_237;input [WEIGHT_SIZE-1:0] Wgt_4_238;input [WEIGHT_SIZE-1:0] Wgt_4_239;input [WEIGHT_SIZE-1:0] Wgt_4_240;input [WEIGHT_SIZE-1:0] Wgt_4_241;input [WEIGHT_SIZE-1:0] Wgt_4_242;input [WEIGHT_SIZE-1:0] Wgt_4_243;input [WEIGHT_SIZE-1:0] Wgt_4_244;input [WEIGHT_SIZE-1:0] Wgt_4_245;input [WEIGHT_SIZE-1:0] Wgt_4_246;input [WEIGHT_SIZE-1:0] Wgt_4_247;input [WEIGHT_SIZE-1:0] Wgt_4_248;input [WEIGHT_SIZE-1:0] Wgt_4_249;input [WEIGHT_SIZE-1:0] Wgt_4_250;input [WEIGHT_SIZE-1:0] Wgt_4_251;input [WEIGHT_SIZE-1:0] Wgt_4_252;input [WEIGHT_SIZE-1:0] Wgt_4_253;input [WEIGHT_SIZE-1:0] Wgt_4_254;input [WEIGHT_SIZE-1:0] Wgt_4_255;input [WEIGHT_SIZE-1:0] Wgt_4_256;input [WEIGHT_SIZE-1:0] Wgt_4_257;input [WEIGHT_SIZE-1:0] Wgt_4_258;input [WEIGHT_SIZE-1:0] Wgt_4_259;input [WEIGHT_SIZE-1:0] Wgt_4_260;input [WEIGHT_SIZE-1:0] Wgt_4_261;input [WEIGHT_SIZE-1:0] Wgt_4_262;input [WEIGHT_SIZE-1:0] Wgt_4_263;input [WEIGHT_SIZE-1:0] Wgt_4_264;input [WEIGHT_SIZE-1:0] Wgt_4_265;input [WEIGHT_SIZE-1:0] Wgt_4_266;input [WEIGHT_SIZE-1:0] Wgt_4_267;input [WEIGHT_SIZE-1:0] Wgt_4_268;input [WEIGHT_SIZE-1:0] Wgt_4_269;input [WEIGHT_SIZE-1:0] Wgt_4_270;input [WEIGHT_SIZE-1:0] Wgt_4_271;input [WEIGHT_SIZE-1:0] Wgt_4_272;input [WEIGHT_SIZE-1:0] Wgt_4_273;input [WEIGHT_SIZE-1:0] Wgt_4_274;input [WEIGHT_SIZE-1:0] Wgt_4_275;input [WEIGHT_SIZE-1:0] Wgt_4_276;input [WEIGHT_SIZE-1:0] Wgt_4_277;input [WEIGHT_SIZE-1:0] Wgt_4_278;input [WEIGHT_SIZE-1:0] Wgt_4_279;input [WEIGHT_SIZE-1:0] Wgt_4_280;input [WEIGHT_SIZE-1:0] Wgt_4_281;input [WEIGHT_SIZE-1:0] Wgt_4_282;input [WEIGHT_SIZE-1:0] Wgt_4_283;input [WEIGHT_SIZE-1:0] Wgt_4_284;input [WEIGHT_SIZE-1:0] Wgt_4_285;input [WEIGHT_SIZE-1:0] Wgt_4_286;input [WEIGHT_SIZE-1:0] Wgt_4_287;input [WEIGHT_SIZE-1:0] Wgt_4_288;input [WEIGHT_SIZE-1:0] Wgt_4_289;input [WEIGHT_SIZE-1:0] Wgt_4_290;input [WEIGHT_SIZE-1:0] Wgt_4_291;input [WEIGHT_SIZE-1:0] Wgt_4_292;input [WEIGHT_SIZE-1:0] Wgt_4_293;input [WEIGHT_SIZE-1:0] Wgt_4_294;input [WEIGHT_SIZE-1:0] Wgt_4_295;input [WEIGHT_SIZE-1:0] Wgt_4_296;input [WEIGHT_SIZE-1:0] Wgt_4_297;input [WEIGHT_SIZE-1:0] Wgt_4_298;input [WEIGHT_SIZE-1:0] Wgt_4_299;input [WEIGHT_SIZE-1:0] Wgt_4_300;input [WEIGHT_SIZE-1:0] Wgt_4_301;input [WEIGHT_SIZE-1:0] Wgt_4_302;input [WEIGHT_SIZE-1:0] Wgt_4_303;input [WEIGHT_SIZE-1:0] Wgt_4_304;input [WEIGHT_SIZE-1:0] Wgt_4_305;input [WEIGHT_SIZE-1:0] Wgt_4_306;input [WEIGHT_SIZE-1:0] Wgt_4_307;input [WEIGHT_SIZE-1:0] Wgt_4_308;input [WEIGHT_SIZE-1:0] Wgt_4_309;input [WEIGHT_SIZE-1:0] Wgt_4_310;input [WEIGHT_SIZE-1:0] Wgt_4_311;input [WEIGHT_SIZE-1:0] Wgt_4_312;input [WEIGHT_SIZE-1:0] Wgt_4_313;input [WEIGHT_SIZE-1:0] Wgt_4_314;input [WEIGHT_SIZE-1:0] Wgt_4_315;input [WEIGHT_SIZE-1:0] Wgt_4_316;input [WEIGHT_SIZE-1:0] Wgt_4_317;input [WEIGHT_SIZE-1:0] Wgt_4_318;input [WEIGHT_SIZE-1:0] Wgt_4_319;input [WEIGHT_SIZE-1:0] Wgt_4_320;input [WEIGHT_SIZE-1:0] Wgt_4_321;input [WEIGHT_SIZE-1:0] Wgt_4_322;input [WEIGHT_SIZE-1:0] Wgt_4_323;input [WEIGHT_SIZE-1:0] Wgt_4_324;input [WEIGHT_SIZE-1:0] Wgt_4_325;input [WEIGHT_SIZE-1:0] Wgt_4_326;input [WEIGHT_SIZE-1:0] Wgt_4_327;input [WEIGHT_SIZE-1:0] Wgt_4_328;input [WEIGHT_SIZE-1:0] Wgt_4_329;input [WEIGHT_SIZE-1:0] Wgt_4_330;input [WEIGHT_SIZE-1:0] Wgt_4_331;input [WEIGHT_SIZE-1:0] Wgt_4_332;input [WEIGHT_SIZE-1:0] Wgt_4_333;input [WEIGHT_SIZE-1:0] Wgt_4_334;input [WEIGHT_SIZE-1:0] Wgt_4_335;input [WEIGHT_SIZE-1:0] Wgt_4_336;input [WEIGHT_SIZE-1:0] Wgt_4_337;input [WEIGHT_SIZE-1:0] Wgt_4_338;input [WEIGHT_SIZE-1:0] Wgt_4_339;input [WEIGHT_SIZE-1:0] Wgt_4_340;input [WEIGHT_SIZE-1:0] Wgt_4_341;input [WEIGHT_SIZE-1:0] Wgt_4_342;input [WEIGHT_SIZE-1:0] Wgt_4_343;input [WEIGHT_SIZE-1:0] Wgt_4_344;input [WEIGHT_SIZE-1:0] Wgt_4_345;input [WEIGHT_SIZE-1:0] Wgt_4_346;input [WEIGHT_SIZE-1:0] Wgt_4_347;input [WEIGHT_SIZE-1:0] Wgt_4_348;input [WEIGHT_SIZE-1:0] Wgt_4_349;input [WEIGHT_SIZE-1:0] Wgt_4_350;input [WEIGHT_SIZE-1:0] Wgt_4_351;input [WEIGHT_SIZE-1:0] Wgt_4_352;input [WEIGHT_SIZE-1:0] Wgt_4_353;input [WEIGHT_SIZE-1:0] Wgt_4_354;input [WEIGHT_SIZE-1:0] Wgt_4_355;input [WEIGHT_SIZE-1:0] Wgt_4_356;input [WEIGHT_SIZE-1:0] Wgt_4_357;input [WEIGHT_SIZE-1:0] Wgt_4_358;input [WEIGHT_SIZE-1:0] Wgt_4_359;input [WEIGHT_SIZE-1:0] Wgt_4_360;input [WEIGHT_SIZE-1:0] Wgt_4_361;input [WEIGHT_SIZE-1:0] Wgt_4_362;input [WEIGHT_SIZE-1:0] Wgt_4_363;input [WEIGHT_SIZE-1:0] Wgt_4_364;input [WEIGHT_SIZE-1:0] Wgt_4_365;input [WEIGHT_SIZE-1:0] Wgt_4_366;input [WEIGHT_SIZE-1:0] Wgt_4_367;input [WEIGHT_SIZE-1:0] Wgt_4_368;input [WEIGHT_SIZE-1:0] Wgt_4_369;input [WEIGHT_SIZE-1:0] Wgt_4_370;input [WEIGHT_SIZE-1:0] Wgt_4_371;input [WEIGHT_SIZE-1:0] Wgt_4_372;input [WEIGHT_SIZE-1:0] Wgt_4_373;input [WEIGHT_SIZE-1:0] Wgt_4_374;input [WEIGHT_SIZE-1:0] Wgt_4_375;input [WEIGHT_SIZE-1:0] Wgt_4_376;input [WEIGHT_SIZE-1:0] Wgt_4_377;input [WEIGHT_SIZE-1:0] Wgt_4_378;input [WEIGHT_SIZE-1:0] Wgt_4_379;input [WEIGHT_SIZE-1:0] Wgt_4_380;input [WEIGHT_SIZE-1:0] Wgt_4_381;input [WEIGHT_SIZE-1:0] Wgt_4_382;input [WEIGHT_SIZE-1:0] Wgt_4_383;input [WEIGHT_SIZE-1:0] Wgt_4_384;input [WEIGHT_SIZE-1:0] Wgt_4_385;input [WEIGHT_SIZE-1:0] Wgt_4_386;input [WEIGHT_SIZE-1:0] Wgt_4_387;input [WEIGHT_SIZE-1:0] Wgt_4_388;input [WEIGHT_SIZE-1:0] Wgt_4_389;input [WEIGHT_SIZE-1:0] Wgt_4_390;input [WEIGHT_SIZE-1:0] Wgt_4_391;input [WEIGHT_SIZE-1:0] Wgt_4_392;input [WEIGHT_SIZE-1:0] Wgt_4_393;input [WEIGHT_SIZE-1:0] Wgt_4_394;input [WEIGHT_SIZE-1:0] Wgt_4_395;input [WEIGHT_SIZE-1:0] Wgt_4_396;input [WEIGHT_SIZE-1:0] Wgt_4_397;input [WEIGHT_SIZE-1:0] Wgt_4_398;input [WEIGHT_SIZE-1:0] Wgt_4_399;input [WEIGHT_SIZE-1:0] Wgt_4_400;input [WEIGHT_SIZE-1:0] Wgt_4_401;input [WEIGHT_SIZE-1:0] Wgt_4_402;input [WEIGHT_SIZE-1:0] Wgt_4_403;input [WEIGHT_SIZE-1:0] Wgt_4_404;input [WEIGHT_SIZE-1:0] Wgt_4_405;input [WEIGHT_SIZE-1:0] Wgt_4_406;input [WEIGHT_SIZE-1:0] Wgt_4_407;input [WEIGHT_SIZE-1:0] Wgt_4_408;input [WEIGHT_SIZE-1:0] Wgt_4_409;input [WEIGHT_SIZE-1:0] Wgt_4_410;input [WEIGHT_SIZE-1:0] Wgt_4_411;input [WEIGHT_SIZE-1:0] Wgt_4_412;input [WEIGHT_SIZE-1:0] Wgt_4_413;input [WEIGHT_SIZE-1:0] Wgt_4_414;input [WEIGHT_SIZE-1:0] Wgt_4_415;input [WEIGHT_SIZE-1:0] Wgt_4_416;input [WEIGHT_SIZE-1:0] Wgt_4_417;input [WEIGHT_SIZE-1:0] Wgt_4_418;input [WEIGHT_SIZE-1:0] Wgt_4_419;input [WEIGHT_SIZE-1:0] Wgt_4_420;input [WEIGHT_SIZE-1:0] Wgt_4_421;input [WEIGHT_SIZE-1:0] Wgt_4_422;input [WEIGHT_SIZE-1:0] Wgt_4_423;input [WEIGHT_SIZE-1:0] Wgt_4_424;input [WEIGHT_SIZE-1:0] Wgt_4_425;input [WEIGHT_SIZE-1:0] Wgt_4_426;input [WEIGHT_SIZE-1:0] Wgt_4_427;input [WEIGHT_SIZE-1:0] Wgt_4_428;input [WEIGHT_SIZE-1:0] Wgt_4_429;input [WEIGHT_SIZE-1:0] Wgt_4_430;input [WEIGHT_SIZE-1:0] Wgt_4_431;input [WEIGHT_SIZE-1:0] Wgt_4_432;input [WEIGHT_SIZE-1:0] Wgt_4_433;input [WEIGHT_SIZE-1:0] Wgt_4_434;input [WEIGHT_SIZE-1:0] Wgt_4_435;input [WEIGHT_SIZE-1:0] Wgt_4_436;input [WEIGHT_SIZE-1:0] Wgt_4_437;input [WEIGHT_SIZE-1:0] Wgt_4_438;input [WEIGHT_SIZE-1:0] Wgt_4_439;input [WEIGHT_SIZE-1:0] Wgt_4_440;input [WEIGHT_SIZE-1:0] Wgt_4_441;input [WEIGHT_SIZE-1:0] Wgt_4_442;input [WEIGHT_SIZE-1:0] Wgt_4_443;input [WEIGHT_SIZE-1:0] Wgt_4_444;input [WEIGHT_SIZE-1:0] Wgt_4_445;input [WEIGHT_SIZE-1:0] Wgt_4_446;input [WEIGHT_SIZE-1:0] Wgt_4_447;input [WEIGHT_SIZE-1:0] Wgt_4_448;input [WEIGHT_SIZE-1:0] Wgt_4_449;input [WEIGHT_SIZE-1:0] Wgt_4_450;input [WEIGHT_SIZE-1:0] Wgt_4_451;input [WEIGHT_SIZE-1:0] Wgt_4_452;input [WEIGHT_SIZE-1:0] Wgt_4_453;input [WEIGHT_SIZE-1:0] Wgt_4_454;input [WEIGHT_SIZE-1:0] Wgt_4_455;input [WEIGHT_SIZE-1:0] Wgt_4_456;input [WEIGHT_SIZE-1:0] Wgt_4_457;input [WEIGHT_SIZE-1:0] Wgt_4_458;input [WEIGHT_SIZE-1:0] Wgt_4_459;input [WEIGHT_SIZE-1:0] Wgt_4_460;input [WEIGHT_SIZE-1:0] Wgt_4_461;input [WEIGHT_SIZE-1:0] Wgt_4_462;input [WEIGHT_SIZE-1:0] Wgt_4_463;input [WEIGHT_SIZE-1:0] Wgt_4_464;input [WEIGHT_SIZE-1:0] Wgt_4_465;input [WEIGHT_SIZE-1:0] Wgt_4_466;input [WEIGHT_SIZE-1:0] Wgt_4_467;input [WEIGHT_SIZE-1:0] Wgt_4_468;input [WEIGHT_SIZE-1:0] Wgt_4_469;input [WEIGHT_SIZE-1:0] Wgt_4_470;input [WEIGHT_SIZE-1:0] Wgt_4_471;input [WEIGHT_SIZE-1:0] Wgt_4_472;input [WEIGHT_SIZE-1:0] Wgt_4_473;input [WEIGHT_SIZE-1:0] Wgt_4_474;input [WEIGHT_SIZE-1:0] Wgt_4_475;input [WEIGHT_SIZE-1:0] Wgt_4_476;input [WEIGHT_SIZE-1:0] Wgt_4_477;input [WEIGHT_SIZE-1:0] Wgt_4_478;input [WEIGHT_SIZE-1:0] Wgt_4_479;input [WEIGHT_SIZE-1:0] Wgt_4_480;input [WEIGHT_SIZE-1:0] Wgt_4_481;input [WEIGHT_SIZE-1:0] Wgt_4_482;input [WEIGHT_SIZE-1:0] Wgt_4_483;input [WEIGHT_SIZE-1:0] Wgt_4_484;input [WEIGHT_SIZE-1:0] Wgt_4_485;input [WEIGHT_SIZE-1:0] Wgt_4_486;input [WEIGHT_SIZE-1:0] Wgt_4_487;input [WEIGHT_SIZE-1:0] Wgt_4_488;input [WEIGHT_SIZE-1:0] Wgt_4_489;input [WEIGHT_SIZE-1:0] Wgt_4_490;input [WEIGHT_SIZE-1:0] Wgt_4_491;input [WEIGHT_SIZE-1:0] Wgt_4_492;input [WEIGHT_SIZE-1:0] Wgt_4_493;input [WEIGHT_SIZE-1:0] Wgt_4_494;input [WEIGHT_SIZE-1:0] Wgt_4_495;input [WEIGHT_SIZE-1:0] Wgt_4_496;input [WEIGHT_SIZE-1:0] Wgt_4_497;input [WEIGHT_SIZE-1:0] Wgt_4_498;input [WEIGHT_SIZE-1:0] Wgt_4_499;input [WEIGHT_SIZE-1:0] Wgt_4_500;input [WEIGHT_SIZE-1:0] Wgt_4_501;input [WEIGHT_SIZE-1:0] Wgt_4_502;input [WEIGHT_SIZE-1:0] Wgt_4_503;input [WEIGHT_SIZE-1:0] Wgt_4_504;input [WEIGHT_SIZE-1:0] Wgt_4_505;input [WEIGHT_SIZE-1:0] Wgt_4_506;input [WEIGHT_SIZE-1:0] Wgt_4_507;input [WEIGHT_SIZE-1:0] Wgt_4_508;input [WEIGHT_SIZE-1:0] Wgt_4_509;input [WEIGHT_SIZE-1:0] Wgt_4_510;input [WEIGHT_SIZE-1:0] Wgt_4_511;input [WEIGHT_SIZE-1:0] Wgt_4_512;input [WEIGHT_SIZE-1:0] Wgt_4_513;input [WEIGHT_SIZE-1:0] Wgt_4_514;input [WEIGHT_SIZE-1:0] Wgt_4_515;input [WEIGHT_SIZE-1:0] Wgt_4_516;input [WEIGHT_SIZE-1:0] Wgt_4_517;input [WEIGHT_SIZE-1:0] Wgt_4_518;input [WEIGHT_SIZE-1:0] Wgt_4_519;input [WEIGHT_SIZE-1:0] Wgt_4_520;input [WEIGHT_SIZE-1:0] Wgt_4_521;input [WEIGHT_SIZE-1:0] Wgt_4_522;input [WEIGHT_SIZE-1:0] Wgt_4_523;input [WEIGHT_SIZE-1:0] Wgt_4_524;input [WEIGHT_SIZE-1:0] Wgt_4_525;input [WEIGHT_SIZE-1:0] Wgt_4_526;input [WEIGHT_SIZE-1:0] Wgt_4_527;input [WEIGHT_SIZE-1:0] Wgt_4_528;input [WEIGHT_SIZE-1:0] Wgt_4_529;input [WEIGHT_SIZE-1:0] Wgt_4_530;input [WEIGHT_SIZE-1:0] Wgt_4_531;input [WEIGHT_SIZE-1:0] Wgt_4_532;input [WEIGHT_SIZE-1:0] Wgt_4_533;input [WEIGHT_SIZE-1:0] Wgt_4_534;input [WEIGHT_SIZE-1:0] Wgt_4_535;input [WEIGHT_SIZE-1:0] Wgt_4_536;input [WEIGHT_SIZE-1:0] Wgt_4_537;input [WEIGHT_SIZE-1:0] Wgt_4_538;input [WEIGHT_SIZE-1:0] Wgt_4_539;input [WEIGHT_SIZE-1:0] Wgt_4_540;input [WEIGHT_SIZE-1:0] Wgt_4_541;input [WEIGHT_SIZE-1:0] Wgt_4_542;input [WEIGHT_SIZE-1:0] Wgt_4_543;input [WEIGHT_SIZE-1:0] Wgt_4_544;input [WEIGHT_SIZE-1:0] Wgt_4_545;input [WEIGHT_SIZE-1:0] Wgt_4_546;input [WEIGHT_SIZE-1:0] Wgt_4_547;input [WEIGHT_SIZE-1:0] Wgt_4_548;input [WEIGHT_SIZE-1:0] Wgt_4_549;input [WEIGHT_SIZE-1:0] Wgt_4_550;input [WEIGHT_SIZE-1:0] Wgt_4_551;input [WEIGHT_SIZE-1:0] Wgt_4_552;input [WEIGHT_SIZE-1:0] Wgt_4_553;input [WEIGHT_SIZE-1:0] Wgt_4_554;input [WEIGHT_SIZE-1:0] Wgt_4_555;input [WEIGHT_SIZE-1:0] Wgt_4_556;input [WEIGHT_SIZE-1:0] Wgt_4_557;input [WEIGHT_SIZE-1:0] Wgt_4_558;input [WEIGHT_SIZE-1:0] Wgt_4_559;input [WEIGHT_SIZE-1:0] Wgt_4_560;input [WEIGHT_SIZE-1:0] Wgt_4_561;input [WEIGHT_SIZE-1:0] Wgt_4_562;input [WEIGHT_SIZE-1:0] Wgt_4_563;input [WEIGHT_SIZE-1:0] Wgt_4_564;input [WEIGHT_SIZE-1:0] Wgt_4_565;input [WEIGHT_SIZE-1:0] Wgt_4_566;input [WEIGHT_SIZE-1:0] Wgt_4_567;input [WEIGHT_SIZE-1:0] Wgt_4_568;input [WEIGHT_SIZE-1:0] Wgt_4_569;input [WEIGHT_SIZE-1:0] Wgt_4_570;input [WEIGHT_SIZE-1:0] Wgt_4_571;input [WEIGHT_SIZE-1:0] Wgt_4_572;input [WEIGHT_SIZE-1:0] Wgt_4_573;input [WEIGHT_SIZE-1:0] Wgt_4_574;input [WEIGHT_SIZE-1:0] Wgt_4_575;input [WEIGHT_SIZE-1:0] Wgt_4_576;input [WEIGHT_SIZE-1:0] Wgt_4_577;input [WEIGHT_SIZE-1:0] Wgt_4_578;input [WEIGHT_SIZE-1:0] Wgt_4_579;input [WEIGHT_SIZE-1:0] Wgt_4_580;input [WEIGHT_SIZE-1:0] Wgt_4_581;input [WEIGHT_SIZE-1:0] Wgt_4_582;input [WEIGHT_SIZE-1:0] Wgt_4_583;input [WEIGHT_SIZE-1:0] Wgt_4_584;input [WEIGHT_SIZE-1:0] Wgt_4_585;input [WEIGHT_SIZE-1:0] Wgt_4_586;input [WEIGHT_SIZE-1:0] Wgt_4_587;input [WEIGHT_SIZE-1:0] Wgt_4_588;input [WEIGHT_SIZE-1:0] Wgt_4_589;input [WEIGHT_SIZE-1:0] Wgt_4_590;input [WEIGHT_SIZE-1:0] Wgt_4_591;input [WEIGHT_SIZE-1:0] Wgt_4_592;input [WEIGHT_SIZE-1:0] Wgt_4_593;input [WEIGHT_SIZE-1:0] Wgt_4_594;input [WEIGHT_SIZE-1:0] Wgt_4_595;input [WEIGHT_SIZE-1:0] Wgt_4_596;input [WEIGHT_SIZE-1:0] Wgt_4_597;input [WEIGHT_SIZE-1:0] Wgt_4_598;input [WEIGHT_SIZE-1:0] Wgt_4_599;input [WEIGHT_SIZE-1:0] Wgt_4_600;input [WEIGHT_SIZE-1:0] Wgt_4_601;input [WEIGHT_SIZE-1:0] Wgt_4_602;input [WEIGHT_SIZE-1:0] Wgt_4_603;input [WEIGHT_SIZE-1:0] Wgt_4_604;input [WEIGHT_SIZE-1:0] Wgt_4_605;input [WEIGHT_SIZE-1:0] Wgt_4_606;input [WEIGHT_SIZE-1:0] Wgt_4_607;input [WEIGHT_SIZE-1:0] Wgt_4_608;input [WEIGHT_SIZE-1:0] Wgt_4_609;input [WEIGHT_SIZE-1:0] Wgt_4_610;input [WEIGHT_SIZE-1:0] Wgt_4_611;input [WEIGHT_SIZE-1:0] Wgt_4_612;input [WEIGHT_SIZE-1:0] Wgt_4_613;input [WEIGHT_SIZE-1:0] Wgt_4_614;input [WEIGHT_SIZE-1:0] Wgt_4_615;input [WEIGHT_SIZE-1:0] Wgt_4_616;input [WEIGHT_SIZE-1:0] Wgt_4_617;input [WEIGHT_SIZE-1:0] Wgt_4_618;input [WEIGHT_SIZE-1:0] Wgt_4_619;input [WEIGHT_SIZE-1:0] Wgt_4_620;input [WEIGHT_SIZE-1:0] Wgt_4_621;input [WEIGHT_SIZE-1:0] Wgt_4_622;input [WEIGHT_SIZE-1:0] Wgt_4_623;input [WEIGHT_SIZE-1:0] Wgt_4_624;input [WEIGHT_SIZE-1:0] Wgt_4_625;input [WEIGHT_SIZE-1:0] Wgt_4_626;input [WEIGHT_SIZE-1:0] Wgt_4_627;input [WEIGHT_SIZE-1:0] Wgt_4_628;input [WEIGHT_SIZE-1:0] Wgt_4_629;input [WEIGHT_SIZE-1:0] Wgt_4_630;input [WEIGHT_SIZE-1:0] Wgt_4_631;input [WEIGHT_SIZE-1:0] Wgt_4_632;input [WEIGHT_SIZE-1:0] Wgt_4_633;input [WEIGHT_SIZE-1:0] Wgt_4_634;input [WEIGHT_SIZE-1:0] Wgt_4_635;input [WEIGHT_SIZE-1:0] Wgt_4_636;input [WEIGHT_SIZE-1:0] Wgt_4_637;input [WEIGHT_SIZE-1:0] Wgt_4_638;input [WEIGHT_SIZE-1:0] Wgt_4_639;input [WEIGHT_SIZE-1:0] Wgt_4_640;input [WEIGHT_SIZE-1:0] Wgt_4_641;input [WEIGHT_SIZE-1:0] Wgt_4_642;input [WEIGHT_SIZE-1:0] Wgt_4_643;input [WEIGHT_SIZE-1:0] Wgt_4_644;input [WEIGHT_SIZE-1:0] Wgt_4_645;input [WEIGHT_SIZE-1:0] Wgt_4_646;input [WEIGHT_SIZE-1:0] Wgt_4_647;input [WEIGHT_SIZE-1:0] Wgt_4_648;input [WEIGHT_SIZE-1:0] Wgt_4_649;input [WEIGHT_SIZE-1:0] Wgt_4_650;input [WEIGHT_SIZE-1:0] Wgt_4_651;input [WEIGHT_SIZE-1:0] Wgt_4_652;input [WEIGHT_SIZE-1:0] Wgt_4_653;input [WEIGHT_SIZE-1:0] Wgt_4_654;input [WEIGHT_SIZE-1:0] Wgt_4_655;input [WEIGHT_SIZE-1:0] Wgt_4_656;input [WEIGHT_SIZE-1:0] Wgt_4_657;input [WEIGHT_SIZE-1:0] Wgt_4_658;input [WEIGHT_SIZE-1:0] Wgt_4_659;input [WEIGHT_SIZE-1:0] Wgt_4_660;input [WEIGHT_SIZE-1:0] Wgt_4_661;input [WEIGHT_SIZE-1:0] Wgt_4_662;input [WEIGHT_SIZE-1:0] Wgt_4_663;input [WEIGHT_SIZE-1:0] Wgt_4_664;input [WEIGHT_SIZE-1:0] Wgt_4_665;input [WEIGHT_SIZE-1:0] Wgt_4_666;input [WEIGHT_SIZE-1:0] Wgt_4_667;input [WEIGHT_SIZE-1:0] Wgt_4_668;input [WEIGHT_SIZE-1:0] Wgt_4_669;input [WEIGHT_SIZE-1:0] Wgt_4_670;input [WEIGHT_SIZE-1:0] Wgt_4_671;input [WEIGHT_SIZE-1:0] Wgt_4_672;input [WEIGHT_SIZE-1:0] Wgt_4_673;input [WEIGHT_SIZE-1:0] Wgt_4_674;input [WEIGHT_SIZE-1:0] Wgt_4_675;input [WEIGHT_SIZE-1:0] Wgt_4_676;input [WEIGHT_SIZE-1:0] Wgt_4_677;input [WEIGHT_SIZE-1:0] Wgt_4_678;input [WEIGHT_SIZE-1:0] Wgt_4_679;input [WEIGHT_SIZE-1:0] Wgt_4_680;input [WEIGHT_SIZE-1:0] Wgt_4_681;input [WEIGHT_SIZE-1:0] Wgt_4_682;input [WEIGHT_SIZE-1:0] Wgt_4_683;input [WEIGHT_SIZE-1:0] Wgt_4_684;input [WEIGHT_SIZE-1:0] Wgt_4_685;input [WEIGHT_SIZE-1:0] Wgt_4_686;input [WEIGHT_SIZE-1:0] Wgt_4_687;input [WEIGHT_SIZE-1:0] Wgt_4_688;input [WEIGHT_SIZE-1:0] Wgt_4_689;input [WEIGHT_SIZE-1:0] Wgt_4_690;input [WEIGHT_SIZE-1:0] Wgt_4_691;input [WEIGHT_SIZE-1:0] Wgt_4_692;input [WEIGHT_SIZE-1:0] Wgt_4_693;input [WEIGHT_SIZE-1:0] Wgt_4_694;input [WEIGHT_SIZE-1:0] Wgt_4_695;input [WEIGHT_SIZE-1:0] Wgt_4_696;input [WEIGHT_SIZE-1:0] Wgt_4_697;input [WEIGHT_SIZE-1:0] Wgt_4_698;input [WEIGHT_SIZE-1:0] Wgt_4_699;input [WEIGHT_SIZE-1:0] Wgt_4_700;input [WEIGHT_SIZE-1:0] Wgt_4_701;input [WEIGHT_SIZE-1:0] Wgt_4_702;input [WEIGHT_SIZE-1:0] Wgt_4_703;input [WEIGHT_SIZE-1:0] Wgt_4_704;input [WEIGHT_SIZE-1:0] Wgt_4_705;input [WEIGHT_SIZE-1:0] Wgt_4_706;input [WEIGHT_SIZE-1:0] Wgt_4_707;input [WEIGHT_SIZE-1:0] Wgt_4_708;input [WEIGHT_SIZE-1:0] Wgt_4_709;input [WEIGHT_SIZE-1:0] Wgt_4_710;input [WEIGHT_SIZE-1:0] Wgt_4_711;input [WEIGHT_SIZE-1:0] Wgt_4_712;input [WEIGHT_SIZE-1:0] Wgt_4_713;input [WEIGHT_SIZE-1:0] Wgt_4_714;input [WEIGHT_SIZE-1:0] Wgt_4_715;input [WEIGHT_SIZE-1:0] Wgt_4_716;input [WEIGHT_SIZE-1:0] Wgt_4_717;input [WEIGHT_SIZE-1:0] Wgt_4_718;input [WEIGHT_SIZE-1:0] Wgt_4_719;input [WEIGHT_SIZE-1:0] Wgt_4_720;input [WEIGHT_SIZE-1:0] Wgt_4_721;input [WEIGHT_SIZE-1:0] Wgt_4_722;input [WEIGHT_SIZE-1:0] Wgt_4_723;input [WEIGHT_SIZE-1:0] Wgt_4_724;input [WEIGHT_SIZE-1:0] Wgt_4_725;input [WEIGHT_SIZE-1:0] Wgt_4_726;input [WEIGHT_SIZE-1:0] Wgt_4_727;input [WEIGHT_SIZE-1:0] Wgt_4_728;input [WEIGHT_SIZE-1:0] Wgt_4_729;input [WEIGHT_SIZE-1:0] Wgt_4_730;input [WEIGHT_SIZE-1:0] Wgt_4_731;input [WEIGHT_SIZE-1:0] Wgt_4_732;input [WEIGHT_SIZE-1:0] Wgt_4_733;input [WEIGHT_SIZE-1:0] Wgt_4_734;input [WEIGHT_SIZE-1:0] Wgt_4_735;input [WEIGHT_SIZE-1:0] Wgt_4_736;input [WEIGHT_SIZE-1:0] Wgt_4_737;input [WEIGHT_SIZE-1:0] Wgt_4_738;input [WEIGHT_SIZE-1:0] Wgt_4_739;input [WEIGHT_SIZE-1:0] Wgt_4_740;input [WEIGHT_SIZE-1:0] Wgt_4_741;input [WEIGHT_SIZE-1:0] Wgt_4_742;input [WEIGHT_SIZE-1:0] Wgt_4_743;input [WEIGHT_SIZE-1:0] Wgt_4_744;input [WEIGHT_SIZE-1:0] Wgt_4_745;input [WEIGHT_SIZE-1:0] Wgt_4_746;input [WEIGHT_SIZE-1:0] Wgt_4_747;input [WEIGHT_SIZE-1:0] Wgt_4_748;input [WEIGHT_SIZE-1:0] Wgt_4_749;input [WEIGHT_SIZE-1:0] Wgt_4_750;input [WEIGHT_SIZE-1:0] Wgt_4_751;input [WEIGHT_SIZE-1:0] Wgt_4_752;input [WEIGHT_SIZE-1:0] Wgt_4_753;input [WEIGHT_SIZE-1:0] Wgt_4_754;input [WEIGHT_SIZE-1:0] Wgt_4_755;input [WEIGHT_SIZE-1:0] Wgt_4_756;input [WEIGHT_SIZE-1:0] Wgt_4_757;input [WEIGHT_SIZE-1:0] Wgt_4_758;input [WEIGHT_SIZE-1:0] Wgt_4_759;input [WEIGHT_SIZE-1:0] Wgt_4_760;input [WEIGHT_SIZE-1:0] Wgt_4_761;input [WEIGHT_SIZE-1:0] Wgt_4_762;input [WEIGHT_SIZE-1:0] Wgt_4_763;input [WEIGHT_SIZE-1:0] Wgt_4_764;input [WEIGHT_SIZE-1:0] Wgt_4_765;input [WEIGHT_SIZE-1:0] Wgt_4_766;input [WEIGHT_SIZE-1:0] Wgt_4_767;input [WEIGHT_SIZE-1:0] Wgt_4_768;input [WEIGHT_SIZE-1:0] Wgt_4_769;input [WEIGHT_SIZE-1:0] Wgt_4_770;input [WEIGHT_SIZE-1:0] Wgt_4_771;input [WEIGHT_SIZE-1:0] Wgt_4_772;input [WEIGHT_SIZE-1:0] Wgt_4_773;input [WEIGHT_SIZE-1:0] Wgt_4_774;input [WEIGHT_SIZE-1:0] Wgt_4_775;input [WEIGHT_SIZE-1:0] Wgt_4_776;input [WEIGHT_SIZE-1:0] Wgt_4_777;input [WEIGHT_SIZE-1:0] Wgt_4_778;input [WEIGHT_SIZE-1:0] Wgt_4_779;input [WEIGHT_SIZE-1:0] Wgt_4_780;input [WEIGHT_SIZE-1:0] Wgt_4_781;input [WEIGHT_SIZE-1:0] Wgt_4_782;input [WEIGHT_SIZE-1:0] Wgt_4_783;input [WEIGHT_SIZE-1:0] Wgt_4_784;input [WEIGHT_SIZE-1:0] Wgt_5_0;input [WEIGHT_SIZE-1:0] Wgt_5_1;input [WEIGHT_SIZE-1:0] Wgt_5_2;input [WEIGHT_SIZE-1:0] Wgt_5_3;input [WEIGHT_SIZE-1:0] Wgt_5_4;input [WEIGHT_SIZE-1:0] Wgt_5_5;input [WEIGHT_SIZE-1:0] Wgt_5_6;input [WEIGHT_SIZE-1:0] Wgt_5_7;input [WEIGHT_SIZE-1:0] Wgt_5_8;input [WEIGHT_SIZE-1:0] Wgt_5_9;input [WEIGHT_SIZE-1:0] Wgt_5_10;input [WEIGHT_SIZE-1:0] Wgt_5_11;input [WEIGHT_SIZE-1:0] Wgt_5_12;input [WEIGHT_SIZE-1:0] Wgt_5_13;input [WEIGHT_SIZE-1:0] Wgt_5_14;input [WEIGHT_SIZE-1:0] Wgt_5_15;input [WEIGHT_SIZE-1:0] Wgt_5_16;input [WEIGHT_SIZE-1:0] Wgt_5_17;input [WEIGHT_SIZE-1:0] Wgt_5_18;input [WEIGHT_SIZE-1:0] Wgt_5_19;input [WEIGHT_SIZE-1:0] Wgt_5_20;input [WEIGHT_SIZE-1:0] Wgt_5_21;input [WEIGHT_SIZE-1:0] Wgt_5_22;input [WEIGHT_SIZE-1:0] Wgt_5_23;input [WEIGHT_SIZE-1:0] Wgt_5_24;input [WEIGHT_SIZE-1:0] Wgt_5_25;input [WEIGHT_SIZE-1:0] Wgt_5_26;input [WEIGHT_SIZE-1:0] Wgt_5_27;input [WEIGHT_SIZE-1:0] Wgt_5_28;input [WEIGHT_SIZE-1:0] Wgt_5_29;input [WEIGHT_SIZE-1:0] Wgt_5_30;input [WEIGHT_SIZE-1:0] Wgt_5_31;input [WEIGHT_SIZE-1:0] Wgt_5_32;input [WEIGHT_SIZE-1:0] Wgt_5_33;input [WEIGHT_SIZE-1:0] Wgt_5_34;input [WEIGHT_SIZE-1:0] Wgt_5_35;input [WEIGHT_SIZE-1:0] Wgt_5_36;input [WEIGHT_SIZE-1:0] Wgt_5_37;input [WEIGHT_SIZE-1:0] Wgt_5_38;input [WEIGHT_SIZE-1:0] Wgt_5_39;input [WEIGHT_SIZE-1:0] Wgt_5_40;input [WEIGHT_SIZE-1:0] Wgt_5_41;input [WEIGHT_SIZE-1:0] Wgt_5_42;input [WEIGHT_SIZE-1:0] Wgt_5_43;input [WEIGHT_SIZE-1:0] Wgt_5_44;input [WEIGHT_SIZE-1:0] Wgt_5_45;input [WEIGHT_SIZE-1:0] Wgt_5_46;input [WEIGHT_SIZE-1:0] Wgt_5_47;input [WEIGHT_SIZE-1:0] Wgt_5_48;input [WEIGHT_SIZE-1:0] Wgt_5_49;input [WEIGHT_SIZE-1:0] Wgt_5_50;input [WEIGHT_SIZE-1:0] Wgt_5_51;input [WEIGHT_SIZE-1:0] Wgt_5_52;input [WEIGHT_SIZE-1:0] Wgt_5_53;input [WEIGHT_SIZE-1:0] Wgt_5_54;input [WEIGHT_SIZE-1:0] Wgt_5_55;input [WEIGHT_SIZE-1:0] Wgt_5_56;input [WEIGHT_SIZE-1:0] Wgt_5_57;input [WEIGHT_SIZE-1:0] Wgt_5_58;input [WEIGHT_SIZE-1:0] Wgt_5_59;input [WEIGHT_SIZE-1:0] Wgt_5_60;input [WEIGHT_SIZE-1:0] Wgt_5_61;input [WEIGHT_SIZE-1:0] Wgt_5_62;input [WEIGHT_SIZE-1:0] Wgt_5_63;input [WEIGHT_SIZE-1:0] Wgt_5_64;input [WEIGHT_SIZE-1:0] Wgt_5_65;input [WEIGHT_SIZE-1:0] Wgt_5_66;input [WEIGHT_SIZE-1:0] Wgt_5_67;input [WEIGHT_SIZE-1:0] Wgt_5_68;input [WEIGHT_SIZE-1:0] Wgt_5_69;input [WEIGHT_SIZE-1:0] Wgt_5_70;input [WEIGHT_SIZE-1:0] Wgt_5_71;input [WEIGHT_SIZE-1:0] Wgt_5_72;input [WEIGHT_SIZE-1:0] Wgt_5_73;input [WEIGHT_SIZE-1:0] Wgt_5_74;input [WEIGHT_SIZE-1:0] Wgt_5_75;input [WEIGHT_SIZE-1:0] Wgt_5_76;input [WEIGHT_SIZE-1:0] Wgt_5_77;input [WEIGHT_SIZE-1:0] Wgt_5_78;input [WEIGHT_SIZE-1:0] Wgt_5_79;input [WEIGHT_SIZE-1:0] Wgt_5_80;input [WEIGHT_SIZE-1:0] Wgt_5_81;input [WEIGHT_SIZE-1:0] Wgt_5_82;input [WEIGHT_SIZE-1:0] Wgt_5_83;input [WEIGHT_SIZE-1:0] Wgt_5_84;input [WEIGHT_SIZE-1:0] Wgt_5_85;input [WEIGHT_SIZE-1:0] Wgt_5_86;input [WEIGHT_SIZE-1:0] Wgt_5_87;input [WEIGHT_SIZE-1:0] Wgt_5_88;input [WEIGHT_SIZE-1:0] Wgt_5_89;input [WEIGHT_SIZE-1:0] Wgt_5_90;input [WEIGHT_SIZE-1:0] Wgt_5_91;input [WEIGHT_SIZE-1:0] Wgt_5_92;input [WEIGHT_SIZE-1:0] Wgt_5_93;input [WEIGHT_SIZE-1:0] Wgt_5_94;input [WEIGHT_SIZE-1:0] Wgt_5_95;input [WEIGHT_SIZE-1:0] Wgt_5_96;input [WEIGHT_SIZE-1:0] Wgt_5_97;input [WEIGHT_SIZE-1:0] Wgt_5_98;input [WEIGHT_SIZE-1:0] Wgt_5_99;input [WEIGHT_SIZE-1:0] Wgt_5_100;input [WEIGHT_SIZE-1:0] Wgt_5_101;input [WEIGHT_SIZE-1:0] Wgt_5_102;input [WEIGHT_SIZE-1:0] Wgt_5_103;input [WEIGHT_SIZE-1:0] Wgt_5_104;input [WEIGHT_SIZE-1:0] Wgt_5_105;input [WEIGHT_SIZE-1:0] Wgt_5_106;input [WEIGHT_SIZE-1:0] Wgt_5_107;input [WEIGHT_SIZE-1:0] Wgt_5_108;input [WEIGHT_SIZE-1:0] Wgt_5_109;input [WEIGHT_SIZE-1:0] Wgt_5_110;input [WEIGHT_SIZE-1:0] Wgt_5_111;input [WEIGHT_SIZE-1:0] Wgt_5_112;input [WEIGHT_SIZE-1:0] Wgt_5_113;input [WEIGHT_SIZE-1:0] Wgt_5_114;input [WEIGHT_SIZE-1:0] Wgt_5_115;input [WEIGHT_SIZE-1:0] Wgt_5_116;input [WEIGHT_SIZE-1:0] Wgt_5_117;input [WEIGHT_SIZE-1:0] Wgt_5_118;input [WEIGHT_SIZE-1:0] Wgt_5_119;input [WEIGHT_SIZE-1:0] Wgt_5_120;input [WEIGHT_SIZE-1:0] Wgt_5_121;input [WEIGHT_SIZE-1:0] Wgt_5_122;input [WEIGHT_SIZE-1:0] Wgt_5_123;input [WEIGHT_SIZE-1:0] Wgt_5_124;input [WEIGHT_SIZE-1:0] Wgt_5_125;input [WEIGHT_SIZE-1:0] Wgt_5_126;input [WEIGHT_SIZE-1:0] Wgt_5_127;input [WEIGHT_SIZE-1:0] Wgt_5_128;input [WEIGHT_SIZE-1:0] Wgt_5_129;input [WEIGHT_SIZE-1:0] Wgt_5_130;input [WEIGHT_SIZE-1:0] Wgt_5_131;input [WEIGHT_SIZE-1:0] Wgt_5_132;input [WEIGHT_SIZE-1:0] Wgt_5_133;input [WEIGHT_SIZE-1:0] Wgt_5_134;input [WEIGHT_SIZE-1:0] Wgt_5_135;input [WEIGHT_SIZE-1:0] Wgt_5_136;input [WEIGHT_SIZE-1:0] Wgt_5_137;input [WEIGHT_SIZE-1:0] Wgt_5_138;input [WEIGHT_SIZE-1:0] Wgt_5_139;input [WEIGHT_SIZE-1:0] Wgt_5_140;input [WEIGHT_SIZE-1:0] Wgt_5_141;input [WEIGHT_SIZE-1:0] Wgt_5_142;input [WEIGHT_SIZE-1:0] Wgt_5_143;input [WEIGHT_SIZE-1:0] Wgt_5_144;input [WEIGHT_SIZE-1:0] Wgt_5_145;input [WEIGHT_SIZE-1:0] Wgt_5_146;input [WEIGHT_SIZE-1:0] Wgt_5_147;input [WEIGHT_SIZE-1:0] Wgt_5_148;input [WEIGHT_SIZE-1:0] Wgt_5_149;input [WEIGHT_SIZE-1:0] Wgt_5_150;input [WEIGHT_SIZE-1:0] Wgt_5_151;input [WEIGHT_SIZE-1:0] Wgt_5_152;input [WEIGHT_SIZE-1:0] Wgt_5_153;input [WEIGHT_SIZE-1:0] Wgt_5_154;input [WEIGHT_SIZE-1:0] Wgt_5_155;input [WEIGHT_SIZE-1:0] Wgt_5_156;input [WEIGHT_SIZE-1:0] Wgt_5_157;input [WEIGHT_SIZE-1:0] Wgt_5_158;input [WEIGHT_SIZE-1:0] Wgt_5_159;input [WEIGHT_SIZE-1:0] Wgt_5_160;input [WEIGHT_SIZE-1:0] Wgt_5_161;input [WEIGHT_SIZE-1:0] Wgt_5_162;input [WEIGHT_SIZE-1:0] Wgt_5_163;input [WEIGHT_SIZE-1:0] Wgt_5_164;input [WEIGHT_SIZE-1:0] Wgt_5_165;input [WEIGHT_SIZE-1:0] Wgt_5_166;input [WEIGHT_SIZE-1:0] Wgt_5_167;input [WEIGHT_SIZE-1:0] Wgt_5_168;input [WEIGHT_SIZE-1:0] Wgt_5_169;input [WEIGHT_SIZE-1:0] Wgt_5_170;input [WEIGHT_SIZE-1:0] Wgt_5_171;input [WEIGHT_SIZE-1:0] Wgt_5_172;input [WEIGHT_SIZE-1:0] Wgt_5_173;input [WEIGHT_SIZE-1:0] Wgt_5_174;input [WEIGHT_SIZE-1:0] Wgt_5_175;input [WEIGHT_SIZE-1:0] Wgt_5_176;input [WEIGHT_SIZE-1:0] Wgt_5_177;input [WEIGHT_SIZE-1:0] Wgt_5_178;input [WEIGHT_SIZE-1:0] Wgt_5_179;input [WEIGHT_SIZE-1:0] Wgt_5_180;input [WEIGHT_SIZE-1:0] Wgt_5_181;input [WEIGHT_SIZE-1:0] Wgt_5_182;input [WEIGHT_SIZE-1:0] Wgt_5_183;input [WEIGHT_SIZE-1:0] Wgt_5_184;input [WEIGHT_SIZE-1:0] Wgt_5_185;input [WEIGHT_SIZE-1:0] Wgt_5_186;input [WEIGHT_SIZE-1:0] Wgt_5_187;input [WEIGHT_SIZE-1:0] Wgt_5_188;input [WEIGHT_SIZE-1:0] Wgt_5_189;input [WEIGHT_SIZE-1:0] Wgt_5_190;input [WEIGHT_SIZE-1:0] Wgt_5_191;input [WEIGHT_SIZE-1:0] Wgt_5_192;input [WEIGHT_SIZE-1:0] Wgt_5_193;input [WEIGHT_SIZE-1:0] Wgt_5_194;input [WEIGHT_SIZE-1:0] Wgt_5_195;input [WEIGHT_SIZE-1:0] Wgt_5_196;input [WEIGHT_SIZE-1:0] Wgt_5_197;input [WEIGHT_SIZE-1:0] Wgt_5_198;input [WEIGHT_SIZE-1:0] Wgt_5_199;input [WEIGHT_SIZE-1:0] Wgt_5_200;input [WEIGHT_SIZE-1:0] Wgt_5_201;input [WEIGHT_SIZE-1:0] Wgt_5_202;input [WEIGHT_SIZE-1:0] Wgt_5_203;input [WEIGHT_SIZE-1:0] Wgt_5_204;input [WEIGHT_SIZE-1:0] Wgt_5_205;input [WEIGHT_SIZE-1:0] Wgt_5_206;input [WEIGHT_SIZE-1:0] Wgt_5_207;input [WEIGHT_SIZE-1:0] Wgt_5_208;input [WEIGHT_SIZE-1:0] Wgt_5_209;input [WEIGHT_SIZE-1:0] Wgt_5_210;input [WEIGHT_SIZE-1:0] Wgt_5_211;input [WEIGHT_SIZE-1:0] Wgt_5_212;input [WEIGHT_SIZE-1:0] Wgt_5_213;input [WEIGHT_SIZE-1:0] Wgt_5_214;input [WEIGHT_SIZE-1:0] Wgt_5_215;input [WEIGHT_SIZE-1:0] Wgt_5_216;input [WEIGHT_SIZE-1:0] Wgt_5_217;input [WEIGHT_SIZE-1:0] Wgt_5_218;input [WEIGHT_SIZE-1:0] Wgt_5_219;input [WEIGHT_SIZE-1:0] Wgt_5_220;input [WEIGHT_SIZE-1:0] Wgt_5_221;input [WEIGHT_SIZE-1:0] Wgt_5_222;input [WEIGHT_SIZE-1:0] Wgt_5_223;input [WEIGHT_SIZE-1:0] Wgt_5_224;input [WEIGHT_SIZE-1:0] Wgt_5_225;input [WEIGHT_SIZE-1:0] Wgt_5_226;input [WEIGHT_SIZE-1:0] Wgt_5_227;input [WEIGHT_SIZE-1:0] Wgt_5_228;input [WEIGHT_SIZE-1:0] Wgt_5_229;input [WEIGHT_SIZE-1:0] Wgt_5_230;input [WEIGHT_SIZE-1:0] Wgt_5_231;input [WEIGHT_SIZE-1:0] Wgt_5_232;input [WEIGHT_SIZE-1:0] Wgt_5_233;input [WEIGHT_SIZE-1:0] Wgt_5_234;input [WEIGHT_SIZE-1:0] Wgt_5_235;input [WEIGHT_SIZE-1:0] Wgt_5_236;input [WEIGHT_SIZE-1:0] Wgt_5_237;input [WEIGHT_SIZE-1:0] Wgt_5_238;input [WEIGHT_SIZE-1:0] Wgt_5_239;input [WEIGHT_SIZE-1:0] Wgt_5_240;input [WEIGHT_SIZE-1:0] Wgt_5_241;input [WEIGHT_SIZE-1:0] Wgt_5_242;input [WEIGHT_SIZE-1:0] Wgt_5_243;input [WEIGHT_SIZE-1:0] Wgt_5_244;input [WEIGHT_SIZE-1:0] Wgt_5_245;input [WEIGHT_SIZE-1:0] Wgt_5_246;input [WEIGHT_SIZE-1:0] Wgt_5_247;input [WEIGHT_SIZE-1:0] Wgt_5_248;input [WEIGHT_SIZE-1:0] Wgt_5_249;input [WEIGHT_SIZE-1:0] Wgt_5_250;input [WEIGHT_SIZE-1:0] Wgt_5_251;input [WEIGHT_SIZE-1:0] Wgt_5_252;input [WEIGHT_SIZE-1:0] Wgt_5_253;input [WEIGHT_SIZE-1:0] Wgt_5_254;input [WEIGHT_SIZE-1:0] Wgt_5_255;input [WEIGHT_SIZE-1:0] Wgt_5_256;input [WEIGHT_SIZE-1:0] Wgt_5_257;input [WEIGHT_SIZE-1:0] Wgt_5_258;input [WEIGHT_SIZE-1:0] Wgt_5_259;input [WEIGHT_SIZE-1:0] Wgt_5_260;input [WEIGHT_SIZE-1:0] Wgt_5_261;input [WEIGHT_SIZE-1:0] Wgt_5_262;input [WEIGHT_SIZE-1:0] Wgt_5_263;input [WEIGHT_SIZE-1:0] Wgt_5_264;input [WEIGHT_SIZE-1:0] Wgt_5_265;input [WEIGHT_SIZE-1:0] Wgt_5_266;input [WEIGHT_SIZE-1:0] Wgt_5_267;input [WEIGHT_SIZE-1:0] Wgt_5_268;input [WEIGHT_SIZE-1:0] Wgt_5_269;input [WEIGHT_SIZE-1:0] Wgt_5_270;input [WEIGHT_SIZE-1:0] Wgt_5_271;input [WEIGHT_SIZE-1:0] Wgt_5_272;input [WEIGHT_SIZE-1:0] Wgt_5_273;input [WEIGHT_SIZE-1:0] Wgt_5_274;input [WEIGHT_SIZE-1:0] Wgt_5_275;input [WEIGHT_SIZE-1:0] Wgt_5_276;input [WEIGHT_SIZE-1:0] Wgt_5_277;input [WEIGHT_SIZE-1:0] Wgt_5_278;input [WEIGHT_SIZE-1:0] Wgt_5_279;input [WEIGHT_SIZE-1:0] Wgt_5_280;input [WEIGHT_SIZE-1:0] Wgt_5_281;input [WEIGHT_SIZE-1:0] Wgt_5_282;input [WEIGHT_SIZE-1:0] Wgt_5_283;input [WEIGHT_SIZE-1:0] Wgt_5_284;input [WEIGHT_SIZE-1:0] Wgt_5_285;input [WEIGHT_SIZE-1:0] Wgt_5_286;input [WEIGHT_SIZE-1:0] Wgt_5_287;input [WEIGHT_SIZE-1:0] Wgt_5_288;input [WEIGHT_SIZE-1:0] Wgt_5_289;input [WEIGHT_SIZE-1:0] Wgt_5_290;input [WEIGHT_SIZE-1:0] Wgt_5_291;input [WEIGHT_SIZE-1:0] Wgt_5_292;input [WEIGHT_SIZE-1:0] Wgt_5_293;input [WEIGHT_SIZE-1:0] Wgt_5_294;input [WEIGHT_SIZE-1:0] Wgt_5_295;input [WEIGHT_SIZE-1:0] Wgt_5_296;input [WEIGHT_SIZE-1:0] Wgt_5_297;input [WEIGHT_SIZE-1:0] Wgt_5_298;input [WEIGHT_SIZE-1:0] Wgt_5_299;input [WEIGHT_SIZE-1:0] Wgt_5_300;input [WEIGHT_SIZE-1:0] Wgt_5_301;input [WEIGHT_SIZE-1:0] Wgt_5_302;input [WEIGHT_SIZE-1:0] Wgt_5_303;input [WEIGHT_SIZE-1:0] Wgt_5_304;input [WEIGHT_SIZE-1:0] Wgt_5_305;input [WEIGHT_SIZE-1:0] Wgt_5_306;input [WEIGHT_SIZE-1:0] Wgt_5_307;input [WEIGHT_SIZE-1:0] Wgt_5_308;input [WEIGHT_SIZE-1:0] Wgt_5_309;input [WEIGHT_SIZE-1:0] Wgt_5_310;input [WEIGHT_SIZE-1:0] Wgt_5_311;input [WEIGHT_SIZE-1:0] Wgt_5_312;input [WEIGHT_SIZE-1:0] Wgt_5_313;input [WEIGHT_SIZE-1:0] Wgt_5_314;input [WEIGHT_SIZE-1:0] Wgt_5_315;input [WEIGHT_SIZE-1:0] Wgt_5_316;input [WEIGHT_SIZE-1:0] Wgt_5_317;input [WEIGHT_SIZE-1:0] Wgt_5_318;input [WEIGHT_SIZE-1:0] Wgt_5_319;input [WEIGHT_SIZE-1:0] Wgt_5_320;input [WEIGHT_SIZE-1:0] Wgt_5_321;input [WEIGHT_SIZE-1:0] Wgt_5_322;input [WEIGHT_SIZE-1:0] Wgt_5_323;input [WEIGHT_SIZE-1:0] Wgt_5_324;input [WEIGHT_SIZE-1:0] Wgt_5_325;input [WEIGHT_SIZE-1:0] Wgt_5_326;input [WEIGHT_SIZE-1:0] Wgt_5_327;input [WEIGHT_SIZE-1:0] Wgt_5_328;input [WEIGHT_SIZE-1:0] Wgt_5_329;input [WEIGHT_SIZE-1:0] Wgt_5_330;input [WEIGHT_SIZE-1:0] Wgt_5_331;input [WEIGHT_SIZE-1:0] Wgt_5_332;input [WEIGHT_SIZE-1:0] Wgt_5_333;input [WEIGHT_SIZE-1:0] Wgt_5_334;input [WEIGHT_SIZE-1:0] Wgt_5_335;input [WEIGHT_SIZE-1:0] Wgt_5_336;input [WEIGHT_SIZE-1:0] Wgt_5_337;input [WEIGHT_SIZE-1:0] Wgt_5_338;input [WEIGHT_SIZE-1:0] Wgt_5_339;input [WEIGHT_SIZE-1:0] Wgt_5_340;input [WEIGHT_SIZE-1:0] Wgt_5_341;input [WEIGHT_SIZE-1:0] Wgt_5_342;input [WEIGHT_SIZE-1:0] Wgt_5_343;input [WEIGHT_SIZE-1:0] Wgt_5_344;input [WEIGHT_SIZE-1:0] Wgt_5_345;input [WEIGHT_SIZE-1:0] Wgt_5_346;input [WEIGHT_SIZE-1:0] Wgt_5_347;input [WEIGHT_SIZE-1:0] Wgt_5_348;input [WEIGHT_SIZE-1:0] Wgt_5_349;input [WEIGHT_SIZE-1:0] Wgt_5_350;input [WEIGHT_SIZE-1:0] Wgt_5_351;input [WEIGHT_SIZE-1:0] Wgt_5_352;input [WEIGHT_SIZE-1:0] Wgt_5_353;input [WEIGHT_SIZE-1:0] Wgt_5_354;input [WEIGHT_SIZE-1:0] Wgt_5_355;input [WEIGHT_SIZE-1:0] Wgt_5_356;input [WEIGHT_SIZE-1:0] Wgt_5_357;input [WEIGHT_SIZE-1:0] Wgt_5_358;input [WEIGHT_SIZE-1:0] Wgt_5_359;input [WEIGHT_SIZE-1:0] Wgt_5_360;input [WEIGHT_SIZE-1:0] Wgt_5_361;input [WEIGHT_SIZE-1:0] Wgt_5_362;input [WEIGHT_SIZE-1:0] Wgt_5_363;input [WEIGHT_SIZE-1:0] Wgt_5_364;input [WEIGHT_SIZE-1:0] Wgt_5_365;input [WEIGHT_SIZE-1:0] Wgt_5_366;input [WEIGHT_SIZE-1:0] Wgt_5_367;input [WEIGHT_SIZE-1:0] Wgt_5_368;input [WEIGHT_SIZE-1:0] Wgt_5_369;input [WEIGHT_SIZE-1:0] Wgt_5_370;input [WEIGHT_SIZE-1:0] Wgt_5_371;input [WEIGHT_SIZE-1:0] Wgt_5_372;input [WEIGHT_SIZE-1:0] Wgt_5_373;input [WEIGHT_SIZE-1:0] Wgt_5_374;input [WEIGHT_SIZE-1:0] Wgt_5_375;input [WEIGHT_SIZE-1:0] Wgt_5_376;input [WEIGHT_SIZE-1:0] Wgt_5_377;input [WEIGHT_SIZE-1:0] Wgt_5_378;input [WEIGHT_SIZE-1:0] Wgt_5_379;input [WEIGHT_SIZE-1:0] Wgt_5_380;input [WEIGHT_SIZE-1:0] Wgt_5_381;input [WEIGHT_SIZE-1:0] Wgt_5_382;input [WEIGHT_SIZE-1:0] Wgt_5_383;input [WEIGHT_SIZE-1:0] Wgt_5_384;input [WEIGHT_SIZE-1:0] Wgt_5_385;input [WEIGHT_SIZE-1:0] Wgt_5_386;input [WEIGHT_SIZE-1:0] Wgt_5_387;input [WEIGHT_SIZE-1:0] Wgt_5_388;input [WEIGHT_SIZE-1:0] Wgt_5_389;input [WEIGHT_SIZE-1:0] Wgt_5_390;input [WEIGHT_SIZE-1:0] Wgt_5_391;input [WEIGHT_SIZE-1:0] Wgt_5_392;input [WEIGHT_SIZE-1:0] Wgt_5_393;input [WEIGHT_SIZE-1:0] Wgt_5_394;input [WEIGHT_SIZE-1:0] Wgt_5_395;input [WEIGHT_SIZE-1:0] Wgt_5_396;input [WEIGHT_SIZE-1:0] Wgt_5_397;input [WEIGHT_SIZE-1:0] Wgt_5_398;input [WEIGHT_SIZE-1:0] Wgt_5_399;input [WEIGHT_SIZE-1:0] Wgt_5_400;input [WEIGHT_SIZE-1:0] Wgt_5_401;input [WEIGHT_SIZE-1:0] Wgt_5_402;input [WEIGHT_SIZE-1:0] Wgt_5_403;input [WEIGHT_SIZE-1:0] Wgt_5_404;input [WEIGHT_SIZE-1:0] Wgt_5_405;input [WEIGHT_SIZE-1:0] Wgt_5_406;input [WEIGHT_SIZE-1:0] Wgt_5_407;input [WEIGHT_SIZE-1:0] Wgt_5_408;input [WEIGHT_SIZE-1:0] Wgt_5_409;input [WEIGHT_SIZE-1:0] Wgt_5_410;input [WEIGHT_SIZE-1:0] Wgt_5_411;input [WEIGHT_SIZE-1:0] Wgt_5_412;input [WEIGHT_SIZE-1:0] Wgt_5_413;input [WEIGHT_SIZE-1:0] Wgt_5_414;input [WEIGHT_SIZE-1:0] Wgt_5_415;input [WEIGHT_SIZE-1:0] Wgt_5_416;input [WEIGHT_SIZE-1:0] Wgt_5_417;input [WEIGHT_SIZE-1:0] Wgt_5_418;input [WEIGHT_SIZE-1:0] Wgt_5_419;input [WEIGHT_SIZE-1:0] Wgt_5_420;input [WEIGHT_SIZE-1:0] Wgt_5_421;input [WEIGHT_SIZE-1:0] Wgt_5_422;input [WEIGHT_SIZE-1:0] Wgt_5_423;input [WEIGHT_SIZE-1:0] Wgt_5_424;input [WEIGHT_SIZE-1:0] Wgt_5_425;input [WEIGHT_SIZE-1:0] Wgt_5_426;input [WEIGHT_SIZE-1:0] Wgt_5_427;input [WEIGHT_SIZE-1:0] Wgt_5_428;input [WEIGHT_SIZE-1:0] Wgt_5_429;input [WEIGHT_SIZE-1:0] Wgt_5_430;input [WEIGHT_SIZE-1:0] Wgt_5_431;input [WEIGHT_SIZE-1:0] Wgt_5_432;input [WEIGHT_SIZE-1:0] Wgt_5_433;input [WEIGHT_SIZE-1:0] Wgt_5_434;input [WEIGHT_SIZE-1:0] Wgt_5_435;input [WEIGHT_SIZE-1:0] Wgt_5_436;input [WEIGHT_SIZE-1:0] Wgt_5_437;input [WEIGHT_SIZE-1:0] Wgt_5_438;input [WEIGHT_SIZE-1:0] Wgt_5_439;input [WEIGHT_SIZE-1:0] Wgt_5_440;input [WEIGHT_SIZE-1:0] Wgt_5_441;input [WEIGHT_SIZE-1:0] Wgt_5_442;input [WEIGHT_SIZE-1:0] Wgt_5_443;input [WEIGHT_SIZE-1:0] Wgt_5_444;input [WEIGHT_SIZE-1:0] Wgt_5_445;input [WEIGHT_SIZE-1:0] Wgt_5_446;input [WEIGHT_SIZE-1:0] Wgt_5_447;input [WEIGHT_SIZE-1:0] Wgt_5_448;input [WEIGHT_SIZE-1:0] Wgt_5_449;input [WEIGHT_SIZE-1:0] Wgt_5_450;input [WEIGHT_SIZE-1:0] Wgt_5_451;input [WEIGHT_SIZE-1:0] Wgt_5_452;input [WEIGHT_SIZE-1:0] Wgt_5_453;input [WEIGHT_SIZE-1:0] Wgt_5_454;input [WEIGHT_SIZE-1:0] Wgt_5_455;input [WEIGHT_SIZE-1:0] Wgt_5_456;input [WEIGHT_SIZE-1:0] Wgt_5_457;input [WEIGHT_SIZE-1:0] Wgt_5_458;input [WEIGHT_SIZE-1:0] Wgt_5_459;input [WEIGHT_SIZE-1:0] Wgt_5_460;input [WEIGHT_SIZE-1:0] Wgt_5_461;input [WEIGHT_SIZE-1:0] Wgt_5_462;input [WEIGHT_SIZE-1:0] Wgt_5_463;input [WEIGHT_SIZE-1:0] Wgt_5_464;input [WEIGHT_SIZE-1:0] Wgt_5_465;input [WEIGHT_SIZE-1:0] Wgt_5_466;input [WEIGHT_SIZE-1:0] Wgt_5_467;input [WEIGHT_SIZE-1:0] Wgt_5_468;input [WEIGHT_SIZE-1:0] Wgt_5_469;input [WEIGHT_SIZE-1:0] Wgt_5_470;input [WEIGHT_SIZE-1:0] Wgt_5_471;input [WEIGHT_SIZE-1:0] Wgt_5_472;input [WEIGHT_SIZE-1:0] Wgt_5_473;input [WEIGHT_SIZE-1:0] Wgt_5_474;input [WEIGHT_SIZE-1:0] Wgt_5_475;input [WEIGHT_SIZE-1:0] Wgt_5_476;input [WEIGHT_SIZE-1:0] Wgt_5_477;input [WEIGHT_SIZE-1:0] Wgt_5_478;input [WEIGHT_SIZE-1:0] Wgt_5_479;input [WEIGHT_SIZE-1:0] Wgt_5_480;input [WEIGHT_SIZE-1:0] Wgt_5_481;input [WEIGHT_SIZE-1:0] Wgt_5_482;input [WEIGHT_SIZE-1:0] Wgt_5_483;input [WEIGHT_SIZE-1:0] Wgt_5_484;input [WEIGHT_SIZE-1:0] Wgt_5_485;input [WEIGHT_SIZE-1:0] Wgt_5_486;input [WEIGHT_SIZE-1:0] Wgt_5_487;input [WEIGHT_SIZE-1:0] Wgt_5_488;input [WEIGHT_SIZE-1:0] Wgt_5_489;input [WEIGHT_SIZE-1:0] Wgt_5_490;input [WEIGHT_SIZE-1:0] Wgt_5_491;input [WEIGHT_SIZE-1:0] Wgt_5_492;input [WEIGHT_SIZE-1:0] Wgt_5_493;input [WEIGHT_SIZE-1:0] Wgt_5_494;input [WEIGHT_SIZE-1:0] Wgt_5_495;input [WEIGHT_SIZE-1:0] Wgt_5_496;input [WEIGHT_SIZE-1:0] Wgt_5_497;input [WEIGHT_SIZE-1:0] Wgt_5_498;input [WEIGHT_SIZE-1:0] Wgt_5_499;input [WEIGHT_SIZE-1:0] Wgt_5_500;input [WEIGHT_SIZE-1:0] Wgt_5_501;input [WEIGHT_SIZE-1:0] Wgt_5_502;input [WEIGHT_SIZE-1:0] Wgt_5_503;input [WEIGHT_SIZE-1:0] Wgt_5_504;input [WEIGHT_SIZE-1:0] Wgt_5_505;input [WEIGHT_SIZE-1:0] Wgt_5_506;input [WEIGHT_SIZE-1:0] Wgt_5_507;input [WEIGHT_SIZE-1:0] Wgt_5_508;input [WEIGHT_SIZE-1:0] Wgt_5_509;input [WEIGHT_SIZE-1:0] Wgt_5_510;input [WEIGHT_SIZE-1:0] Wgt_5_511;input [WEIGHT_SIZE-1:0] Wgt_5_512;input [WEIGHT_SIZE-1:0] Wgt_5_513;input [WEIGHT_SIZE-1:0] Wgt_5_514;input [WEIGHT_SIZE-1:0] Wgt_5_515;input [WEIGHT_SIZE-1:0] Wgt_5_516;input [WEIGHT_SIZE-1:0] Wgt_5_517;input [WEIGHT_SIZE-1:0] Wgt_5_518;input [WEIGHT_SIZE-1:0] Wgt_5_519;input [WEIGHT_SIZE-1:0] Wgt_5_520;input [WEIGHT_SIZE-1:0] Wgt_5_521;input [WEIGHT_SIZE-1:0] Wgt_5_522;input [WEIGHT_SIZE-1:0] Wgt_5_523;input [WEIGHT_SIZE-1:0] Wgt_5_524;input [WEIGHT_SIZE-1:0] Wgt_5_525;input [WEIGHT_SIZE-1:0] Wgt_5_526;input [WEIGHT_SIZE-1:0] Wgt_5_527;input [WEIGHT_SIZE-1:0] Wgt_5_528;input [WEIGHT_SIZE-1:0] Wgt_5_529;input [WEIGHT_SIZE-1:0] Wgt_5_530;input [WEIGHT_SIZE-1:0] Wgt_5_531;input [WEIGHT_SIZE-1:0] Wgt_5_532;input [WEIGHT_SIZE-1:0] Wgt_5_533;input [WEIGHT_SIZE-1:0] Wgt_5_534;input [WEIGHT_SIZE-1:0] Wgt_5_535;input [WEIGHT_SIZE-1:0] Wgt_5_536;input [WEIGHT_SIZE-1:0] Wgt_5_537;input [WEIGHT_SIZE-1:0] Wgt_5_538;input [WEIGHT_SIZE-1:0] Wgt_5_539;input [WEIGHT_SIZE-1:0] Wgt_5_540;input [WEIGHT_SIZE-1:0] Wgt_5_541;input [WEIGHT_SIZE-1:0] Wgt_5_542;input [WEIGHT_SIZE-1:0] Wgt_5_543;input [WEIGHT_SIZE-1:0] Wgt_5_544;input [WEIGHT_SIZE-1:0] Wgt_5_545;input [WEIGHT_SIZE-1:0] Wgt_5_546;input [WEIGHT_SIZE-1:0] Wgt_5_547;input [WEIGHT_SIZE-1:0] Wgt_5_548;input [WEIGHT_SIZE-1:0] Wgt_5_549;input [WEIGHT_SIZE-1:0] Wgt_5_550;input [WEIGHT_SIZE-1:0] Wgt_5_551;input [WEIGHT_SIZE-1:0] Wgt_5_552;input [WEIGHT_SIZE-1:0] Wgt_5_553;input [WEIGHT_SIZE-1:0] Wgt_5_554;input [WEIGHT_SIZE-1:0] Wgt_5_555;input [WEIGHT_SIZE-1:0] Wgt_5_556;input [WEIGHT_SIZE-1:0] Wgt_5_557;input [WEIGHT_SIZE-1:0] Wgt_5_558;input [WEIGHT_SIZE-1:0] Wgt_5_559;input [WEIGHT_SIZE-1:0] Wgt_5_560;input [WEIGHT_SIZE-1:0] Wgt_5_561;input [WEIGHT_SIZE-1:0] Wgt_5_562;input [WEIGHT_SIZE-1:0] Wgt_5_563;input [WEIGHT_SIZE-1:0] Wgt_5_564;input [WEIGHT_SIZE-1:0] Wgt_5_565;input [WEIGHT_SIZE-1:0] Wgt_5_566;input [WEIGHT_SIZE-1:0] Wgt_5_567;input [WEIGHT_SIZE-1:0] Wgt_5_568;input [WEIGHT_SIZE-1:0] Wgt_5_569;input [WEIGHT_SIZE-1:0] Wgt_5_570;input [WEIGHT_SIZE-1:0] Wgt_5_571;input [WEIGHT_SIZE-1:0] Wgt_5_572;input [WEIGHT_SIZE-1:0] Wgt_5_573;input [WEIGHT_SIZE-1:0] Wgt_5_574;input [WEIGHT_SIZE-1:0] Wgt_5_575;input [WEIGHT_SIZE-1:0] Wgt_5_576;input [WEIGHT_SIZE-1:0] Wgt_5_577;input [WEIGHT_SIZE-1:0] Wgt_5_578;input [WEIGHT_SIZE-1:0] Wgt_5_579;input [WEIGHT_SIZE-1:0] Wgt_5_580;input [WEIGHT_SIZE-1:0] Wgt_5_581;input [WEIGHT_SIZE-1:0] Wgt_5_582;input [WEIGHT_SIZE-1:0] Wgt_5_583;input [WEIGHT_SIZE-1:0] Wgt_5_584;input [WEIGHT_SIZE-1:0] Wgt_5_585;input [WEIGHT_SIZE-1:0] Wgt_5_586;input [WEIGHT_SIZE-1:0] Wgt_5_587;input [WEIGHT_SIZE-1:0] Wgt_5_588;input [WEIGHT_SIZE-1:0] Wgt_5_589;input [WEIGHT_SIZE-1:0] Wgt_5_590;input [WEIGHT_SIZE-1:0] Wgt_5_591;input [WEIGHT_SIZE-1:0] Wgt_5_592;input [WEIGHT_SIZE-1:0] Wgt_5_593;input [WEIGHT_SIZE-1:0] Wgt_5_594;input [WEIGHT_SIZE-1:0] Wgt_5_595;input [WEIGHT_SIZE-1:0] Wgt_5_596;input [WEIGHT_SIZE-1:0] Wgt_5_597;input [WEIGHT_SIZE-1:0] Wgt_5_598;input [WEIGHT_SIZE-1:0] Wgt_5_599;input [WEIGHT_SIZE-1:0] Wgt_5_600;input [WEIGHT_SIZE-1:0] Wgt_5_601;input [WEIGHT_SIZE-1:0] Wgt_5_602;input [WEIGHT_SIZE-1:0] Wgt_5_603;input [WEIGHT_SIZE-1:0] Wgt_5_604;input [WEIGHT_SIZE-1:0] Wgt_5_605;input [WEIGHT_SIZE-1:0] Wgt_5_606;input [WEIGHT_SIZE-1:0] Wgt_5_607;input [WEIGHT_SIZE-1:0] Wgt_5_608;input [WEIGHT_SIZE-1:0] Wgt_5_609;input [WEIGHT_SIZE-1:0] Wgt_5_610;input [WEIGHT_SIZE-1:0] Wgt_5_611;input [WEIGHT_SIZE-1:0] Wgt_5_612;input [WEIGHT_SIZE-1:0] Wgt_5_613;input [WEIGHT_SIZE-1:0] Wgt_5_614;input [WEIGHT_SIZE-1:0] Wgt_5_615;input [WEIGHT_SIZE-1:0] Wgt_5_616;input [WEIGHT_SIZE-1:0] Wgt_5_617;input [WEIGHT_SIZE-1:0] Wgt_5_618;input [WEIGHT_SIZE-1:0] Wgt_5_619;input [WEIGHT_SIZE-1:0] Wgt_5_620;input [WEIGHT_SIZE-1:0] Wgt_5_621;input [WEIGHT_SIZE-1:0] Wgt_5_622;input [WEIGHT_SIZE-1:0] Wgt_5_623;input [WEIGHT_SIZE-1:0] Wgt_5_624;input [WEIGHT_SIZE-1:0] Wgt_5_625;input [WEIGHT_SIZE-1:0] Wgt_5_626;input [WEIGHT_SIZE-1:0] Wgt_5_627;input [WEIGHT_SIZE-1:0] Wgt_5_628;input [WEIGHT_SIZE-1:0] Wgt_5_629;input [WEIGHT_SIZE-1:0] Wgt_5_630;input [WEIGHT_SIZE-1:0] Wgt_5_631;input [WEIGHT_SIZE-1:0] Wgt_5_632;input [WEIGHT_SIZE-1:0] Wgt_5_633;input [WEIGHT_SIZE-1:0] Wgt_5_634;input [WEIGHT_SIZE-1:0] Wgt_5_635;input [WEIGHT_SIZE-1:0] Wgt_5_636;input [WEIGHT_SIZE-1:0] Wgt_5_637;input [WEIGHT_SIZE-1:0] Wgt_5_638;input [WEIGHT_SIZE-1:0] Wgt_5_639;input [WEIGHT_SIZE-1:0] Wgt_5_640;input [WEIGHT_SIZE-1:0] Wgt_5_641;input [WEIGHT_SIZE-1:0] Wgt_5_642;input [WEIGHT_SIZE-1:0] Wgt_5_643;input [WEIGHT_SIZE-1:0] Wgt_5_644;input [WEIGHT_SIZE-1:0] Wgt_5_645;input [WEIGHT_SIZE-1:0] Wgt_5_646;input [WEIGHT_SIZE-1:0] Wgt_5_647;input [WEIGHT_SIZE-1:0] Wgt_5_648;input [WEIGHT_SIZE-1:0] Wgt_5_649;input [WEIGHT_SIZE-1:0] Wgt_5_650;input [WEIGHT_SIZE-1:0] Wgt_5_651;input [WEIGHT_SIZE-1:0] Wgt_5_652;input [WEIGHT_SIZE-1:0] Wgt_5_653;input [WEIGHT_SIZE-1:0] Wgt_5_654;input [WEIGHT_SIZE-1:0] Wgt_5_655;input [WEIGHT_SIZE-1:0] Wgt_5_656;input [WEIGHT_SIZE-1:0] Wgt_5_657;input [WEIGHT_SIZE-1:0] Wgt_5_658;input [WEIGHT_SIZE-1:0] Wgt_5_659;input [WEIGHT_SIZE-1:0] Wgt_5_660;input [WEIGHT_SIZE-1:0] Wgt_5_661;input [WEIGHT_SIZE-1:0] Wgt_5_662;input [WEIGHT_SIZE-1:0] Wgt_5_663;input [WEIGHT_SIZE-1:0] Wgt_5_664;input [WEIGHT_SIZE-1:0] Wgt_5_665;input [WEIGHT_SIZE-1:0] Wgt_5_666;input [WEIGHT_SIZE-1:0] Wgt_5_667;input [WEIGHT_SIZE-1:0] Wgt_5_668;input [WEIGHT_SIZE-1:0] Wgt_5_669;input [WEIGHT_SIZE-1:0] Wgt_5_670;input [WEIGHT_SIZE-1:0] Wgt_5_671;input [WEIGHT_SIZE-1:0] Wgt_5_672;input [WEIGHT_SIZE-1:0] Wgt_5_673;input [WEIGHT_SIZE-1:0] Wgt_5_674;input [WEIGHT_SIZE-1:0] Wgt_5_675;input [WEIGHT_SIZE-1:0] Wgt_5_676;input [WEIGHT_SIZE-1:0] Wgt_5_677;input [WEIGHT_SIZE-1:0] Wgt_5_678;input [WEIGHT_SIZE-1:0] Wgt_5_679;input [WEIGHT_SIZE-1:0] Wgt_5_680;input [WEIGHT_SIZE-1:0] Wgt_5_681;input [WEIGHT_SIZE-1:0] Wgt_5_682;input [WEIGHT_SIZE-1:0] Wgt_5_683;input [WEIGHT_SIZE-1:0] Wgt_5_684;input [WEIGHT_SIZE-1:0] Wgt_5_685;input [WEIGHT_SIZE-1:0] Wgt_5_686;input [WEIGHT_SIZE-1:0] Wgt_5_687;input [WEIGHT_SIZE-1:0] Wgt_5_688;input [WEIGHT_SIZE-1:0] Wgt_5_689;input [WEIGHT_SIZE-1:0] Wgt_5_690;input [WEIGHT_SIZE-1:0] Wgt_5_691;input [WEIGHT_SIZE-1:0] Wgt_5_692;input [WEIGHT_SIZE-1:0] Wgt_5_693;input [WEIGHT_SIZE-1:0] Wgt_5_694;input [WEIGHT_SIZE-1:0] Wgt_5_695;input [WEIGHT_SIZE-1:0] Wgt_5_696;input [WEIGHT_SIZE-1:0] Wgt_5_697;input [WEIGHT_SIZE-1:0] Wgt_5_698;input [WEIGHT_SIZE-1:0] Wgt_5_699;input [WEIGHT_SIZE-1:0] Wgt_5_700;input [WEIGHT_SIZE-1:0] Wgt_5_701;input [WEIGHT_SIZE-1:0] Wgt_5_702;input [WEIGHT_SIZE-1:0] Wgt_5_703;input [WEIGHT_SIZE-1:0] Wgt_5_704;input [WEIGHT_SIZE-1:0] Wgt_5_705;input [WEIGHT_SIZE-1:0] Wgt_5_706;input [WEIGHT_SIZE-1:0] Wgt_5_707;input [WEIGHT_SIZE-1:0] Wgt_5_708;input [WEIGHT_SIZE-1:0] Wgt_5_709;input [WEIGHT_SIZE-1:0] Wgt_5_710;input [WEIGHT_SIZE-1:0] Wgt_5_711;input [WEIGHT_SIZE-1:0] Wgt_5_712;input [WEIGHT_SIZE-1:0] Wgt_5_713;input [WEIGHT_SIZE-1:0] Wgt_5_714;input [WEIGHT_SIZE-1:0] Wgt_5_715;input [WEIGHT_SIZE-1:0] Wgt_5_716;input [WEIGHT_SIZE-1:0] Wgt_5_717;input [WEIGHT_SIZE-1:0] Wgt_5_718;input [WEIGHT_SIZE-1:0] Wgt_5_719;input [WEIGHT_SIZE-1:0] Wgt_5_720;input [WEIGHT_SIZE-1:0] Wgt_5_721;input [WEIGHT_SIZE-1:0] Wgt_5_722;input [WEIGHT_SIZE-1:0] Wgt_5_723;input [WEIGHT_SIZE-1:0] Wgt_5_724;input [WEIGHT_SIZE-1:0] Wgt_5_725;input [WEIGHT_SIZE-1:0] Wgt_5_726;input [WEIGHT_SIZE-1:0] Wgt_5_727;input [WEIGHT_SIZE-1:0] Wgt_5_728;input [WEIGHT_SIZE-1:0] Wgt_5_729;input [WEIGHT_SIZE-1:0] Wgt_5_730;input [WEIGHT_SIZE-1:0] Wgt_5_731;input [WEIGHT_SIZE-1:0] Wgt_5_732;input [WEIGHT_SIZE-1:0] Wgt_5_733;input [WEIGHT_SIZE-1:0] Wgt_5_734;input [WEIGHT_SIZE-1:0] Wgt_5_735;input [WEIGHT_SIZE-1:0] Wgt_5_736;input [WEIGHT_SIZE-1:0] Wgt_5_737;input [WEIGHT_SIZE-1:0] Wgt_5_738;input [WEIGHT_SIZE-1:0] Wgt_5_739;input [WEIGHT_SIZE-1:0] Wgt_5_740;input [WEIGHT_SIZE-1:0] Wgt_5_741;input [WEIGHT_SIZE-1:0] Wgt_5_742;input [WEIGHT_SIZE-1:0] Wgt_5_743;input [WEIGHT_SIZE-1:0] Wgt_5_744;input [WEIGHT_SIZE-1:0] Wgt_5_745;input [WEIGHT_SIZE-1:0] Wgt_5_746;input [WEIGHT_SIZE-1:0] Wgt_5_747;input [WEIGHT_SIZE-1:0] Wgt_5_748;input [WEIGHT_SIZE-1:0] Wgt_5_749;input [WEIGHT_SIZE-1:0] Wgt_5_750;input [WEIGHT_SIZE-1:0] Wgt_5_751;input [WEIGHT_SIZE-1:0] Wgt_5_752;input [WEIGHT_SIZE-1:0] Wgt_5_753;input [WEIGHT_SIZE-1:0] Wgt_5_754;input [WEIGHT_SIZE-1:0] Wgt_5_755;input [WEIGHT_SIZE-1:0] Wgt_5_756;input [WEIGHT_SIZE-1:0] Wgt_5_757;input [WEIGHT_SIZE-1:0] Wgt_5_758;input [WEIGHT_SIZE-1:0] Wgt_5_759;input [WEIGHT_SIZE-1:0] Wgt_5_760;input [WEIGHT_SIZE-1:0] Wgt_5_761;input [WEIGHT_SIZE-1:0] Wgt_5_762;input [WEIGHT_SIZE-1:0] Wgt_5_763;input [WEIGHT_SIZE-1:0] Wgt_5_764;input [WEIGHT_SIZE-1:0] Wgt_5_765;input [WEIGHT_SIZE-1:0] Wgt_5_766;input [WEIGHT_SIZE-1:0] Wgt_5_767;input [WEIGHT_SIZE-1:0] Wgt_5_768;input [WEIGHT_SIZE-1:0] Wgt_5_769;input [WEIGHT_SIZE-1:0] Wgt_5_770;input [WEIGHT_SIZE-1:0] Wgt_5_771;input [WEIGHT_SIZE-1:0] Wgt_5_772;input [WEIGHT_SIZE-1:0] Wgt_5_773;input [WEIGHT_SIZE-1:0] Wgt_5_774;input [WEIGHT_SIZE-1:0] Wgt_5_775;input [WEIGHT_SIZE-1:0] Wgt_5_776;input [WEIGHT_SIZE-1:0] Wgt_5_777;input [WEIGHT_SIZE-1:0] Wgt_5_778;input [WEIGHT_SIZE-1:0] Wgt_5_779;input [WEIGHT_SIZE-1:0] Wgt_5_780;input [WEIGHT_SIZE-1:0] Wgt_5_781;input [WEIGHT_SIZE-1:0] Wgt_5_782;input [WEIGHT_SIZE-1:0] Wgt_5_783;input [WEIGHT_SIZE-1:0] Wgt_5_784;input [WEIGHT_SIZE-1:0] Wgt_6_0;input [WEIGHT_SIZE-1:0] Wgt_6_1;input [WEIGHT_SIZE-1:0] Wgt_6_2;input [WEIGHT_SIZE-1:0] Wgt_6_3;input [WEIGHT_SIZE-1:0] Wgt_6_4;input [WEIGHT_SIZE-1:0] Wgt_6_5;input [WEIGHT_SIZE-1:0] Wgt_6_6;input [WEIGHT_SIZE-1:0] Wgt_6_7;input [WEIGHT_SIZE-1:0] Wgt_6_8;input [WEIGHT_SIZE-1:0] Wgt_6_9;input [WEIGHT_SIZE-1:0] Wgt_6_10;input [WEIGHT_SIZE-1:0] Wgt_6_11;input [WEIGHT_SIZE-1:0] Wgt_6_12;input [WEIGHT_SIZE-1:0] Wgt_6_13;input [WEIGHT_SIZE-1:0] Wgt_6_14;input [WEIGHT_SIZE-1:0] Wgt_6_15;input [WEIGHT_SIZE-1:0] Wgt_6_16;input [WEIGHT_SIZE-1:0] Wgt_6_17;input [WEIGHT_SIZE-1:0] Wgt_6_18;input [WEIGHT_SIZE-1:0] Wgt_6_19;input [WEIGHT_SIZE-1:0] Wgt_6_20;input [WEIGHT_SIZE-1:0] Wgt_6_21;input [WEIGHT_SIZE-1:0] Wgt_6_22;input [WEIGHT_SIZE-1:0] Wgt_6_23;input [WEIGHT_SIZE-1:0] Wgt_6_24;input [WEIGHT_SIZE-1:0] Wgt_6_25;input [WEIGHT_SIZE-1:0] Wgt_6_26;input [WEIGHT_SIZE-1:0] Wgt_6_27;input [WEIGHT_SIZE-1:0] Wgt_6_28;input [WEIGHT_SIZE-1:0] Wgt_6_29;input [WEIGHT_SIZE-1:0] Wgt_6_30;input [WEIGHT_SIZE-1:0] Wgt_6_31;input [WEIGHT_SIZE-1:0] Wgt_6_32;input [WEIGHT_SIZE-1:0] Wgt_6_33;input [WEIGHT_SIZE-1:0] Wgt_6_34;input [WEIGHT_SIZE-1:0] Wgt_6_35;input [WEIGHT_SIZE-1:0] Wgt_6_36;input [WEIGHT_SIZE-1:0] Wgt_6_37;input [WEIGHT_SIZE-1:0] Wgt_6_38;input [WEIGHT_SIZE-1:0] Wgt_6_39;input [WEIGHT_SIZE-1:0] Wgt_6_40;input [WEIGHT_SIZE-1:0] Wgt_6_41;input [WEIGHT_SIZE-1:0] Wgt_6_42;input [WEIGHT_SIZE-1:0] Wgt_6_43;input [WEIGHT_SIZE-1:0] Wgt_6_44;input [WEIGHT_SIZE-1:0] Wgt_6_45;input [WEIGHT_SIZE-1:0] Wgt_6_46;input [WEIGHT_SIZE-1:0] Wgt_6_47;input [WEIGHT_SIZE-1:0] Wgt_6_48;input [WEIGHT_SIZE-1:0] Wgt_6_49;input [WEIGHT_SIZE-1:0] Wgt_6_50;input [WEIGHT_SIZE-1:0] Wgt_6_51;input [WEIGHT_SIZE-1:0] Wgt_6_52;input [WEIGHT_SIZE-1:0] Wgt_6_53;input [WEIGHT_SIZE-1:0] Wgt_6_54;input [WEIGHT_SIZE-1:0] Wgt_6_55;input [WEIGHT_SIZE-1:0] Wgt_6_56;input [WEIGHT_SIZE-1:0] Wgt_6_57;input [WEIGHT_SIZE-1:0] Wgt_6_58;input [WEIGHT_SIZE-1:0] Wgt_6_59;input [WEIGHT_SIZE-1:0] Wgt_6_60;input [WEIGHT_SIZE-1:0] Wgt_6_61;input [WEIGHT_SIZE-1:0] Wgt_6_62;input [WEIGHT_SIZE-1:0] Wgt_6_63;input [WEIGHT_SIZE-1:0] Wgt_6_64;input [WEIGHT_SIZE-1:0] Wgt_6_65;input [WEIGHT_SIZE-1:0] Wgt_6_66;input [WEIGHT_SIZE-1:0] Wgt_6_67;input [WEIGHT_SIZE-1:0] Wgt_6_68;input [WEIGHT_SIZE-1:0] Wgt_6_69;input [WEIGHT_SIZE-1:0] Wgt_6_70;input [WEIGHT_SIZE-1:0] Wgt_6_71;input [WEIGHT_SIZE-1:0] Wgt_6_72;input [WEIGHT_SIZE-1:0] Wgt_6_73;input [WEIGHT_SIZE-1:0] Wgt_6_74;input [WEIGHT_SIZE-1:0] Wgt_6_75;input [WEIGHT_SIZE-1:0] Wgt_6_76;input [WEIGHT_SIZE-1:0] Wgt_6_77;input [WEIGHT_SIZE-1:0] Wgt_6_78;input [WEIGHT_SIZE-1:0] Wgt_6_79;input [WEIGHT_SIZE-1:0] Wgt_6_80;input [WEIGHT_SIZE-1:0] Wgt_6_81;input [WEIGHT_SIZE-1:0] Wgt_6_82;input [WEIGHT_SIZE-1:0] Wgt_6_83;input [WEIGHT_SIZE-1:0] Wgt_6_84;input [WEIGHT_SIZE-1:0] Wgt_6_85;input [WEIGHT_SIZE-1:0] Wgt_6_86;input [WEIGHT_SIZE-1:0] Wgt_6_87;input [WEIGHT_SIZE-1:0] Wgt_6_88;input [WEIGHT_SIZE-1:0] Wgt_6_89;input [WEIGHT_SIZE-1:0] Wgt_6_90;input [WEIGHT_SIZE-1:0] Wgt_6_91;input [WEIGHT_SIZE-1:0] Wgt_6_92;input [WEIGHT_SIZE-1:0] Wgt_6_93;input [WEIGHT_SIZE-1:0] Wgt_6_94;input [WEIGHT_SIZE-1:0] Wgt_6_95;input [WEIGHT_SIZE-1:0] Wgt_6_96;input [WEIGHT_SIZE-1:0] Wgt_6_97;input [WEIGHT_SIZE-1:0] Wgt_6_98;input [WEIGHT_SIZE-1:0] Wgt_6_99;input [WEIGHT_SIZE-1:0] Wgt_6_100;input [WEIGHT_SIZE-1:0] Wgt_6_101;input [WEIGHT_SIZE-1:0] Wgt_6_102;input [WEIGHT_SIZE-1:0] Wgt_6_103;input [WEIGHT_SIZE-1:0] Wgt_6_104;input [WEIGHT_SIZE-1:0] Wgt_6_105;input [WEIGHT_SIZE-1:0] Wgt_6_106;input [WEIGHT_SIZE-1:0] Wgt_6_107;input [WEIGHT_SIZE-1:0] Wgt_6_108;input [WEIGHT_SIZE-1:0] Wgt_6_109;input [WEIGHT_SIZE-1:0] Wgt_6_110;input [WEIGHT_SIZE-1:0] Wgt_6_111;input [WEIGHT_SIZE-1:0] Wgt_6_112;input [WEIGHT_SIZE-1:0] Wgt_6_113;input [WEIGHT_SIZE-1:0] Wgt_6_114;input [WEIGHT_SIZE-1:0] Wgt_6_115;input [WEIGHT_SIZE-1:0] Wgt_6_116;input [WEIGHT_SIZE-1:0] Wgt_6_117;input [WEIGHT_SIZE-1:0] Wgt_6_118;input [WEIGHT_SIZE-1:0] Wgt_6_119;input [WEIGHT_SIZE-1:0] Wgt_6_120;input [WEIGHT_SIZE-1:0] Wgt_6_121;input [WEIGHT_SIZE-1:0] Wgt_6_122;input [WEIGHT_SIZE-1:0] Wgt_6_123;input [WEIGHT_SIZE-1:0] Wgt_6_124;input [WEIGHT_SIZE-1:0] Wgt_6_125;input [WEIGHT_SIZE-1:0] Wgt_6_126;input [WEIGHT_SIZE-1:0] Wgt_6_127;input [WEIGHT_SIZE-1:0] Wgt_6_128;input [WEIGHT_SIZE-1:0] Wgt_6_129;input [WEIGHT_SIZE-1:0] Wgt_6_130;input [WEIGHT_SIZE-1:0] Wgt_6_131;input [WEIGHT_SIZE-1:0] Wgt_6_132;input [WEIGHT_SIZE-1:0] Wgt_6_133;input [WEIGHT_SIZE-1:0] Wgt_6_134;input [WEIGHT_SIZE-1:0] Wgt_6_135;input [WEIGHT_SIZE-1:0] Wgt_6_136;input [WEIGHT_SIZE-1:0] Wgt_6_137;input [WEIGHT_SIZE-1:0] Wgt_6_138;input [WEIGHT_SIZE-1:0] Wgt_6_139;input [WEIGHT_SIZE-1:0] Wgt_6_140;input [WEIGHT_SIZE-1:0] Wgt_6_141;input [WEIGHT_SIZE-1:0] Wgt_6_142;input [WEIGHT_SIZE-1:0] Wgt_6_143;input [WEIGHT_SIZE-1:0] Wgt_6_144;input [WEIGHT_SIZE-1:0] Wgt_6_145;input [WEIGHT_SIZE-1:0] Wgt_6_146;input [WEIGHT_SIZE-1:0] Wgt_6_147;input [WEIGHT_SIZE-1:0] Wgt_6_148;input [WEIGHT_SIZE-1:0] Wgt_6_149;input [WEIGHT_SIZE-1:0] Wgt_6_150;input [WEIGHT_SIZE-1:0] Wgt_6_151;input [WEIGHT_SIZE-1:0] Wgt_6_152;input [WEIGHT_SIZE-1:0] Wgt_6_153;input [WEIGHT_SIZE-1:0] Wgt_6_154;input [WEIGHT_SIZE-1:0] Wgt_6_155;input [WEIGHT_SIZE-1:0] Wgt_6_156;input [WEIGHT_SIZE-1:0] Wgt_6_157;input [WEIGHT_SIZE-1:0] Wgt_6_158;input [WEIGHT_SIZE-1:0] Wgt_6_159;input [WEIGHT_SIZE-1:0] Wgt_6_160;input [WEIGHT_SIZE-1:0] Wgt_6_161;input [WEIGHT_SIZE-1:0] Wgt_6_162;input [WEIGHT_SIZE-1:0] Wgt_6_163;input [WEIGHT_SIZE-1:0] Wgt_6_164;input [WEIGHT_SIZE-1:0] Wgt_6_165;input [WEIGHT_SIZE-1:0] Wgt_6_166;input [WEIGHT_SIZE-1:0] Wgt_6_167;input [WEIGHT_SIZE-1:0] Wgt_6_168;input [WEIGHT_SIZE-1:0] Wgt_6_169;input [WEIGHT_SIZE-1:0] Wgt_6_170;input [WEIGHT_SIZE-1:0] Wgt_6_171;input [WEIGHT_SIZE-1:0] Wgt_6_172;input [WEIGHT_SIZE-1:0] Wgt_6_173;input [WEIGHT_SIZE-1:0] Wgt_6_174;input [WEIGHT_SIZE-1:0] Wgt_6_175;input [WEIGHT_SIZE-1:0] Wgt_6_176;input [WEIGHT_SIZE-1:0] Wgt_6_177;input [WEIGHT_SIZE-1:0] Wgt_6_178;input [WEIGHT_SIZE-1:0] Wgt_6_179;input [WEIGHT_SIZE-1:0] Wgt_6_180;input [WEIGHT_SIZE-1:0] Wgt_6_181;input [WEIGHT_SIZE-1:0] Wgt_6_182;input [WEIGHT_SIZE-1:0] Wgt_6_183;input [WEIGHT_SIZE-1:0] Wgt_6_184;input [WEIGHT_SIZE-1:0] Wgt_6_185;input [WEIGHT_SIZE-1:0] Wgt_6_186;input [WEIGHT_SIZE-1:0] Wgt_6_187;input [WEIGHT_SIZE-1:0] Wgt_6_188;input [WEIGHT_SIZE-1:0] Wgt_6_189;input [WEIGHT_SIZE-1:0] Wgt_6_190;input [WEIGHT_SIZE-1:0] Wgt_6_191;input [WEIGHT_SIZE-1:0] Wgt_6_192;input [WEIGHT_SIZE-1:0] Wgt_6_193;input [WEIGHT_SIZE-1:0] Wgt_6_194;input [WEIGHT_SIZE-1:0] Wgt_6_195;input [WEIGHT_SIZE-1:0] Wgt_6_196;input [WEIGHT_SIZE-1:0] Wgt_6_197;input [WEIGHT_SIZE-1:0] Wgt_6_198;input [WEIGHT_SIZE-1:0] Wgt_6_199;input [WEIGHT_SIZE-1:0] Wgt_6_200;input [WEIGHT_SIZE-1:0] Wgt_6_201;input [WEIGHT_SIZE-1:0] Wgt_6_202;input [WEIGHT_SIZE-1:0] Wgt_6_203;input [WEIGHT_SIZE-1:0] Wgt_6_204;input [WEIGHT_SIZE-1:0] Wgt_6_205;input [WEIGHT_SIZE-1:0] Wgt_6_206;input [WEIGHT_SIZE-1:0] Wgt_6_207;input [WEIGHT_SIZE-1:0] Wgt_6_208;input [WEIGHT_SIZE-1:0] Wgt_6_209;input [WEIGHT_SIZE-1:0] Wgt_6_210;input [WEIGHT_SIZE-1:0] Wgt_6_211;input [WEIGHT_SIZE-1:0] Wgt_6_212;input [WEIGHT_SIZE-1:0] Wgt_6_213;input [WEIGHT_SIZE-1:0] Wgt_6_214;input [WEIGHT_SIZE-1:0] Wgt_6_215;input [WEIGHT_SIZE-1:0] Wgt_6_216;input [WEIGHT_SIZE-1:0] Wgt_6_217;input [WEIGHT_SIZE-1:0] Wgt_6_218;input [WEIGHT_SIZE-1:0] Wgt_6_219;input [WEIGHT_SIZE-1:0] Wgt_6_220;input [WEIGHT_SIZE-1:0] Wgt_6_221;input [WEIGHT_SIZE-1:0] Wgt_6_222;input [WEIGHT_SIZE-1:0] Wgt_6_223;input [WEIGHT_SIZE-1:0] Wgt_6_224;input [WEIGHT_SIZE-1:0] Wgt_6_225;input [WEIGHT_SIZE-1:0] Wgt_6_226;input [WEIGHT_SIZE-1:0] Wgt_6_227;input [WEIGHT_SIZE-1:0] Wgt_6_228;input [WEIGHT_SIZE-1:0] Wgt_6_229;input [WEIGHT_SIZE-1:0] Wgt_6_230;input [WEIGHT_SIZE-1:0] Wgt_6_231;input [WEIGHT_SIZE-1:0] Wgt_6_232;input [WEIGHT_SIZE-1:0] Wgt_6_233;input [WEIGHT_SIZE-1:0] Wgt_6_234;input [WEIGHT_SIZE-1:0] Wgt_6_235;input [WEIGHT_SIZE-1:0] Wgt_6_236;input [WEIGHT_SIZE-1:0] Wgt_6_237;input [WEIGHT_SIZE-1:0] Wgt_6_238;input [WEIGHT_SIZE-1:0] Wgt_6_239;input [WEIGHT_SIZE-1:0] Wgt_6_240;input [WEIGHT_SIZE-1:0] Wgt_6_241;input [WEIGHT_SIZE-1:0] Wgt_6_242;input [WEIGHT_SIZE-1:0] Wgt_6_243;input [WEIGHT_SIZE-1:0] Wgt_6_244;input [WEIGHT_SIZE-1:0] Wgt_6_245;input [WEIGHT_SIZE-1:0] Wgt_6_246;input [WEIGHT_SIZE-1:0] Wgt_6_247;input [WEIGHT_SIZE-1:0] Wgt_6_248;input [WEIGHT_SIZE-1:0] Wgt_6_249;input [WEIGHT_SIZE-1:0] Wgt_6_250;input [WEIGHT_SIZE-1:0] Wgt_6_251;input [WEIGHT_SIZE-1:0] Wgt_6_252;input [WEIGHT_SIZE-1:0] Wgt_6_253;input [WEIGHT_SIZE-1:0] Wgt_6_254;input [WEIGHT_SIZE-1:0] Wgt_6_255;input [WEIGHT_SIZE-1:0] Wgt_6_256;input [WEIGHT_SIZE-1:0] Wgt_6_257;input [WEIGHT_SIZE-1:0] Wgt_6_258;input [WEIGHT_SIZE-1:0] Wgt_6_259;input [WEIGHT_SIZE-1:0] Wgt_6_260;input [WEIGHT_SIZE-1:0] Wgt_6_261;input [WEIGHT_SIZE-1:0] Wgt_6_262;input [WEIGHT_SIZE-1:0] Wgt_6_263;input [WEIGHT_SIZE-1:0] Wgt_6_264;input [WEIGHT_SIZE-1:0] Wgt_6_265;input [WEIGHT_SIZE-1:0] Wgt_6_266;input [WEIGHT_SIZE-1:0] Wgt_6_267;input [WEIGHT_SIZE-1:0] Wgt_6_268;input [WEIGHT_SIZE-1:0] Wgt_6_269;input [WEIGHT_SIZE-1:0] Wgt_6_270;input [WEIGHT_SIZE-1:0] Wgt_6_271;input [WEIGHT_SIZE-1:0] Wgt_6_272;input [WEIGHT_SIZE-1:0] Wgt_6_273;input [WEIGHT_SIZE-1:0] Wgt_6_274;input [WEIGHT_SIZE-1:0] Wgt_6_275;input [WEIGHT_SIZE-1:0] Wgt_6_276;input [WEIGHT_SIZE-1:0] Wgt_6_277;input [WEIGHT_SIZE-1:0] Wgt_6_278;input [WEIGHT_SIZE-1:0] Wgt_6_279;input [WEIGHT_SIZE-1:0] Wgt_6_280;input [WEIGHT_SIZE-1:0] Wgt_6_281;input [WEIGHT_SIZE-1:0] Wgt_6_282;input [WEIGHT_SIZE-1:0] Wgt_6_283;input [WEIGHT_SIZE-1:0] Wgt_6_284;input [WEIGHT_SIZE-1:0] Wgt_6_285;input [WEIGHT_SIZE-1:0] Wgt_6_286;input [WEIGHT_SIZE-1:0] Wgt_6_287;input [WEIGHT_SIZE-1:0] Wgt_6_288;input [WEIGHT_SIZE-1:0] Wgt_6_289;input [WEIGHT_SIZE-1:0] Wgt_6_290;input [WEIGHT_SIZE-1:0] Wgt_6_291;input [WEIGHT_SIZE-1:0] Wgt_6_292;input [WEIGHT_SIZE-1:0] Wgt_6_293;input [WEIGHT_SIZE-1:0] Wgt_6_294;input [WEIGHT_SIZE-1:0] Wgt_6_295;input [WEIGHT_SIZE-1:0] Wgt_6_296;input [WEIGHT_SIZE-1:0] Wgt_6_297;input [WEIGHT_SIZE-1:0] Wgt_6_298;input [WEIGHT_SIZE-1:0] Wgt_6_299;input [WEIGHT_SIZE-1:0] Wgt_6_300;input [WEIGHT_SIZE-1:0] Wgt_6_301;input [WEIGHT_SIZE-1:0] Wgt_6_302;input [WEIGHT_SIZE-1:0] Wgt_6_303;input [WEIGHT_SIZE-1:0] Wgt_6_304;input [WEIGHT_SIZE-1:0] Wgt_6_305;input [WEIGHT_SIZE-1:0] Wgt_6_306;input [WEIGHT_SIZE-1:0] Wgt_6_307;input [WEIGHT_SIZE-1:0] Wgt_6_308;input [WEIGHT_SIZE-1:0] Wgt_6_309;input [WEIGHT_SIZE-1:0] Wgt_6_310;input [WEIGHT_SIZE-1:0] Wgt_6_311;input [WEIGHT_SIZE-1:0] Wgt_6_312;input [WEIGHT_SIZE-1:0] Wgt_6_313;input [WEIGHT_SIZE-1:0] Wgt_6_314;input [WEIGHT_SIZE-1:0] Wgt_6_315;input [WEIGHT_SIZE-1:0] Wgt_6_316;input [WEIGHT_SIZE-1:0] Wgt_6_317;input [WEIGHT_SIZE-1:0] Wgt_6_318;input [WEIGHT_SIZE-1:0] Wgt_6_319;input [WEIGHT_SIZE-1:0] Wgt_6_320;input [WEIGHT_SIZE-1:0] Wgt_6_321;input [WEIGHT_SIZE-1:0] Wgt_6_322;input [WEIGHT_SIZE-1:0] Wgt_6_323;input [WEIGHT_SIZE-1:0] Wgt_6_324;input [WEIGHT_SIZE-1:0] Wgt_6_325;input [WEIGHT_SIZE-1:0] Wgt_6_326;input [WEIGHT_SIZE-1:0] Wgt_6_327;input [WEIGHT_SIZE-1:0] Wgt_6_328;input [WEIGHT_SIZE-1:0] Wgt_6_329;input [WEIGHT_SIZE-1:0] Wgt_6_330;input [WEIGHT_SIZE-1:0] Wgt_6_331;input [WEIGHT_SIZE-1:0] Wgt_6_332;input [WEIGHT_SIZE-1:0] Wgt_6_333;input [WEIGHT_SIZE-1:0] Wgt_6_334;input [WEIGHT_SIZE-1:0] Wgt_6_335;input [WEIGHT_SIZE-1:0] Wgt_6_336;input [WEIGHT_SIZE-1:0] Wgt_6_337;input [WEIGHT_SIZE-1:0] Wgt_6_338;input [WEIGHT_SIZE-1:0] Wgt_6_339;input [WEIGHT_SIZE-1:0] Wgt_6_340;input [WEIGHT_SIZE-1:0] Wgt_6_341;input [WEIGHT_SIZE-1:0] Wgt_6_342;input [WEIGHT_SIZE-1:0] Wgt_6_343;input [WEIGHT_SIZE-1:0] Wgt_6_344;input [WEIGHT_SIZE-1:0] Wgt_6_345;input [WEIGHT_SIZE-1:0] Wgt_6_346;input [WEIGHT_SIZE-1:0] Wgt_6_347;input [WEIGHT_SIZE-1:0] Wgt_6_348;input [WEIGHT_SIZE-1:0] Wgt_6_349;input [WEIGHT_SIZE-1:0] Wgt_6_350;input [WEIGHT_SIZE-1:0] Wgt_6_351;input [WEIGHT_SIZE-1:0] Wgt_6_352;input [WEIGHT_SIZE-1:0] Wgt_6_353;input [WEIGHT_SIZE-1:0] Wgt_6_354;input [WEIGHT_SIZE-1:0] Wgt_6_355;input [WEIGHT_SIZE-1:0] Wgt_6_356;input [WEIGHT_SIZE-1:0] Wgt_6_357;input [WEIGHT_SIZE-1:0] Wgt_6_358;input [WEIGHT_SIZE-1:0] Wgt_6_359;input [WEIGHT_SIZE-1:0] Wgt_6_360;input [WEIGHT_SIZE-1:0] Wgt_6_361;input [WEIGHT_SIZE-1:0] Wgt_6_362;input [WEIGHT_SIZE-1:0] Wgt_6_363;input [WEIGHT_SIZE-1:0] Wgt_6_364;input [WEIGHT_SIZE-1:0] Wgt_6_365;input [WEIGHT_SIZE-1:0] Wgt_6_366;input [WEIGHT_SIZE-1:0] Wgt_6_367;input [WEIGHT_SIZE-1:0] Wgt_6_368;input [WEIGHT_SIZE-1:0] Wgt_6_369;input [WEIGHT_SIZE-1:0] Wgt_6_370;input [WEIGHT_SIZE-1:0] Wgt_6_371;input [WEIGHT_SIZE-1:0] Wgt_6_372;input [WEIGHT_SIZE-1:0] Wgt_6_373;input [WEIGHT_SIZE-1:0] Wgt_6_374;input [WEIGHT_SIZE-1:0] Wgt_6_375;input [WEIGHT_SIZE-1:0] Wgt_6_376;input [WEIGHT_SIZE-1:0] Wgt_6_377;input [WEIGHT_SIZE-1:0] Wgt_6_378;input [WEIGHT_SIZE-1:0] Wgt_6_379;input [WEIGHT_SIZE-1:0] Wgt_6_380;input [WEIGHT_SIZE-1:0] Wgt_6_381;input [WEIGHT_SIZE-1:0] Wgt_6_382;input [WEIGHT_SIZE-1:0] Wgt_6_383;input [WEIGHT_SIZE-1:0] Wgt_6_384;input [WEIGHT_SIZE-1:0] Wgt_6_385;input [WEIGHT_SIZE-1:0] Wgt_6_386;input [WEIGHT_SIZE-1:0] Wgt_6_387;input [WEIGHT_SIZE-1:0] Wgt_6_388;input [WEIGHT_SIZE-1:0] Wgt_6_389;input [WEIGHT_SIZE-1:0] Wgt_6_390;input [WEIGHT_SIZE-1:0] Wgt_6_391;input [WEIGHT_SIZE-1:0] Wgt_6_392;input [WEIGHT_SIZE-1:0] Wgt_6_393;input [WEIGHT_SIZE-1:0] Wgt_6_394;input [WEIGHT_SIZE-1:0] Wgt_6_395;input [WEIGHT_SIZE-1:0] Wgt_6_396;input [WEIGHT_SIZE-1:0] Wgt_6_397;input [WEIGHT_SIZE-1:0] Wgt_6_398;input [WEIGHT_SIZE-1:0] Wgt_6_399;input [WEIGHT_SIZE-1:0] Wgt_6_400;input [WEIGHT_SIZE-1:0] Wgt_6_401;input [WEIGHT_SIZE-1:0] Wgt_6_402;input [WEIGHT_SIZE-1:0] Wgt_6_403;input [WEIGHT_SIZE-1:0] Wgt_6_404;input [WEIGHT_SIZE-1:0] Wgt_6_405;input [WEIGHT_SIZE-1:0] Wgt_6_406;input [WEIGHT_SIZE-1:0] Wgt_6_407;input [WEIGHT_SIZE-1:0] Wgt_6_408;input [WEIGHT_SIZE-1:0] Wgt_6_409;input [WEIGHT_SIZE-1:0] Wgt_6_410;input [WEIGHT_SIZE-1:0] Wgt_6_411;input [WEIGHT_SIZE-1:0] Wgt_6_412;input [WEIGHT_SIZE-1:0] Wgt_6_413;input [WEIGHT_SIZE-1:0] Wgt_6_414;input [WEIGHT_SIZE-1:0] Wgt_6_415;input [WEIGHT_SIZE-1:0] Wgt_6_416;input [WEIGHT_SIZE-1:0] Wgt_6_417;input [WEIGHT_SIZE-1:0] Wgt_6_418;input [WEIGHT_SIZE-1:0] Wgt_6_419;input [WEIGHT_SIZE-1:0] Wgt_6_420;input [WEIGHT_SIZE-1:0] Wgt_6_421;input [WEIGHT_SIZE-1:0] Wgt_6_422;input [WEIGHT_SIZE-1:0] Wgt_6_423;input [WEIGHT_SIZE-1:0] Wgt_6_424;input [WEIGHT_SIZE-1:0] Wgt_6_425;input [WEIGHT_SIZE-1:0] Wgt_6_426;input [WEIGHT_SIZE-1:0] Wgt_6_427;input [WEIGHT_SIZE-1:0] Wgt_6_428;input [WEIGHT_SIZE-1:0] Wgt_6_429;input [WEIGHT_SIZE-1:0] Wgt_6_430;input [WEIGHT_SIZE-1:0] Wgt_6_431;input [WEIGHT_SIZE-1:0] Wgt_6_432;input [WEIGHT_SIZE-1:0] Wgt_6_433;input [WEIGHT_SIZE-1:0] Wgt_6_434;input [WEIGHT_SIZE-1:0] Wgt_6_435;input [WEIGHT_SIZE-1:0] Wgt_6_436;input [WEIGHT_SIZE-1:0] Wgt_6_437;input [WEIGHT_SIZE-1:0] Wgt_6_438;input [WEIGHT_SIZE-1:0] Wgt_6_439;input [WEIGHT_SIZE-1:0] Wgt_6_440;input [WEIGHT_SIZE-1:0] Wgt_6_441;input [WEIGHT_SIZE-1:0] Wgt_6_442;input [WEIGHT_SIZE-1:0] Wgt_6_443;input [WEIGHT_SIZE-1:0] Wgt_6_444;input [WEIGHT_SIZE-1:0] Wgt_6_445;input [WEIGHT_SIZE-1:0] Wgt_6_446;input [WEIGHT_SIZE-1:0] Wgt_6_447;input [WEIGHT_SIZE-1:0] Wgt_6_448;input [WEIGHT_SIZE-1:0] Wgt_6_449;input [WEIGHT_SIZE-1:0] Wgt_6_450;input [WEIGHT_SIZE-1:0] Wgt_6_451;input [WEIGHT_SIZE-1:0] Wgt_6_452;input [WEIGHT_SIZE-1:0] Wgt_6_453;input [WEIGHT_SIZE-1:0] Wgt_6_454;input [WEIGHT_SIZE-1:0] Wgt_6_455;input [WEIGHT_SIZE-1:0] Wgt_6_456;input [WEIGHT_SIZE-1:0] Wgt_6_457;input [WEIGHT_SIZE-1:0] Wgt_6_458;input [WEIGHT_SIZE-1:0] Wgt_6_459;input [WEIGHT_SIZE-1:0] Wgt_6_460;input [WEIGHT_SIZE-1:0] Wgt_6_461;input [WEIGHT_SIZE-1:0] Wgt_6_462;input [WEIGHT_SIZE-1:0] Wgt_6_463;input [WEIGHT_SIZE-1:0] Wgt_6_464;input [WEIGHT_SIZE-1:0] Wgt_6_465;input [WEIGHT_SIZE-1:0] Wgt_6_466;input [WEIGHT_SIZE-1:0] Wgt_6_467;input [WEIGHT_SIZE-1:0] Wgt_6_468;input [WEIGHT_SIZE-1:0] Wgt_6_469;input [WEIGHT_SIZE-1:0] Wgt_6_470;input [WEIGHT_SIZE-1:0] Wgt_6_471;input [WEIGHT_SIZE-1:0] Wgt_6_472;input [WEIGHT_SIZE-1:0] Wgt_6_473;input [WEIGHT_SIZE-1:0] Wgt_6_474;input [WEIGHT_SIZE-1:0] Wgt_6_475;input [WEIGHT_SIZE-1:0] Wgt_6_476;input [WEIGHT_SIZE-1:0] Wgt_6_477;input [WEIGHT_SIZE-1:0] Wgt_6_478;input [WEIGHT_SIZE-1:0] Wgt_6_479;input [WEIGHT_SIZE-1:0] Wgt_6_480;input [WEIGHT_SIZE-1:0] Wgt_6_481;input [WEIGHT_SIZE-1:0] Wgt_6_482;input [WEIGHT_SIZE-1:0] Wgt_6_483;input [WEIGHT_SIZE-1:0] Wgt_6_484;input [WEIGHT_SIZE-1:0] Wgt_6_485;input [WEIGHT_SIZE-1:0] Wgt_6_486;input [WEIGHT_SIZE-1:0] Wgt_6_487;input [WEIGHT_SIZE-1:0] Wgt_6_488;input [WEIGHT_SIZE-1:0] Wgt_6_489;input [WEIGHT_SIZE-1:0] Wgt_6_490;input [WEIGHT_SIZE-1:0] Wgt_6_491;input [WEIGHT_SIZE-1:0] Wgt_6_492;input [WEIGHT_SIZE-1:0] Wgt_6_493;input [WEIGHT_SIZE-1:0] Wgt_6_494;input [WEIGHT_SIZE-1:0] Wgt_6_495;input [WEIGHT_SIZE-1:0] Wgt_6_496;input [WEIGHT_SIZE-1:0] Wgt_6_497;input [WEIGHT_SIZE-1:0] Wgt_6_498;input [WEIGHT_SIZE-1:0] Wgt_6_499;input [WEIGHT_SIZE-1:0] Wgt_6_500;input [WEIGHT_SIZE-1:0] Wgt_6_501;input [WEIGHT_SIZE-1:0] Wgt_6_502;input [WEIGHT_SIZE-1:0] Wgt_6_503;input [WEIGHT_SIZE-1:0] Wgt_6_504;input [WEIGHT_SIZE-1:0] Wgt_6_505;input [WEIGHT_SIZE-1:0] Wgt_6_506;input [WEIGHT_SIZE-1:0] Wgt_6_507;input [WEIGHT_SIZE-1:0] Wgt_6_508;input [WEIGHT_SIZE-1:0] Wgt_6_509;input [WEIGHT_SIZE-1:0] Wgt_6_510;input [WEIGHT_SIZE-1:0] Wgt_6_511;input [WEIGHT_SIZE-1:0] Wgt_6_512;input [WEIGHT_SIZE-1:0] Wgt_6_513;input [WEIGHT_SIZE-1:0] Wgt_6_514;input [WEIGHT_SIZE-1:0] Wgt_6_515;input [WEIGHT_SIZE-1:0] Wgt_6_516;input [WEIGHT_SIZE-1:0] Wgt_6_517;input [WEIGHT_SIZE-1:0] Wgt_6_518;input [WEIGHT_SIZE-1:0] Wgt_6_519;input [WEIGHT_SIZE-1:0] Wgt_6_520;input [WEIGHT_SIZE-1:0] Wgt_6_521;input [WEIGHT_SIZE-1:0] Wgt_6_522;input [WEIGHT_SIZE-1:0] Wgt_6_523;input [WEIGHT_SIZE-1:0] Wgt_6_524;input [WEIGHT_SIZE-1:0] Wgt_6_525;input [WEIGHT_SIZE-1:0] Wgt_6_526;input [WEIGHT_SIZE-1:0] Wgt_6_527;input [WEIGHT_SIZE-1:0] Wgt_6_528;input [WEIGHT_SIZE-1:0] Wgt_6_529;input [WEIGHT_SIZE-1:0] Wgt_6_530;input [WEIGHT_SIZE-1:0] Wgt_6_531;input [WEIGHT_SIZE-1:0] Wgt_6_532;input [WEIGHT_SIZE-1:0] Wgt_6_533;input [WEIGHT_SIZE-1:0] Wgt_6_534;input [WEIGHT_SIZE-1:0] Wgt_6_535;input [WEIGHT_SIZE-1:0] Wgt_6_536;input [WEIGHT_SIZE-1:0] Wgt_6_537;input [WEIGHT_SIZE-1:0] Wgt_6_538;input [WEIGHT_SIZE-1:0] Wgt_6_539;input [WEIGHT_SIZE-1:0] Wgt_6_540;input [WEIGHT_SIZE-1:0] Wgt_6_541;input [WEIGHT_SIZE-1:0] Wgt_6_542;input [WEIGHT_SIZE-1:0] Wgt_6_543;input [WEIGHT_SIZE-1:0] Wgt_6_544;input [WEIGHT_SIZE-1:0] Wgt_6_545;input [WEIGHT_SIZE-1:0] Wgt_6_546;input [WEIGHT_SIZE-1:0] Wgt_6_547;input [WEIGHT_SIZE-1:0] Wgt_6_548;input [WEIGHT_SIZE-1:0] Wgt_6_549;input [WEIGHT_SIZE-1:0] Wgt_6_550;input [WEIGHT_SIZE-1:0] Wgt_6_551;input [WEIGHT_SIZE-1:0] Wgt_6_552;input [WEIGHT_SIZE-1:0] Wgt_6_553;input [WEIGHT_SIZE-1:0] Wgt_6_554;input [WEIGHT_SIZE-1:0] Wgt_6_555;input [WEIGHT_SIZE-1:0] Wgt_6_556;input [WEIGHT_SIZE-1:0] Wgt_6_557;input [WEIGHT_SIZE-1:0] Wgt_6_558;input [WEIGHT_SIZE-1:0] Wgt_6_559;input [WEIGHT_SIZE-1:0] Wgt_6_560;input [WEIGHT_SIZE-1:0] Wgt_6_561;input [WEIGHT_SIZE-1:0] Wgt_6_562;input [WEIGHT_SIZE-1:0] Wgt_6_563;input [WEIGHT_SIZE-1:0] Wgt_6_564;input [WEIGHT_SIZE-1:0] Wgt_6_565;input [WEIGHT_SIZE-1:0] Wgt_6_566;input [WEIGHT_SIZE-1:0] Wgt_6_567;input [WEIGHT_SIZE-1:0] Wgt_6_568;input [WEIGHT_SIZE-1:0] Wgt_6_569;input [WEIGHT_SIZE-1:0] Wgt_6_570;input [WEIGHT_SIZE-1:0] Wgt_6_571;input [WEIGHT_SIZE-1:0] Wgt_6_572;input [WEIGHT_SIZE-1:0] Wgt_6_573;input [WEIGHT_SIZE-1:0] Wgt_6_574;input [WEIGHT_SIZE-1:0] Wgt_6_575;input [WEIGHT_SIZE-1:0] Wgt_6_576;input [WEIGHT_SIZE-1:0] Wgt_6_577;input [WEIGHT_SIZE-1:0] Wgt_6_578;input [WEIGHT_SIZE-1:0] Wgt_6_579;input [WEIGHT_SIZE-1:0] Wgt_6_580;input [WEIGHT_SIZE-1:0] Wgt_6_581;input [WEIGHT_SIZE-1:0] Wgt_6_582;input [WEIGHT_SIZE-1:0] Wgt_6_583;input [WEIGHT_SIZE-1:0] Wgt_6_584;input [WEIGHT_SIZE-1:0] Wgt_6_585;input [WEIGHT_SIZE-1:0] Wgt_6_586;input [WEIGHT_SIZE-1:0] Wgt_6_587;input [WEIGHT_SIZE-1:0] Wgt_6_588;input [WEIGHT_SIZE-1:0] Wgt_6_589;input [WEIGHT_SIZE-1:0] Wgt_6_590;input [WEIGHT_SIZE-1:0] Wgt_6_591;input [WEIGHT_SIZE-1:0] Wgt_6_592;input [WEIGHT_SIZE-1:0] Wgt_6_593;input [WEIGHT_SIZE-1:0] Wgt_6_594;input [WEIGHT_SIZE-1:0] Wgt_6_595;input [WEIGHT_SIZE-1:0] Wgt_6_596;input [WEIGHT_SIZE-1:0] Wgt_6_597;input [WEIGHT_SIZE-1:0] Wgt_6_598;input [WEIGHT_SIZE-1:0] Wgt_6_599;input [WEIGHT_SIZE-1:0] Wgt_6_600;input [WEIGHT_SIZE-1:0] Wgt_6_601;input [WEIGHT_SIZE-1:0] Wgt_6_602;input [WEIGHT_SIZE-1:0] Wgt_6_603;input [WEIGHT_SIZE-1:0] Wgt_6_604;input [WEIGHT_SIZE-1:0] Wgt_6_605;input [WEIGHT_SIZE-1:0] Wgt_6_606;input [WEIGHT_SIZE-1:0] Wgt_6_607;input [WEIGHT_SIZE-1:0] Wgt_6_608;input [WEIGHT_SIZE-1:0] Wgt_6_609;input [WEIGHT_SIZE-1:0] Wgt_6_610;input [WEIGHT_SIZE-1:0] Wgt_6_611;input [WEIGHT_SIZE-1:0] Wgt_6_612;input [WEIGHT_SIZE-1:0] Wgt_6_613;input [WEIGHT_SIZE-1:0] Wgt_6_614;input [WEIGHT_SIZE-1:0] Wgt_6_615;input [WEIGHT_SIZE-1:0] Wgt_6_616;input [WEIGHT_SIZE-1:0] Wgt_6_617;input [WEIGHT_SIZE-1:0] Wgt_6_618;input [WEIGHT_SIZE-1:0] Wgt_6_619;input [WEIGHT_SIZE-1:0] Wgt_6_620;input [WEIGHT_SIZE-1:0] Wgt_6_621;input [WEIGHT_SIZE-1:0] Wgt_6_622;input [WEIGHT_SIZE-1:0] Wgt_6_623;input [WEIGHT_SIZE-1:0] Wgt_6_624;input [WEIGHT_SIZE-1:0] Wgt_6_625;input [WEIGHT_SIZE-1:0] Wgt_6_626;input [WEIGHT_SIZE-1:0] Wgt_6_627;input [WEIGHT_SIZE-1:0] Wgt_6_628;input [WEIGHT_SIZE-1:0] Wgt_6_629;input [WEIGHT_SIZE-1:0] Wgt_6_630;input [WEIGHT_SIZE-1:0] Wgt_6_631;input [WEIGHT_SIZE-1:0] Wgt_6_632;input [WEIGHT_SIZE-1:0] Wgt_6_633;input [WEIGHT_SIZE-1:0] Wgt_6_634;input [WEIGHT_SIZE-1:0] Wgt_6_635;input [WEIGHT_SIZE-1:0] Wgt_6_636;input [WEIGHT_SIZE-1:0] Wgt_6_637;input [WEIGHT_SIZE-1:0] Wgt_6_638;input [WEIGHT_SIZE-1:0] Wgt_6_639;input [WEIGHT_SIZE-1:0] Wgt_6_640;input [WEIGHT_SIZE-1:0] Wgt_6_641;input [WEIGHT_SIZE-1:0] Wgt_6_642;input [WEIGHT_SIZE-1:0] Wgt_6_643;input [WEIGHT_SIZE-1:0] Wgt_6_644;input [WEIGHT_SIZE-1:0] Wgt_6_645;input [WEIGHT_SIZE-1:0] Wgt_6_646;input [WEIGHT_SIZE-1:0] Wgt_6_647;input [WEIGHT_SIZE-1:0] Wgt_6_648;input [WEIGHT_SIZE-1:0] Wgt_6_649;input [WEIGHT_SIZE-1:0] Wgt_6_650;input [WEIGHT_SIZE-1:0] Wgt_6_651;input [WEIGHT_SIZE-1:0] Wgt_6_652;input [WEIGHT_SIZE-1:0] Wgt_6_653;input [WEIGHT_SIZE-1:0] Wgt_6_654;input [WEIGHT_SIZE-1:0] Wgt_6_655;input [WEIGHT_SIZE-1:0] Wgt_6_656;input [WEIGHT_SIZE-1:0] Wgt_6_657;input [WEIGHT_SIZE-1:0] Wgt_6_658;input [WEIGHT_SIZE-1:0] Wgt_6_659;input [WEIGHT_SIZE-1:0] Wgt_6_660;input [WEIGHT_SIZE-1:0] Wgt_6_661;input [WEIGHT_SIZE-1:0] Wgt_6_662;input [WEIGHT_SIZE-1:0] Wgt_6_663;input [WEIGHT_SIZE-1:0] Wgt_6_664;input [WEIGHT_SIZE-1:0] Wgt_6_665;input [WEIGHT_SIZE-1:0] Wgt_6_666;input [WEIGHT_SIZE-1:0] Wgt_6_667;input [WEIGHT_SIZE-1:0] Wgt_6_668;input [WEIGHT_SIZE-1:0] Wgt_6_669;input [WEIGHT_SIZE-1:0] Wgt_6_670;input [WEIGHT_SIZE-1:0] Wgt_6_671;input [WEIGHT_SIZE-1:0] Wgt_6_672;input [WEIGHT_SIZE-1:0] Wgt_6_673;input [WEIGHT_SIZE-1:0] Wgt_6_674;input [WEIGHT_SIZE-1:0] Wgt_6_675;input [WEIGHT_SIZE-1:0] Wgt_6_676;input [WEIGHT_SIZE-1:0] Wgt_6_677;input [WEIGHT_SIZE-1:0] Wgt_6_678;input [WEIGHT_SIZE-1:0] Wgt_6_679;input [WEIGHT_SIZE-1:0] Wgt_6_680;input [WEIGHT_SIZE-1:0] Wgt_6_681;input [WEIGHT_SIZE-1:0] Wgt_6_682;input [WEIGHT_SIZE-1:0] Wgt_6_683;input [WEIGHT_SIZE-1:0] Wgt_6_684;input [WEIGHT_SIZE-1:0] Wgt_6_685;input [WEIGHT_SIZE-1:0] Wgt_6_686;input [WEIGHT_SIZE-1:0] Wgt_6_687;input [WEIGHT_SIZE-1:0] Wgt_6_688;input [WEIGHT_SIZE-1:0] Wgt_6_689;input [WEIGHT_SIZE-1:0] Wgt_6_690;input [WEIGHT_SIZE-1:0] Wgt_6_691;input [WEIGHT_SIZE-1:0] Wgt_6_692;input [WEIGHT_SIZE-1:0] Wgt_6_693;input [WEIGHT_SIZE-1:0] Wgt_6_694;input [WEIGHT_SIZE-1:0] Wgt_6_695;input [WEIGHT_SIZE-1:0] Wgt_6_696;input [WEIGHT_SIZE-1:0] Wgt_6_697;input [WEIGHT_SIZE-1:0] Wgt_6_698;input [WEIGHT_SIZE-1:0] Wgt_6_699;input [WEIGHT_SIZE-1:0] Wgt_6_700;input [WEIGHT_SIZE-1:0] Wgt_6_701;input [WEIGHT_SIZE-1:0] Wgt_6_702;input [WEIGHT_SIZE-1:0] Wgt_6_703;input [WEIGHT_SIZE-1:0] Wgt_6_704;input [WEIGHT_SIZE-1:0] Wgt_6_705;input [WEIGHT_SIZE-1:0] Wgt_6_706;input [WEIGHT_SIZE-1:0] Wgt_6_707;input [WEIGHT_SIZE-1:0] Wgt_6_708;input [WEIGHT_SIZE-1:0] Wgt_6_709;input [WEIGHT_SIZE-1:0] Wgt_6_710;input [WEIGHT_SIZE-1:0] Wgt_6_711;input [WEIGHT_SIZE-1:0] Wgt_6_712;input [WEIGHT_SIZE-1:0] Wgt_6_713;input [WEIGHT_SIZE-1:0] Wgt_6_714;input [WEIGHT_SIZE-1:0] Wgt_6_715;input [WEIGHT_SIZE-1:0] Wgt_6_716;input [WEIGHT_SIZE-1:0] Wgt_6_717;input [WEIGHT_SIZE-1:0] Wgt_6_718;input [WEIGHT_SIZE-1:0] Wgt_6_719;input [WEIGHT_SIZE-1:0] Wgt_6_720;input [WEIGHT_SIZE-1:0] Wgt_6_721;input [WEIGHT_SIZE-1:0] Wgt_6_722;input [WEIGHT_SIZE-1:0] Wgt_6_723;input [WEIGHT_SIZE-1:0] Wgt_6_724;input [WEIGHT_SIZE-1:0] Wgt_6_725;input [WEIGHT_SIZE-1:0] Wgt_6_726;input [WEIGHT_SIZE-1:0] Wgt_6_727;input [WEIGHT_SIZE-1:0] Wgt_6_728;input [WEIGHT_SIZE-1:0] Wgt_6_729;input [WEIGHT_SIZE-1:0] Wgt_6_730;input [WEIGHT_SIZE-1:0] Wgt_6_731;input [WEIGHT_SIZE-1:0] Wgt_6_732;input [WEIGHT_SIZE-1:0] Wgt_6_733;input [WEIGHT_SIZE-1:0] Wgt_6_734;input [WEIGHT_SIZE-1:0] Wgt_6_735;input [WEIGHT_SIZE-1:0] Wgt_6_736;input [WEIGHT_SIZE-1:0] Wgt_6_737;input [WEIGHT_SIZE-1:0] Wgt_6_738;input [WEIGHT_SIZE-1:0] Wgt_6_739;input [WEIGHT_SIZE-1:0] Wgt_6_740;input [WEIGHT_SIZE-1:0] Wgt_6_741;input [WEIGHT_SIZE-1:0] Wgt_6_742;input [WEIGHT_SIZE-1:0] Wgt_6_743;input [WEIGHT_SIZE-1:0] Wgt_6_744;input [WEIGHT_SIZE-1:0] Wgt_6_745;input [WEIGHT_SIZE-1:0] Wgt_6_746;input [WEIGHT_SIZE-1:0] Wgt_6_747;input [WEIGHT_SIZE-1:0] Wgt_6_748;input [WEIGHT_SIZE-1:0] Wgt_6_749;input [WEIGHT_SIZE-1:0] Wgt_6_750;input [WEIGHT_SIZE-1:0] Wgt_6_751;input [WEIGHT_SIZE-1:0] Wgt_6_752;input [WEIGHT_SIZE-1:0] Wgt_6_753;input [WEIGHT_SIZE-1:0] Wgt_6_754;input [WEIGHT_SIZE-1:0] Wgt_6_755;input [WEIGHT_SIZE-1:0] Wgt_6_756;input [WEIGHT_SIZE-1:0] Wgt_6_757;input [WEIGHT_SIZE-1:0] Wgt_6_758;input [WEIGHT_SIZE-1:0] Wgt_6_759;input [WEIGHT_SIZE-1:0] Wgt_6_760;input [WEIGHT_SIZE-1:0] Wgt_6_761;input [WEIGHT_SIZE-1:0] Wgt_6_762;input [WEIGHT_SIZE-1:0] Wgt_6_763;input [WEIGHT_SIZE-1:0] Wgt_6_764;input [WEIGHT_SIZE-1:0] Wgt_6_765;input [WEIGHT_SIZE-1:0] Wgt_6_766;input [WEIGHT_SIZE-1:0] Wgt_6_767;input [WEIGHT_SIZE-1:0] Wgt_6_768;input [WEIGHT_SIZE-1:0] Wgt_6_769;input [WEIGHT_SIZE-1:0] Wgt_6_770;input [WEIGHT_SIZE-1:0] Wgt_6_771;input [WEIGHT_SIZE-1:0] Wgt_6_772;input [WEIGHT_SIZE-1:0] Wgt_6_773;input [WEIGHT_SIZE-1:0] Wgt_6_774;input [WEIGHT_SIZE-1:0] Wgt_6_775;input [WEIGHT_SIZE-1:0] Wgt_6_776;input [WEIGHT_SIZE-1:0] Wgt_6_777;input [WEIGHT_SIZE-1:0] Wgt_6_778;input [WEIGHT_SIZE-1:0] Wgt_6_779;input [WEIGHT_SIZE-1:0] Wgt_6_780;input [WEIGHT_SIZE-1:0] Wgt_6_781;input [WEIGHT_SIZE-1:0] Wgt_6_782;input [WEIGHT_SIZE-1:0] Wgt_6_783;input [WEIGHT_SIZE-1:0] Wgt_6_784;input [WEIGHT_SIZE-1:0] Wgt_7_0;input [WEIGHT_SIZE-1:0] Wgt_7_1;input [WEIGHT_SIZE-1:0] Wgt_7_2;input [WEIGHT_SIZE-1:0] Wgt_7_3;input [WEIGHT_SIZE-1:0] Wgt_7_4;input [WEIGHT_SIZE-1:0] Wgt_7_5;input [WEIGHT_SIZE-1:0] Wgt_7_6;input [WEIGHT_SIZE-1:0] Wgt_7_7;input [WEIGHT_SIZE-1:0] Wgt_7_8;input [WEIGHT_SIZE-1:0] Wgt_7_9;input [WEIGHT_SIZE-1:0] Wgt_7_10;input [WEIGHT_SIZE-1:0] Wgt_7_11;input [WEIGHT_SIZE-1:0] Wgt_7_12;input [WEIGHT_SIZE-1:0] Wgt_7_13;input [WEIGHT_SIZE-1:0] Wgt_7_14;input [WEIGHT_SIZE-1:0] Wgt_7_15;input [WEIGHT_SIZE-1:0] Wgt_7_16;input [WEIGHT_SIZE-1:0] Wgt_7_17;input [WEIGHT_SIZE-1:0] Wgt_7_18;input [WEIGHT_SIZE-1:0] Wgt_7_19;input [WEIGHT_SIZE-1:0] Wgt_7_20;input [WEIGHT_SIZE-1:0] Wgt_7_21;input [WEIGHT_SIZE-1:0] Wgt_7_22;input [WEIGHT_SIZE-1:0] Wgt_7_23;input [WEIGHT_SIZE-1:0] Wgt_7_24;input [WEIGHT_SIZE-1:0] Wgt_7_25;input [WEIGHT_SIZE-1:0] Wgt_7_26;input [WEIGHT_SIZE-1:0] Wgt_7_27;input [WEIGHT_SIZE-1:0] Wgt_7_28;input [WEIGHT_SIZE-1:0] Wgt_7_29;input [WEIGHT_SIZE-1:0] Wgt_7_30;input [WEIGHT_SIZE-1:0] Wgt_7_31;input [WEIGHT_SIZE-1:0] Wgt_7_32;input [WEIGHT_SIZE-1:0] Wgt_7_33;input [WEIGHT_SIZE-1:0] Wgt_7_34;input [WEIGHT_SIZE-1:0] Wgt_7_35;input [WEIGHT_SIZE-1:0] Wgt_7_36;input [WEIGHT_SIZE-1:0] Wgt_7_37;input [WEIGHT_SIZE-1:0] Wgt_7_38;input [WEIGHT_SIZE-1:0] Wgt_7_39;input [WEIGHT_SIZE-1:0] Wgt_7_40;input [WEIGHT_SIZE-1:0] Wgt_7_41;input [WEIGHT_SIZE-1:0] Wgt_7_42;input [WEIGHT_SIZE-1:0] Wgt_7_43;input [WEIGHT_SIZE-1:0] Wgt_7_44;input [WEIGHT_SIZE-1:0] Wgt_7_45;input [WEIGHT_SIZE-1:0] Wgt_7_46;input [WEIGHT_SIZE-1:0] Wgt_7_47;input [WEIGHT_SIZE-1:0] Wgt_7_48;input [WEIGHT_SIZE-1:0] Wgt_7_49;input [WEIGHT_SIZE-1:0] Wgt_7_50;input [WEIGHT_SIZE-1:0] Wgt_7_51;input [WEIGHT_SIZE-1:0] Wgt_7_52;input [WEIGHT_SIZE-1:0] Wgt_7_53;input [WEIGHT_SIZE-1:0] Wgt_7_54;input [WEIGHT_SIZE-1:0] Wgt_7_55;input [WEIGHT_SIZE-1:0] Wgt_7_56;input [WEIGHT_SIZE-1:0] Wgt_7_57;input [WEIGHT_SIZE-1:0] Wgt_7_58;input [WEIGHT_SIZE-1:0] Wgt_7_59;input [WEIGHT_SIZE-1:0] Wgt_7_60;input [WEIGHT_SIZE-1:0] Wgt_7_61;input [WEIGHT_SIZE-1:0] Wgt_7_62;input [WEIGHT_SIZE-1:0] Wgt_7_63;input [WEIGHT_SIZE-1:0] Wgt_7_64;input [WEIGHT_SIZE-1:0] Wgt_7_65;input [WEIGHT_SIZE-1:0] Wgt_7_66;input [WEIGHT_SIZE-1:0] Wgt_7_67;input [WEIGHT_SIZE-1:0] Wgt_7_68;input [WEIGHT_SIZE-1:0] Wgt_7_69;input [WEIGHT_SIZE-1:0] Wgt_7_70;input [WEIGHT_SIZE-1:0] Wgt_7_71;input [WEIGHT_SIZE-1:0] Wgt_7_72;input [WEIGHT_SIZE-1:0] Wgt_7_73;input [WEIGHT_SIZE-1:0] Wgt_7_74;input [WEIGHT_SIZE-1:0] Wgt_7_75;input [WEIGHT_SIZE-1:0] Wgt_7_76;input [WEIGHT_SIZE-1:0] Wgt_7_77;input [WEIGHT_SIZE-1:0] Wgt_7_78;input [WEIGHT_SIZE-1:0] Wgt_7_79;input [WEIGHT_SIZE-1:0] Wgt_7_80;input [WEIGHT_SIZE-1:0] Wgt_7_81;input [WEIGHT_SIZE-1:0] Wgt_7_82;input [WEIGHT_SIZE-1:0] Wgt_7_83;input [WEIGHT_SIZE-1:0] Wgt_7_84;input [WEIGHT_SIZE-1:0] Wgt_7_85;input [WEIGHT_SIZE-1:0] Wgt_7_86;input [WEIGHT_SIZE-1:0] Wgt_7_87;input [WEIGHT_SIZE-1:0] Wgt_7_88;input [WEIGHT_SIZE-1:0] Wgt_7_89;input [WEIGHT_SIZE-1:0] Wgt_7_90;input [WEIGHT_SIZE-1:0] Wgt_7_91;input [WEIGHT_SIZE-1:0] Wgt_7_92;input [WEIGHT_SIZE-1:0] Wgt_7_93;input [WEIGHT_SIZE-1:0] Wgt_7_94;input [WEIGHT_SIZE-1:0] Wgt_7_95;input [WEIGHT_SIZE-1:0] Wgt_7_96;input [WEIGHT_SIZE-1:0] Wgt_7_97;input [WEIGHT_SIZE-1:0] Wgt_7_98;input [WEIGHT_SIZE-1:0] Wgt_7_99;input [WEIGHT_SIZE-1:0] Wgt_7_100;input [WEIGHT_SIZE-1:0] Wgt_7_101;input [WEIGHT_SIZE-1:0] Wgt_7_102;input [WEIGHT_SIZE-1:0] Wgt_7_103;input [WEIGHT_SIZE-1:0] Wgt_7_104;input [WEIGHT_SIZE-1:0] Wgt_7_105;input [WEIGHT_SIZE-1:0] Wgt_7_106;input [WEIGHT_SIZE-1:0] Wgt_7_107;input [WEIGHT_SIZE-1:0] Wgt_7_108;input [WEIGHT_SIZE-1:0] Wgt_7_109;input [WEIGHT_SIZE-1:0] Wgt_7_110;input [WEIGHT_SIZE-1:0] Wgt_7_111;input [WEIGHT_SIZE-1:0] Wgt_7_112;input [WEIGHT_SIZE-1:0] Wgt_7_113;input [WEIGHT_SIZE-1:0] Wgt_7_114;input [WEIGHT_SIZE-1:0] Wgt_7_115;input [WEIGHT_SIZE-1:0] Wgt_7_116;input [WEIGHT_SIZE-1:0] Wgt_7_117;input [WEIGHT_SIZE-1:0] Wgt_7_118;input [WEIGHT_SIZE-1:0] Wgt_7_119;input [WEIGHT_SIZE-1:0] Wgt_7_120;input [WEIGHT_SIZE-1:0] Wgt_7_121;input [WEIGHT_SIZE-1:0] Wgt_7_122;input [WEIGHT_SIZE-1:0] Wgt_7_123;input [WEIGHT_SIZE-1:0] Wgt_7_124;input [WEIGHT_SIZE-1:0] Wgt_7_125;input [WEIGHT_SIZE-1:0] Wgt_7_126;input [WEIGHT_SIZE-1:0] Wgt_7_127;input [WEIGHT_SIZE-1:0] Wgt_7_128;input [WEIGHT_SIZE-1:0] Wgt_7_129;input [WEIGHT_SIZE-1:0] Wgt_7_130;input [WEIGHT_SIZE-1:0] Wgt_7_131;input [WEIGHT_SIZE-1:0] Wgt_7_132;input [WEIGHT_SIZE-1:0] Wgt_7_133;input [WEIGHT_SIZE-1:0] Wgt_7_134;input [WEIGHT_SIZE-1:0] Wgt_7_135;input [WEIGHT_SIZE-1:0] Wgt_7_136;input [WEIGHT_SIZE-1:0] Wgt_7_137;input [WEIGHT_SIZE-1:0] Wgt_7_138;input [WEIGHT_SIZE-1:0] Wgt_7_139;input [WEIGHT_SIZE-1:0] Wgt_7_140;input [WEIGHT_SIZE-1:0] Wgt_7_141;input [WEIGHT_SIZE-1:0] Wgt_7_142;input [WEIGHT_SIZE-1:0] Wgt_7_143;input [WEIGHT_SIZE-1:0] Wgt_7_144;input [WEIGHT_SIZE-1:0] Wgt_7_145;input [WEIGHT_SIZE-1:0] Wgt_7_146;input [WEIGHT_SIZE-1:0] Wgt_7_147;input [WEIGHT_SIZE-1:0] Wgt_7_148;input [WEIGHT_SIZE-1:0] Wgt_7_149;input [WEIGHT_SIZE-1:0] Wgt_7_150;input [WEIGHT_SIZE-1:0] Wgt_7_151;input [WEIGHT_SIZE-1:0] Wgt_7_152;input [WEIGHT_SIZE-1:0] Wgt_7_153;input [WEIGHT_SIZE-1:0] Wgt_7_154;input [WEIGHT_SIZE-1:0] Wgt_7_155;input [WEIGHT_SIZE-1:0] Wgt_7_156;input [WEIGHT_SIZE-1:0] Wgt_7_157;input [WEIGHT_SIZE-1:0] Wgt_7_158;input [WEIGHT_SIZE-1:0] Wgt_7_159;input [WEIGHT_SIZE-1:0] Wgt_7_160;input [WEIGHT_SIZE-1:0] Wgt_7_161;input [WEIGHT_SIZE-1:0] Wgt_7_162;input [WEIGHT_SIZE-1:0] Wgt_7_163;input [WEIGHT_SIZE-1:0] Wgt_7_164;input [WEIGHT_SIZE-1:0] Wgt_7_165;input [WEIGHT_SIZE-1:0] Wgt_7_166;input [WEIGHT_SIZE-1:0] Wgt_7_167;input [WEIGHT_SIZE-1:0] Wgt_7_168;input [WEIGHT_SIZE-1:0] Wgt_7_169;input [WEIGHT_SIZE-1:0] Wgt_7_170;input [WEIGHT_SIZE-1:0] Wgt_7_171;input [WEIGHT_SIZE-1:0] Wgt_7_172;input [WEIGHT_SIZE-1:0] Wgt_7_173;input [WEIGHT_SIZE-1:0] Wgt_7_174;input [WEIGHT_SIZE-1:0] Wgt_7_175;input [WEIGHT_SIZE-1:0] Wgt_7_176;input [WEIGHT_SIZE-1:0] Wgt_7_177;input [WEIGHT_SIZE-1:0] Wgt_7_178;input [WEIGHT_SIZE-1:0] Wgt_7_179;input [WEIGHT_SIZE-1:0] Wgt_7_180;input [WEIGHT_SIZE-1:0] Wgt_7_181;input [WEIGHT_SIZE-1:0] Wgt_7_182;input [WEIGHT_SIZE-1:0] Wgt_7_183;input [WEIGHT_SIZE-1:0] Wgt_7_184;input [WEIGHT_SIZE-1:0] Wgt_7_185;input [WEIGHT_SIZE-1:0] Wgt_7_186;input [WEIGHT_SIZE-1:0] Wgt_7_187;input [WEIGHT_SIZE-1:0] Wgt_7_188;input [WEIGHT_SIZE-1:0] Wgt_7_189;input [WEIGHT_SIZE-1:0] Wgt_7_190;input [WEIGHT_SIZE-1:0] Wgt_7_191;input [WEIGHT_SIZE-1:0] Wgt_7_192;input [WEIGHT_SIZE-1:0] Wgt_7_193;input [WEIGHT_SIZE-1:0] Wgt_7_194;input [WEIGHT_SIZE-1:0] Wgt_7_195;input [WEIGHT_SIZE-1:0] Wgt_7_196;input [WEIGHT_SIZE-1:0] Wgt_7_197;input [WEIGHT_SIZE-1:0] Wgt_7_198;input [WEIGHT_SIZE-1:0] Wgt_7_199;input [WEIGHT_SIZE-1:0] Wgt_7_200;input [WEIGHT_SIZE-1:0] Wgt_7_201;input [WEIGHT_SIZE-1:0] Wgt_7_202;input [WEIGHT_SIZE-1:0] Wgt_7_203;input [WEIGHT_SIZE-1:0] Wgt_7_204;input [WEIGHT_SIZE-1:0] Wgt_7_205;input [WEIGHT_SIZE-1:0] Wgt_7_206;input [WEIGHT_SIZE-1:0] Wgt_7_207;input [WEIGHT_SIZE-1:0] Wgt_7_208;input [WEIGHT_SIZE-1:0] Wgt_7_209;input [WEIGHT_SIZE-1:0] Wgt_7_210;input [WEIGHT_SIZE-1:0] Wgt_7_211;input [WEIGHT_SIZE-1:0] Wgt_7_212;input [WEIGHT_SIZE-1:0] Wgt_7_213;input [WEIGHT_SIZE-1:0] Wgt_7_214;input [WEIGHT_SIZE-1:0] Wgt_7_215;input [WEIGHT_SIZE-1:0] Wgt_7_216;input [WEIGHT_SIZE-1:0] Wgt_7_217;input [WEIGHT_SIZE-1:0] Wgt_7_218;input [WEIGHT_SIZE-1:0] Wgt_7_219;input [WEIGHT_SIZE-1:0] Wgt_7_220;input [WEIGHT_SIZE-1:0] Wgt_7_221;input [WEIGHT_SIZE-1:0] Wgt_7_222;input [WEIGHT_SIZE-1:0] Wgt_7_223;input [WEIGHT_SIZE-1:0] Wgt_7_224;input [WEIGHT_SIZE-1:0] Wgt_7_225;input [WEIGHT_SIZE-1:0] Wgt_7_226;input [WEIGHT_SIZE-1:0] Wgt_7_227;input [WEIGHT_SIZE-1:0] Wgt_7_228;input [WEIGHT_SIZE-1:0] Wgt_7_229;input [WEIGHT_SIZE-1:0] Wgt_7_230;input [WEIGHT_SIZE-1:0] Wgt_7_231;input [WEIGHT_SIZE-1:0] Wgt_7_232;input [WEIGHT_SIZE-1:0] Wgt_7_233;input [WEIGHT_SIZE-1:0] Wgt_7_234;input [WEIGHT_SIZE-1:0] Wgt_7_235;input [WEIGHT_SIZE-1:0] Wgt_7_236;input [WEIGHT_SIZE-1:0] Wgt_7_237;input [WEIGHT_SIZE-1:0] Wgt_7_238;input [WEIGHT_SIZE-1:0] Wgt_7_239;input [WEIGHT_SIZE-1:0] Wgt_7_240;input [WEIGHT_SIZE-1:0] Wgt_7_241;input [WEIGHT_SIZE-1:0] Wgt_7_242;input [WEIGHT_SIZE-1:0] Wgt_7_243;input [WEIGHT_SIZE-1:0] Wgt_7_244;input [WEIGHT_SIZE-1:0] Wgt_7_245;input [WEIGHT_SIZE-1:0] Wgt_7_246;input [WEIGHT_SIZE-1:0] Wgt_7_247;input [WEIGHT_SIZE-1:0] Wgt_7_248;input [WEIGHT_SIZE-1:0] Wgt_7_249;input [WEIGHT_SIZE-1:0] Wgt_7_250;input [WEIGHT_SIZE-1:0] Wgt_7_251;input [WEIGHT_SIZE-1:0] Wgt_7_252;input [WEIGHT_SIZE-1:0] Wgt_7_253;input [WEIGHT_SIZE-1:0] Wgt_7_254;input [WEIGHT_SIZE-1:0] Wgt_7_255;input [WEIGHT_SIZE-1:0] Wgt_7_256;input [WEIGHT_SIZE-1:0] Wgt_7_257;input [WEIGHT_SIZE-1:0] Wgt_7_258;input [WEIGHT_SIZE-1:0] Wgt_7_259;input [WEIGHT_SIZE-1:0] Wgt_7_260;input [WEIGHT_SIZE-1:0] Wgt_7_261;input [WEIGHT_SIZE-1:0] Wgt_7_262;input [WEIGHT_SIZE-1:0] Wgt_7_263;input [WEIGHT_SIZE-1:0] Wgt_7_264;input [WEIGHT_SIZE-1:0] Wgt_7_265;input [WEIGHT_SIZE-1:0] Wgt_7_266;input [WEIGHT_SIZE-1:0] Wgt_7_267;input [WEIGHT_SIZE-1:0] Wgt_7_268;input [WEIGHT_SIZE-1:0] Wgt_7_269;input [WEIGHT_SIZE-1:0] Wgt_7_270;input [WEIGHT_SIZE-1:0] Wgt_7_271;input [WEIGHT_SIZE-1:0] Wgt_7_272;input [WEIGHT_SIZE-1:0] Wgt_7_273;input [WEIGHT_SIZE-1:0] Wgt_7_274;input [WEIGHT_SIZE-1:0] Wgt_7_275;input [WEIGHT_SIZE-1:0] Wgt_7_276;input [WEIGHT_SIZE-1:0] Wgt_7_277;input [WEIGHT_SIZE-1:0] Wgt_7_278;input [WEIGHT_SIZE-1:0] Wgt_7_279;input [WEIGHT_SIZE-1:0] Wgt_7_280;input [WEIGHT_SIZE-1:0] Wgt_7_281;input [WEIGHT_SIZE-1:0] Wgt_7_282;input [WEIGHT_SIZE-1:0] Wgt_7_283;input [WEIGHT_SIZE-1:0] Wgt_7_284;input [WEIGHT_SIZE-1:0] Wgt_7_285;input [WEIGHT_SIZE-1:0] Wgt_7_286;input [WEIGHT_SIZE-1:0] Wgt_7_287;input [WEIGHT_SIZE-1:0] Wgt_7_288;input [WEIGHT_SIZE-1:0] Wgt_7_289;input [WEIGHT_SIZE-1:0] Wgt_7_290;input [WEIGHT_SIZE-1:0] Wgt_7_291;input [WEIGHT_SIZE-1:0] Wgt_7_292;input [WEIGHT_SIZE-1:0] Wgt_7_293;input [WEIGHT_SIZE-1:0] Wgt_7_294;input [WEIGHT_SIZE-1:0] Wgt_7_295;input [WEIGHT_SIZE-1:0] Wgt_7_296;input [WEIGHT_SIZE-1:0] Wgt_7_297;input [WEIGHT_SIZE-1:0] Wgt_7_298;input [WEIGHT_SIZE-1:0] Wgt_7_299;input [WEIGHT_SIZE-1:0] Wgt_7_300;input [WEIGHT_SIZE-1:0] Wgt_7_301;input [WEIGHT_SIZE-1:0] Wgt_7_302;input [WEIGHT_SIZE-1:0] Wgt_7_303;input [WEIGHT_SIZE-1:0] Wgt_7_304;input [WEIGHT_SIZE-1:0] Wgt_7_305;input [WEIGHT_SIZE-1:0] Wgt_7_306;input [WEIGHT_SIZE-1:0] Wgt_7_307;input [WEIGHT_SIZE-1:0] Wgt_7_308;input [WEIGHT_SIZE-1:0] Wgt_7_309;input [WEIGHT_SIZE-1:0] Wgt_7_310;input [WEIGHT_SIZE-1:0] Wgt_7_311;input [WEIGHT_SIZE-1:0] Wgt_7_312;input [WEIGHT_SIZE-1:0] Wgt_7_313;input [WEIGHT_SIZE-1:0] Wgt_7_314;input [WEIGHT_SIZE-1:0] Wgt_7_315;input [WEIGHT_SIZE-1:0] Wgt_7_316;input [WEIGHT_SIZE-1:0] Wgt_7_317;input [WEIGHT_SIZE-1:0] Wgt_7_318;input [WEIGHT_SIZE-1:0] Wgt_7_319;input [WEIGHT_SIZE-1:0] Wgt_7_320;input [WEIGHT_SIZE-1:0] Wgt_7_321;input [WEIGHT_SIZE-1:0] Wgt_7_322;input [WEIGHT_SIZE-1:0] Wgt_7_323;input [WEIGHT_SIZE-1:0] Wgt_7_324;input [WEIGHT_SIZE-1:0] Wgt_7_325;input [WEIGHT_SIZE-1:0] Wgt_7_326;input [WEIGHT_SIZE-1:0] Wgt_7_327;input [WEIGHT_SIZE-1:0] Wgt_7_328;input [WEIGHT_SIZE-1:0] Wgt_7_329;input [WEIGHT_SIZE-1:0] Wgt_7_330;input [WEIGHT_SIZE-1:0] Wgt_7_331;input [WEIGHT_SIZE-1:0] Wgt_7_332;input [WEIGHT_SIZE-1:0] Wgt_7_333;input [WEIGHT_SIZE-1:0] Wgt_7_334;input [WEIGHT_SIZE-1:0] Wgt_7_335;input [WEIGHT_SIZE-1:0] Wgt_7_336;input [WEIGHT_SIZE-1:0] Wgt_7_337;input [WEIGHT_SIZE-1:0] Wgt_7_338;input [WEIGHT_SIZE-1:0] Wgt_7_339;input [WEIGHT_SIZE-1:0] Wgt_7_340;input [WEIGHT_SIZE-1:0] Wgt_7_341;input [WEIGHT_SIZE-1:0] Wgt_7_342;input [WEIGHT_SIZE-1:0] Wgt_7_343;input [WEIGHT_SIZE-1:0] Wgt_7_344;input [WEIGHT_SIZE-1:0] Wgt_7_345;input [WEIGHT_SIZE-1:0] Wgt_7_346;input [WEIGHT_SIZE-1:0] Wgt_7_347;input [WEIGHT_SIZE-1:0] Wgt_7_348;input [WEIGHT_SIZE-1:0] Wgt_7_349;input [WEIGHT_SIZE-1:0] Wgt_7_350;input [WEIGHT_SIZE-1:0] Wgt_7_351;input [WEIGHT_SIZE-1:0] Wgt_7_352;input [WEIGHT_SIZE-1:0] Wgt_7_353;input [WEIGHT_SIZE-1:0] Wgt_7_354;input [WEIGHT_SIZE-1:0] Wgt_7_355;input [WEIGHT_SIZE-1:0] Wgt_7_356;input [WEIGHT_SIZE-1:0] Wgt_7_357;input [WEIGHT_SIZE-1:0] Wgt_7_358;input [WEIGHT_SIZE-1:0] Wgt_7_359;input [WEIGHT_SIZE-1:0] Wgt_7_360;input [WEIGHT_SIZE-1:0] Wgt_7_361;input [WEIGHT_SIZE-1:0] Wgt_7_362;input [WEIGHT_SIZE-1:0] Wgt_7_363;input [WEIGHT_SIZE-1:0] Wgt_7_364;input [WEIGHT_SIZE-1:0] Wgt_7_365;input [WEIGHT_SIZE-1:0] Wgt_7_366;input [WEIGHT_SIZE-1:0] Wgt_7_367;input [WEIGHT_SIZE-1:0] Wgt_7_368;input [WEIGHT_SIZE-1:0] Wgt_7_369;input [WEIGHT_SIZE-1:0] Wgt_7_370;input [WEIGHT_SIZE-1:0] Wgt_7_371;input [WEIGHT_SIZE-1:0] Wgt_7_372;input [WEIGHT_SIZE-1:0] Wgt_7_373;input [WEIGHT_SIZE-1:0] Wgt_7_374;input [WEIGHT_SIZE-1:0] Wgt_7_375;input [WEIGHT_SIZE-1:0] Wgt_7_376;input [WEIGHT_SIZE-1:0] Wgt_7_377;input [WEIGHT_SIZE-1:0] Wgt_7_378;input [WEIGHT_SIZE-1:0] Wgt_7_379;input [WEIGHT_SIZE-1:0] Wgt_7_380;input [WEIGHT_SIZE-1:0] Wgt_7_381;input [WEIGHT_SIZE-1:0] Wgt_7_382;input [WEIGHT_SIZE-1:0] Wgt_7_383;input [WEIGHT_SIZE-1:0] Wgt_7_384;input [WEIGHT_SIZE-1:0] Wgt_7_385;input [WEIGHT_SIZE-1:0] Wgt_7_386;input [WEIGHT_SIZE-1:0] Wgt_7_387;input [WEIGHT_SIZE-1:0] Wgt_7_388;input [WEIGHT_SIZE-1:0] Wgt_7_389;input [WEIGHT_SIZE-1:0] Wgt_7_390;input [WEIGHT_SIZE-1:0] Wgt_7_391;input [WEIGHT_SIZE-1:0] Wgt_7_392;input [WEIGHT_SIZE-1:0] Wgt_7_393;input [WEIGHT_SIZE-1:0] Wgt_7_394;input [WEIGHT_SIZE-1:0] Wgt_7_395;input [WEIGHT_SIZE-1:0] Wgt_7_396;input [WEIGHT_SIZE-1:0] Wgt_7_397;input [WEIGHT_SIZE-1:0] Wgt_7_398;input [WEIGHT_SIZE-1:0] Wgt_7_399;input [WEIGHT_SIZE-1:0] Wgt_7_400;input [WEIGHT_SIZE-1:0] Wgt_7_401;input [WEIGHT_SIZE-1:0] Wgt_7_402;input [WEIGHT_SIZE-1:0] Wgt_7_403;input [WEIGHT_SIZE-1:0] Wgt_7_404;input [WEIGHT_SIZE-1:0] Wgt_7_405;input [WEIGHT_SIZE-1:0] Wgt_7_406;input [WEIGHT_SIZE-1:0] Wgt_7_407;input [WEIGHT_SIZE-1:0] Wgt_7_408;input [WEIGHT_SIZE-1:0] Wgt_7_409;input [WEIGHT_SIZE-1:0] Wgt_7_410;input [WEIGHT_SIZE-1:0] Wgt_7_411;input [WEIGHT_SIZE-1:0] Wgt_7_412;input [WEIGHT_SIZE-1:0] Wgt_7_413;input [WEIGHT_SIZE-1:0] Wgt_7_414;input [WEIGHT_SIZE-1:0] Wgt_7_415;input [WEIGHT_SIZE-1:0] Wgt_7_416;input [WEIGHT_SIZE-1:0] Wgt_7_417;input [WEIGHT_SIZE-1:0] Wgt_7_418;input [WEIGHT_SIZE-1:0] Wgt_7_419;input [WEIGHT_SIZE-1:0] Wgt_7_420;input [WEIGHT_SIZE-1:0] Wgt_7_421;input [WEIGHT_SIZE-1:0] Wgt_7_422;input [WEIGHT_SIZE-1:0] Wgt_7_423;input [WEIGHT_SIZE-1:0] Wgt_7_424;input [WEIGHT_SIZE-1:0] Wgt_7_425;input [WEIGHT_SIZE-1:0] Wgt_7_426;input [WEIGHT_SIZE-1:0] Wgt_7_427;input [WEIGHT_SIZE-1:0] Wgt_7_428;input [WEIGHT_SIZE-1:0] Wgt_7_429;input [WEIGHT_SIZE-1:0] Wgt_7_430;input [WEIGHT_SIZE-1:0] Wgt_7_431;input [WEIGHT_SIZE-1:0] Wgt_7_432;input [WEIGHT_SIZE-1:0] Wgt_7_433;input [WEIGHT_SIZE-1:0] Wgt_7_434;input [WEIGHT_SIZE-1:0] Wgt_7_435;input [WEIGHT_SIZE-1:0] Wgt_7_436;input [WEIGHT_SIZE-1:0] Wgt_7_437;input [WEIGHT_SIZE-1:0] Wgt_7_438;input [WEIGHT_SIZE-1:0] Wgt_7_439;input [WEIGHT_SIZE-1:0] Wgt_7_440;input [WEIGHT_SIZE-1:0] Wgt_7_441;input [WEIGHT_SIZE-1:0] Wgt_7_442;input [WEIGHT_SIZE-1:0] Wgt_7_443;input [WEIGHT_SIZE-1:0] Wgt_7_444;input [WEIGHT_SIZE-1:0] Wgt_7_445;input [WEIGHT_SIZE-1:0] Wgt_7_446;input [WEIGHT_SIZE-1:0] Wgt_7_447;input [WEIGHT_SIZE-1:0] Wgt_7_448;input [WEIGHT_SIZE-1:0] Wgt_7_449;input [WEIGHT_SIZE-1:0] Wgt_7_450;input [WEIGHT_SIZE-1:0] Wgt_7_451;input [WEIGHT_SIZE-1:0] Wgt_7_452;input [WEIGHT_SIZE-1:0] Wgt_7_453;input [WEIGHT_SIZE-1:0] Wgt_7_454;input [WEIGHT_SIZE-1:0] Wgt_7_455;input [WEIGHT_SIZE-1:0] Wgt_7_456;input [WEIGHT_SIZE-1:0] Wgt_7_457;input [WEIGHT_SIZE-1:0] Wgt_7_458;input [WEIGHT_SIZE-1:0] Wgt_7_459;input [WEIGHT_SIZE-1:0] Wgt_7_460;input [WEIGHT_SIZE-1:0] Wgt_7_461;input [WEIGHT_SIZE-1:0] Wgt_7_462;input [WEIGHT_SIZE-1:0] Wgt_7_463;input [WEIGHT_SIZE-1:0] Wgt_7_464;input [WEIGHT_SIZE-1:0] Wgt_7_465;input [WEIGHT_SIZE-1:0] Wgt_7_466;input [WEIGHT_SIZE-1:0] Wgt_7_467;input [WEIGHT_SIZE-1:0] Wgt_7_468;input [WEIGHT_SIZE-1:0] Wgt_7_469;input [WEIGHT_SIZE-1:0] Wgt_7_470;input [WEIGHT_SIZE-1:0] Wgt_7_471;input [WEIGHT_SIZE-1:0] Wgt_7_472;input [WEIGHT_SIZE-1:0] Wgt_7_473;input [WEIGHT_SIZE-1:0] Wgt_7_474;input [WEIGHT_SIZE-1:0] Wgt_7_475;input [WEIGHT_SIZE-1:0] Wgt_7_476;input [WEIGHT_SIZE-1:0] Wgt_7_477;input [WEIGHT_SIZE-1:0] Wgt_7_478;input [WEIGHT_SIZE-1:0] Wgt_7_479;input [WEIGHT_SIZE-1:0] Wgt_7_480;input [WEIGHT_SIZE-1:0] Wgt_7_481;input [WEIGHT_SIZE-1:0] Wgt_7_482;input [WEIGHT_SIZE-1:0] Wgt_7_483;input [WEIGHT_SIZE-1:0] Wgt_7_484;input [WEIGHT_SIZE-1:0] Wgt_7_485;input [WEIGHT_SIZE-1:0] Wgt_7_486;input [WEIGHT_SIZE-1:0] Wgt_7_487;input [WEIGHT_SIZE-1:0] Wgt_7_488;input [WEIGHT_SIZE-1:0] Wgt_7_489;input [WEIGHT_SIZE-1:0] Wgt_7_490;input [WEIGHT_SIZE-1:0] Wgt_7_491;input [WEIGHT_SIZE-1:0] Wgt_7_492;input [WEIGHT_SIZE-1:0] Wgt_7_493;input [WEIGHT_SIZE-1:0] Wgt_7_494;input [WEIGHT_SIZE-1:0] Wgt_7_495;input [WEIGHT_SIZE-1:0] Wgt_7_496;input [WEIGHT_SIZE-1:0] Wgt_7_497;input [WEIGHT_SIZE-1:0] Wgt_7_498;input [WEIGHT_SIZE-1:0] Wgt_7_499;input [WEIGHT_SIZE-1:0] Wgt_7_500;input [WEIGHT_SIZE-1:0] Wgt_7_501;input [WEIGHT_SIZE-1:0] Wgt_7_502;input [WEIGHT_SIZE-1:0] Wgt_7_503;input [WEIGHT_SIZE-1:0] Wgt_7_504;input [WEIGHT_SIZE-1:0] Wgt_7_505;input [WEIGHT_SIZE-1:0] Wgt_7_506;input [WEIGHT_SIZE-1:0] Wgt_7_507;input [WEIGHT_SIZE-1:0] Wgt_7_508;input [WEIGHT_SIZE-1:0] Wgt_7_509;input [WEIGHT_SIZE-1:0] Wgt_7_510;input [WEIGHT_SIZE-1:0] Wgt_7_511;input [WEIGHT_SIZE-1:0] Wgt_7_512;input [WEIGHT_SIZE-1:0] Wgt_7_513;input [WEIGHT_SIZE-1:0] Wgt_7_514;input [WEIGHT_SIZE-1:0] Wgt_7_515;input [WEIGHT_SIZE-1:0] Wgt_7_516;input [WEIGHT_SIZE-1:0] Wgt_7_517;input [WEIGHT_SIZE-1:0] Wgt_7_518;input [WEIGHT_SIZE-1:0] Wgt_7_519;input [WEIGHT_SIZE-1:0] Wgt_7_520;input [WEIGHT_SIZE-1:0] Wgt_7_521;input [WEIGHT_SIZE-1:0] Wgt_7_522;input [WEIGHT_SIZE-1:0] Wgt_7_523;input [WEIGHT_SIZE-1:0] Wgt_7_524;input [WEIGHT_SIZE-1:0] Wgt_7_525;input [WEIGHT_SIZE-1:0] Wgt_7_526;input [WEIGHT_SIZE-1:0] Wgt_7_527;input [WEIGHT_SIZE-1:0] Wgt_7_528;input [WEIGHT_SIZE-1:0] Wgt_7_529;input [WEIGHT_SIZE-1:0] Wgt_7_530;input [WEIGHT_SIZE-1:0] Wgt_7_531;input [WEIGHT_SIZE-1:0] Wgt_7_532;input [WEIGHT_SIZE-1:0] Wgt_7_533;input [WEIGHT_SIZE-1:0] Wgt_7_534;input [WEIGHT_SIZE-1:0] Wgt_7_535;input [WEIGHT_SIZE-1:0] Wgt_7_536;input [WEIGHT_SIZE-1:0] Wgt_7_537;input [WEIGHT_SIZE-1:0] Wgt_7_538;input [WEIGHT_SIZE-1:0] Wgt_7_539;input [WEIGHT_SIZE-1:0] Wgt_7_540;input [WEIGHT_SIZE-1:0] Wgt_7_541;input [WEIGHT_SIZE-1:0] Wgt_7_542;input [WEIGHT_SIZE-1:0] Wgt_7_543;input [WEIGHT_SIZE-1:0] Wgt_7_544;input [WEIGHT_SIZE-1:0] Wgt_7_545;input [WEIGHT_SIZE-1:0] Wgt_7_546;input [WEIGHT_SIZE-1:0] Wgt_7_547;input [WEIGHT_SIZE-1:0] Wgt_7_548;input [WEIGHT_SIZE-1:0] Wgt_7_549;input [WEIGHT_SIZE-1:0] Wgt_7_550;input [WEIGHT_SIZE-1:0] Wgt_7_551;input [WEIGHT_SIZE-1:0] Wgt_7_552;input [WEIGHT_SIZE-1:0] Wgt_7_553;input [WEIGHT_SIZE-1:0] Wgt_7_554;input [WEIGHT_SIZE-1:0] Wgt_7_555;input [WEIGHT_SIZE-1:0] Wgt_7_556;input [WEIGHT_SIZE-1:0] Wgt_7_557;input [WEIGHT_SIZE-1:0] Wgt_7_558;input [WEIGHT_SIZE-1:0] Wgt_7_559;input [WEIGHT_SIZE-1:0] Wgt_7_560;input [WEIGHT_SIZE-1:0] Wgt_7_561;input [WEIGHT_SIZE-1:0] Wgt_7_562;input [WEIGHT_SIZE-1:0] Wgt_7_563;input [WEIGHT_SIZE-1:0] Wgt_7_564;input [WEIGHT_SIZE-1:0] Wgt_7_565;input [WEIGHT_SIZE-1:0] Wgt_7_566;input [WEIGHT_SIZE-1:0] Wgt_7_567;input [WEIGHT_SIZE-1:0] Wgt_7_568;input [WEIGHT_SIZE-1:0] Wgt_7_569;input [WEIGHT_SIZE-1:0] Wgt_7_570;input [WEIGHT_SIZE-1:0] Wgt_7_571;input [WEIGHT_SIZE-1:0] Wgt_7_572;input [WEIGHT_SIZE-1:0] Wgt_7_573;input [WEIGHT_SIZE-1:0] Wgt_7_574;input [WEIGHT_SIZE-1:0] Wgt_7_575;input [WEIGHT_SIZE-1:0] Wgt_7_576;input [WEIGHT_SIZE-1:0] Wgt_7_577;input [WEIGHT_SIZE-1:0] Wgt_7_578;input [WEIGHT_SIZE-1:0] Wgt_7_579;input [WEIGHT_SIZE-1:0] Wgt_7_580;input [WEIGHT_SIZE-1:0] Wgt_7_581;input [WEIGHT_SIZE-1:0] Wgt_7_582;input [WEIGHT_SIZE-1:0] Wgt_7_583;input [WEIGHT_SIZE-1:0] Wgt_7_584;input [WEIGHT_SIZE-1:0] Wgt_7_585;input [WEIGHT_SIZE-1:0] Wgt_7_586;input [WEIGHT_SIZE-1:0] Wgt_7_587;input [WEIGHT_SIZE-1:0] Wgt_7_588;input [WEIGHT_SIZE-1:0] Wgt_7_589;input [WEIGHT_SIZE-1:0] Wgt_7_590;input [WEIGHT_SIZE-1:0] Wgt_7_591;input [WEIGHT_SIZE-1:0] Wgt_7_592;input [WEIGHT_SIZE-1:0] Wgt_7_593;input [WEIGHT_SIZE-1:0] Wgt_7_594;input [WEIGHT_SIZE-1:0] Wgt_7_595;input [WEIGHT_SIZE-1:0] Wgt_7_596;input [WEIGHT_SIZE-1:0] Wgt_7_597;input [WEIGHT_SIZE-1:0] Wgt_7_598;input [WEIGHT_SIZE-1:0] Wgt_7_599;input [WEIGHT_SIZE-1:0] Wgt_7_600;input [WEIGHT_SIZE-1:0] Wgt_7_601;input [WEIGHT_SIZE-1:0] Wgt_7_602;input [WEIGHT_SIZE-1:0] Wgt_7_603;input [WEIGHT_SIZE-1:0] Wgt_7_604;input [WEIGHT_SIZE-1:0] Wgt_7_605;input [WEIGHT_SIZE-1:0] Wgt_7_606;input [WEIGHT_SIZE-1:0] Wgt_7_607;input [WEIGHT_SIZE-1:0] Wgt_7_608;input [WEIGHT_SIZE-1:0] Wgt_7_609;input [WEIGHT_SIZE-1:0] Wgt_7_610;input [WEIGHT_SIZE-1:0] Wgt_7_611;input [WEIGHT_SIZE-1:0] Wgt_7_612;input [WEIGHT_SIZE-1:0] Wgt_7_613;input [WEIGHT_SIZE-1:0] Wgt_7_614;input [WEIGHT_SIZE-1:0] Wgt_7_615;input [WEIGHT_SIZE-1:0] Wgt_7_616;input [WEIGHT_SIZE-1:0] Wgt_7_617;input [WEIGHT_SIZE-1:0] Wgt_7_618;input [WEIGHT_SIZE-1:0] Wgt_7_619;input [WEIGHT_SIZE-1:0] Wgt_7_620;input [WEIGHT_SIZE-1:0] Wgt_7_621;input [WEIGHT_SIZE-1:0] Wgt_7_622;input [WEIGHT_SIZE-1:0] Wgt_7_623;input [WEIGHT_SIZE-1:0] Wgt_7_624;input [WEIGHT_SIZE-1:0] Wgt_7_625;input [WEIGHT_SIZE-1:0] Wgt_7_626;input [WEIGHT_SIZE-1:0] Wgt_7_627;input [WEIGHT_SIZE-1:0] Wgt_7_628;input [WEIGHT_SIZE-1:0] Wgt_7_629;input [WEIGHT_SIZE-1:0] Wgt_7_630;input [WEIGHT_SIZE-1:0] Wgt_7_631;input [WEIGHT_SIZE-1:0] Wgt_7_632;input [WEIGHT_SIZE-1:0] Wgt_7_633;input [WEIGHT_SIZE-1:0] Wgt_7_634;input [WEIGHT_SIZE-1:0] Wgt_7_635;input [WEIGHT_SIZE-1:0] Wgt_7_636;input [WEIGHT_SIZE-1:0] Wgt_7_637;input [WEIGHT_SIZE-1:0] Wgt_7_638;input [WEIGHT_SIZE-1:0] Wgt_7_639;input [WEIGHT_SIZE-1:0] Wgt_7_640;input [WEIGHT_SIZE-1:0] Wgt_7_641;input [WEIGHT_SIZE-1:0] Wgt_7_642;input [WEIGHT_SIZE-1:0] Wgt_7_643;input [WEIGHT_SIZE-1:0] Wgt_7_644;input [WEIGHT_SIZE-1:0] Wgt_7_645;input [WEIGHT_SIZE-1:0] Wgt_7_646;input [WEIGHT_SIZE-1:0] Wgt_7_647;input [WEIGHT_SIZE-1:0] Wgt_7_648;input [WEIGHT_SIZE-1:0] Wgt_7_649;input [WEIGHT_SIZE-1:0] Wgt_7_650;input [WEIGHT_SIZE-1:0] Wgt_7_651;input [WEIGHT_SIZE-1:0] Wgt_7_652;input [WEIGHT_SIZE-1:0] Wgt_7_653;input [WEIGHT_SIZE-1:0] Wgt_7_654;input [WEIGHT_SIZE-1:0] Wgt_7_655;input [WEIGHT_SIZE-1:0] Wgt_7_656;input [WEIGHT_SIZE-1:0] Wgt_7_657;input [WEIGHT_SIZE-1:0] Wgt_7_658;input [WEIGHT_SIZE-1:0] Wgt_7_659;input [WEIGHT_SIZE-1:0] Wgt_7_660;input [WEIGHT_SIZE-1:0] Wgt_7_661;input [WEIGHT_SIZE-1:0] Wgt_7_662;input [WEIGHT_SIZE-1:0] Wgt_7_663;input [WEIGHT_SIZE-1:0] Wgt_7_664;input [WEIGHT_SIZE-1:0] Wgt_7_665;input [WEIGHT_SIZE-1:0] Wgt_7_666;input [WEIGHT_SIZE-1:0] Wgt_7_667;input [WEIGHT_SIZE-1:0] Wgt_7_668;input [WEIGHT_SIZE-1:0] Wgt_7_669;input [WEIGHT_SIZE-1:0] Wgt_7_670;input [WEIGHT_SIZE-1:0] Wgt_7_671;input [WEIGHT_SIZE-1:0] Wgt_7_672;input [WEIGHT_SIZE-1:0] Wgt_7_673;input [WEIGHT_SIZE-1:0] Wgt_7_674;input [WEIGHT_SIZE-1:0] Wgt_7_675;input [WEIGHT_SIZE-1:0] Wgt_7_676;input [WEIGHT_SIZE-1:0] Wgt_7_677;input [WEIGHT_SIZE-1:0] Wgt_7_678;input [WEIGHT_SIZE-1:0] Wgt_7_679;input [WEIGHT_SIZE-1:0] Wgt_7_680;input [WEIGHT_SIZE-1:0] Wgt_7_681;input [WEIGHT_SIZE-1:0] Wgt_7_682;input [WEIGHT_SIZE-1:0] Wgt_7_683;input [WEIGHT_SIZE-1:0] Wgt_7_684;input [WEIGHT_SIZE-1:0] Wgt_7_685;input [WEIGHT_SIZE-1:0] Wgt_7_686;input [WEIGHT_SIZE-1:0] Wgt_7_687;input [WEIGHT_SIZE-1:0] Wgt_7_688;input [WEIGHT_SIZE-1:0] Wgt_7_689;input [WEIGHT_SIZE-1:0] Wgt_7_690;input [WEIGHT_SIZE-1:0] Wgt_7_691;input [WEIGHT_SIZE-1:0] Wgt_7_692;input [WEIGHT_SIZE-1:0] Wgt_7_693;input [WEIGHT_SIZE-1:0] Wgt_7_694;input [WEIGHT_SIZE-1:0] Wgt_7_695;input [WEIGHT_SIZE-1:0] Wgt_7_696;input [WEIGHT_SIZE-1:0] Wgt_7_697;input [WEIGHT_SIZE-1:0] Wgt_7_698;input [WEIGHT_SIZE-1:0] Wgt_7_699;input [WEIGHT_SIZE-1:0] Wgt_7_700;input [WEIGHT_SIZE-1:0] Wgt_7_701;input [WEIGHT_SIZE-1:0] Wgt_7_702;input [WEIGHT_SIZE-1:0] Wgt_7_703;input [WEIGHT_SIZE-1:0] Wgt_7_704;input [WEIGHT_SIZE-1:0] Wgt_7_705;input [WEIGHT_SIZE-1:0] Wgt_7_706;input [WEIGHT_SIZE-1:0] Wgt_7_707;input [WEIGHT_SIZE-1:0] Wgt_7_708;input [WEIGHT_SIZE-1:0] Wgt_7_709;input [WEIGHT_SIZE-1:0] Wgt_7_710;input [WEIGHT_SIZE-1:0] Wgt_7_711;input [WEIGHT_SIZE-1:0] Wgt_7_712;input [WEIGHT_SIZE-1:0] Wgt_7_713;input [WEIGHT_SIZE-1:0] Wgt_7_714;input [WEIGHT_SIZE-1:0] Wgt_7_715;input [WEIGHT_SIZE-1:0] Wgt_7_716;input [WEIGHT_SIZE-1:0] Wgt_7_717;input [WEIGHT_SIZE-1:0] Wgt_7_718;input [WEIGHT_SIZE-1:0] Wgt_7_719;input [WEIGHT_SIZE-1:0] Wgt_7_720;input [WEIGHT_SIZE-1:0] Wgt_7_721;input [WEIGHT_SIZE-1:0] Wgt_7_722;input [WEIGHT_SIZE-1:0] Wgt_7_723;input [WEIGHT_SIZE-1:0] Wgt_7_724;input [WEIGHT_SIZE-1:0] Wgt_7_725;input [WEIGHT_SIZE-1:0] Wgt_7_726;input [WEIGHT_SIZE-1:0] Wgt_7_727;input [WEIGHT_SIZE-1:0] Wgt_7_728;input [WEIGHT_SIZE-1:0] Wgt_7_729;input [WEIGHT_SIZE-1:0] Wgt_7_730;input [WEIGHT_SIZE-1:0] Wgt_7_731;input [WEIGHT_SIZE-1:0] Wgt_7_732;input [WEIGHT_SIZE-1:0] Wgt_7_733;input [WEIGHT_SIZE-1:0] Wgt_7_734;input [WEIGHT_SIZE-1:0] Wgt_7_735;input [WEIGHT_SIZE-1:0] Wgt_7_736;input [WEIGHT_SIZE-1:0] Wgt_7_737;input [WEIGHT_SIZE-1:0] Wgt_7_738;input [WEIGHT_SIZE-1:0] Wgt_7_739;input [WEIGHT_SIZE-1:0] Wgt_7_740;input [WEIGHT_SIZE-1:0] Wgt_7_741;input [WEIGHT_SIZE-1:0] Wgt_7_742;input [WEIGHT_SIZE-1:0] Wgt_7_743;input [WEIGHT_SIZE-1:0] Wgt_7_744;input [WEIGHT_SIZE-1:0] Wgt_7_745;input [WEIGHT_SIZE-1:0] Wgt_7_746;input [WEIGHT_SIZE-1:0] Wgt_7_747;input [WEIGHT_SIZE-1:0] Wgt_7_748;input [WEIGHT_SIZE-1:0] Wgt_7_749;input [WEIGHT_SIZE-1:0] Wgt_7_750;input [WEIGHT_SIZE-1:0] Wgt_7_751;input [WEIGHT_SIZE-1:0] Wgt_7_752;input [WEIGHT_SIZE-1:0] Wgt_7_753;input [WEIGHT_SIZE-1:0] Wgt_7_754;input [WEIGHT_SIZE-1:0] Wgt_7_755;input [WEIGHT_SIZE-1:0] Wgt_7_756;input [WEIGHT_SIZE-1:0] Wgt_7_757;input [WEIGHT_SIZE-1:0] Wgt_7_758;input [WEIGHT_SIZE-1:0] Wgt_7_759;input [WEIGHT_SIZE-1:0] Wgt_7_760;input [WEIGHT_SIZE-1:0] Wgt_7_761;input [WEIGHT_SIZE-1:0] Wgt_7_762;input [WEIGHT_SIZE-1:0] Wgt_7_763;input [WEIGHT_SIZE-1:0] Wgt_7_764;input [WEIGHT_SIZE-1:0] Wgt_7_765;input [WEIGHT_SIZE-1:0] Wgt_7_766;input [WEIGHT_SIZE-1:0] Wgt_7_767;input [WEIGHT_SIZE-1:0] Wgt_7_768;input [WEIGHT_SIZE-1:0] Wgt_7_769;input [WEIGHT_SIZE-1:0] Wgt_7_770;input [WEIGHT_SIZE-1:0] Wgt_7_771;input [WEIGHT_SIZE-1:0] Wgt_7_772;input [WEIGHT_SIZE-1:0] Wgt_7_773;input [WEIGHT_SIZE-1:0] Wgt_7_774;input [WEIGHT_SIZE-1:0] Wgt_7_775;input [WEIGHT_SIZE-1:0] Wgt_7_776;input [WEIGHT_SIZE-1:0] Wgt_7_777;input [WEIGHT_SIZE-1:0] Wgt_7_778;input [WEIGHT_SIZE-1:0] Wgt_7_779;input [WEIGHT_SIZE-1:0] Wgt_7_780;input [WEIGHT_SIZE-1:0] Wgt_7_781;input [WEIGHT_SIZE-1:0] Wgt_7_782;input [WEIGHT_SIZE-1:0] Wgt_7_783;input [WEIGHT_SIZE-1:0] Wgt_7_784;input [WEIGHT_SIZE-1:0] Wgt_8_0;input [WEIGHT_SIZE-1:0] Wgt_8_1;input [WEIGHT_SIZE-1:0] Wgt_8_2;input [WEIGHT_SIZE-1:0] Wgt_8_3;input [WEIGHT_SIZE-1:0] Wgt_8_4;input [WEIGHT_SIZE-1:0] Wgt_8_5;input [WEIGHT_SIZE-1:0] Wgt_8_6;input [WEIGHT_SIZE-1:0] Wgt_8_7;input [WEIGHT_SIZE-1:0] Wgt_8_8;input [WEIGHT_SIZE-1:0] Wgt_8_9;input [WEIGHT_SIZE-1:0] Wgt_8_10;input [WEIGHT_SIZE-1:0] Wgt_8_11;input [WEIGHT_SIZE-1:0] Wgt_8_12;input [WEIGHT_SIZE-1:0] Wgt_8_13;input [WEIGHT_SIZE-1:0] Wgt_8_14;input [WEIGHT_SIZE-1:0] Wgt_8_15;input [WEIGHT_SIZE-1:0] Wgt_8_16;input [WEIGHT_SIZE-1:0] Wgt_8_17;input [WEIGHT_SIZE-1:0] Wgt_8_18;input [WEIGHT_SIZE-1:0] Wgt_8_19;input [WEIGHT_SIZE-1:0] Wgt_8_20;input [WEIGHT_SIZE-1:0] Wgt_8_21;input [WEIGHT_SIZE-1:0] Wgt_8_22;input [WEIGHT_SIZE-1:0] Wgt_8_23;input [WEIGHT_SIZE-1:0] Wgt_8_24;input [WEIGHT_SIZE-1:0] Wgt_8_25;input [WEIGHT_SIZE-1:0] Wgt_8_26;input [WEIGHT_SIZE-1:0] Wgt_8_27;input [WEIGHT_SIZE-1:0] Wgt_8_28;input [WEIGHT_SIZE-1:0] Wgt_8_29;input [WEIGHT_SIZE-1:0] Wgt_8_30;input [WEIGHT_SIZE-1:0] Wgt_8_31;input [WEIGHT_SIZE-1:0] Wgt_8_32;input [WEIGHT_SIZE-1:0] Wgt_8_33;input [WEIGHT_SIZE-1:0] Wgt_8_34;input [WEIGHT_SIZE-1:0] Wgt_8_35;input [WEIGHT_SIZE-1:0] Wgt_8_36;input [WEIGHT_SIZE-1:0] Wgt_8_37;input [WEIGHT_SIZE-1:0] Wgt_8_38;input [WEIGHT_SIZE-1:0] Wgt_8_39;input [WEIGHT_SIZE-1:0] Wgt_8_40;input [WEIGHT_SIZE-1:0] Wgt_8_41;input [WEIGHT_SIZE-1:0] Wgt_8_42;input [WEIGHT_SIZE-1:0] Wgt_8_43;input [WEIGHT_SIZE-1:0] Wgt_8_44;input [WEIGHT_SIZE-1:0] Wgt_8_45;input [WEIGHT_SIZE-1:0] Wgt_8_46;input [WEIGHT_SIZE-1:0] Wgt_8_47;input [WEIGHT_SIZE-1:0] Wgt_8_48;input [WEIGHT_SIZE-1:0] Wgt_8_49;input [WEIGHT_SIZE-1:0] Wgt_8_50;input [WEIGHT_SIZE-1:0] Wgt_8_51;input [WEIGHT_SIZE-1:0] Wgt_8_52;input [WEIGHT_SIZE-1:0] Wgt_8_53;input [WEIGHT_SIZE-1:0] Wgt_8_54;input [WEIGHT_SIZE-1:0] Wgt_8_55;input [WEIGHT_SIZE-1:0] Wgt_8_56;input [WEIGHT_SIZE-1:0] Wgt_8_57;input [WEIGHT_SIZE-1:0] Wgt_8_58;input [WEIGHT_SIZE-1:0] Wgt_8_59;input [WEIGHT_SIZE-1:0] Wgt_8_60;input [WEIGHT_SIZE-1:0] Wgt_8_61;input [WEIGHT_SIZE-1:0] Wgt_8_62;input [WEIGHT_SIZE-1:0] Wgt_8_63;input [WEIGHT_SIZE-1:0] Wgt_8_64;input [WEIGHT_SIZE-1:0] Wgt_8_65;input [WEIGHT_SIZE-1:0] Wgt_8_66;input [WEIGHT_SIZE-1:0] Wgt_8_67;input [WEIGHT_SIZE-1:0] Wgt_8_68;input [WEIGHT_SIZE-1:0] Wgt_8_69;input [WEIGHT_SIZE-1:0] Wgt_8_70;input [WEIGHT_SIZE-1:0] Wgt_8_71;input [WEIGHT_SIZE-1:0] Wgt_8_72;input [WEIGHT_SIZE-1:0] Wgt_8_73;input [WEIGHT_SIZE-1:0] Wgt_8_74;input [WEIGHT_SIZE-1:0] Wgt_8_75;input [WEIGHT_SIZE-1:0] Wgt_8_76;input [WEIGHT_SIZE-1:0] Wgt_8_77;input [WEIGHT_SIZE-1:0] Wgt_8_78;input [WEIGHT_SIZE-1:0] Wgt_8_79;input [WEIGHT_SIZE-1:0] Wgt_8_80;input [WEIGHT_SIZE-1:0] Wgt_8_81;input [WEIGHT_SIZE-1:0] Wgt_8_82;input [WEIGHT_SIZE-1:0] Wgt_8_83;input [WEIGHT_SIZE-1:0] Wgt_8_84;input [WEIGHT_SIZE-1:0] Wgt_8_85;input [WEIGHT_SIZE-1:0] Wgt_8_86;input [WEIGHT_SIZE-1:0] Wgt_8_87;input [WEIGHT_SIZE-1:0] Wgt_8_88;input [WEIGHT_SIZE-1:0] Wgt_8_89;input [WEIGHT_SIZE-1:0] Wgt_8_90;input [WEIGHT_SIZE-1:0] Wgt_8_91;input [WEIGHT_SIZE-1:0] Wgt_8_92;input [WEIGHT_SIZE-1:0] Wgt_8_93;input [WEIGHT_SIZE-1:0] Wgt_8_94;input [WEIGHT_SIZE-1:0] Wgt_8_95;input [WEIGHT_SIZE-1:0] Wgt_8_96;input [WEIGHT_SIZE-1:0] Wgt_8_97;input [WEIGHT_SIZE-1:0] Wgt_8_98;input [WEIGHT_SIZE-1:0] Wgt_8_99;input [WEIGHT_SIZE-1:0] Wgt_8_100;input [WEIGHT_SIZE-1:0] Wgt_8_101;input [WEIGHT_SIZE-1:0] Wgt_8_102;input [WEIGHT_SIZE-1:0] Wgt_8_103;input [WEIGHT_SIZE-1:0] Wgt_8_104;input [WEIGHT_SIZE-1:0] Wgt_8_105;input [WEIGHT_SIZE-1:0] Wgt_8_106;input [WEIGHT_SIZE-1:0] Wgt_8_107;input [WEIGHT_SIZE-1:0] Wgt_8_108;input [WEIGHT_SIZE-1:0] Wgt_8_109;input [WEIGHT_SIZE-1:0] Wgt_8_110;input [WEIGHT_SIZE-1:0] Wgt_8_111;input [WEIGHT_SIZE-1:0] Wgt_8_112;input [WEIGHT_SIZE-1:0] Wgt_8_113;input [WEIGHT_SIZE-1:0] Wgt_8_114;input [WEIGHT_SIZE-1:0] Wgt_8_115;input [WEIGHT_SIZE-1:0] Wgt_8_116;input [WEIGHT_SIZE-1:0] Wgt_8_117;input [WEIGHT_SIZE-1:0] Wgt_8_118;input [WEIGHT_SIZE-1:0] Wgt_8_119;input [WEIGHT_SIZE-1:0] Wgt_8_120;input [WEIGHT_SIZE-1:0] Wgt_8_121;input [WEIGHT_SIZE-1:0] Wgt_8_122;input [WEIGHT_SIZE-1:0] Wgt_8_123;input [WEIGHT_SIZE-1:0] Wgt_8_124;input [WEIGHT_SIZE-1:0] Wgt_8_125;input [WEIGHT_SIZE-1:0] Wgt_8_126;input [WEIGHT_SIZE-1:0] Wgt_8_127;input [WEIGHT_SIZE-1:0] Wgt_8_128;input [WEIGHT_SIZE-1:0] Wgt_8_129;input [WEIGHT_SIZE-1:0] Wgt_8_130;input [WEIGHT_SIZE-1:0] Wgt_8_131;input [WEIGHT_SIZE-1:0] Wgt_8_132;input [WEIGHT_SIZE-1:0] Wgt_8_133;input [WEIGHT_SIZE-1:0] Wgt_8_134;input [WEIGHT_SIZE-1:0] Wgt_8_135;input [WEIGHT_SIZE-1:0] Wgt_8_136;input [WEIGHT_SIZE-1:0] Wgt_8_137;input [WEIGHT_SIZE-1:0] Wgt_8_138;input [WEIGHT_SIZE-1:0] Wgt_8_139;input [WEIGHT_SIZE-1:0] Wgt_8_140;input [WEIGHT_SIZE-1:0] Wgt_8_141;input [WEIGHT_SIZE-1:0] Wgt_8_142;input [WEIGHT_SIZE-1:0] Wgt_8_143;input [WEIGHT_SIZE-1:0] Wgt_8_144;input [WEIGHT_SIZE-1:0] Wgt_8_145;input [WEIGHT_SIZE-1:0] Wgt_8_146;input [WEIGHT_SIZE-1:0] Wgt_8_147;input [WEIGHT_SIZE-1:0] Wgt_8_148;input [WEIGHT_SIZE-1:0] Wgt_8_149;input [WEIGHT_SIZE-1:0] Wgt_8_150;input [WEIGHT_SIZE-1:0] Wgt_8_151;input [WEIGHT_SIZE-1:0] Wgt_8_152;input [WEIGHT_SIZE-1:0] Wgt_8_153;input [WEIGHT_SIZE-1:0] Wgt_8_154;input [WEIGHT_SIZE-1:0] Wgt_8_155;input [WEIGHT_SIZE-1:0] Wgt_8_156;input [WEIGHT_SIZE-1:0] Wgt_8_157;input [WEIGHT_SIZE-1:0] Wgt_8_158;input [WEIGHT_SIZE-1:0] Wgt_8_159;input [WEIGHT_SIZE-1:0] Wgt_8_160;input [WEIGHT_SIZE-1:0] Wgt_8_161;input [WEIGHT_SIZE-1:0] Wgt_8_162;input [WEIGHT_SIZE-1:0] Wgt_8_163;input [WEIGHT_SIZE-1:0] Wgt_8_164;input [WEIGHT_SIZE-1:0] Wgt_8_165;input [WEIGHT_SIZE-1:0] Wgt_8_166;input [WEIGHT_SIZE-1:0] Wgt_8_167;input [WEIGHT_SIZE-1:0] Wgt_8_168;input [WEIGHT_SIZE-1:0] Wgt_8_169;input [WEIGHT_SIZE-1:0] Wgt_8_170;input [WEIGHT_SIZE-1:0] Wgt_8_171;input [WEIGHT_SIZE-1:0] Wgt_8_172;input [WEIGHT_SIZE-1:0] Wgt_8_173;input [WEIGHT_SIZE-1:0] Wgt_8_174;input [WEIGHT_SIZE-1:0] Wgt_8_175;input [WEIGHT_SIZE-1:0] Wgt_8_176;input [WEIGHT_SIZE-1:0] Wgt_8_177;input [WEIGHT_SIZE-1:0] Wgt_8_178;input [WEIGHT_SIZE-1:0] Wgt_8_179;input [WEIGHT_SIZE-1:0] Wgt_8_180;input [WEIGHT_SIZE-1:0] Wgt_8_181;input [WEIGHT_SIZE-1:0] Wgt_8_182;input [WEIGHT_SIZE-1:0] Wgt_8_183;input [WEIGHT_SIZE-1:0] Wgt_8_184;input [WEIGHT_SIZE-1:0] Wgt_8_185;input [WEIGHT_SIZE-1:0] Wgt_8_186;input [WEIGHT_SIZE-1:0] Wgt_8_187;input [WEIGHT_SIZE-1:0] Wgt_8_188;input [WEIGHT_SIZE-1:0] Wgt_8_189;input [WEIGHT_SIZE-1:0] Wgt_8_190;input [WEIGHT_SIZE-1:0] Wgt_8_191;input [WEIGHT_SIZE-1:0] Wgt_8_192;input [WEIGHT_SIZE-1:0] Wgt_8_193;input [WEIGHT_SIZE-1:0] Wgt_8_194;input [WEIGHT_SIZE-1:0] Wgt_8_195;input [WEIGHT_SIZE-1:0] Wgt_8_196;input [WEIGHT_SIZE-1:0] Wgt_8_197;input [WEIGHT_SIZE-1:0] Wgt_8_198;input [WEIGHT_SIZE-1:0] Wgt_8_199;input [WEIGHT_SIZE-1:0] Wgt_8_200;input [WEIGHT_SIZE-1:0] Wgt_8_201;input [WEIGHT_SIZE-1:0] Wgt_8_202;input [WEIGHT_SIZE-1:0] Wgt_8_203;input [WEIGHT_SIZE-1:0] Wgt_8_204;input [WEIGHT_SIZE-1:0] Wgt_8_205;input [WEIGHT_SIZE-1:0] Wgt_8_206;input [WEIGHT_SIZE-1:0] Wgt_8_207;input [WEIGHT_SIZE-1:0] Wgt_8_208;input [WEIGHT_SIZE-1:0] Wgt_8_209;input [WEIGHT_SIZE-1:0] Wgt_8_210;input [WEIGHT_SIZE-1:0] Wgt_8_211;input [WEIGHT_SIZE-1:0] Wgt_8_212;input [WEIGHT_SIZE-1:0] Wgt_8_213;input [WEIGHT_SIZE-1:0] Wgt_8_214;input [WEIGHT_SIZE-1:0] Wgt_8_215;input [WEIGHT_SIZE-1:0] Wgt_8_216;input [WEIGHT_SIZE-1:0] Wgt_8_217;input [WEIGHT_SIZE-1:0] Wgt_8_218;input [WEIGHT_SIZE-1:0] Wgt_8_219;input [WEIGHT_SIZE-1:0] Wgt_8_220;input [WEIGHT_SIZE-1:0] Wgt_8_221;input [WEIGHT_SIZE-1:0] Wgt_8_222;input [WEIGHT_SIZE-1:0] Wgt_8_223;input [WEIGHT_SIZE-1:0] Wgt_8_224;input [WEIGHT_SIZE-1:0] Wgt_8_225;input [WEIGHT_SIZE-1:0] Wgt_8_226;input [WEIGHT_SIZE-1:0] Wgt_8_227;input [WEIGHT_SIZE-1:0] Wgt_8_228;input [WEIGHT_SIZE-1:0] Wgt_8_229;input [WEIGHT_SIZE-1:0] Wgt_8_230;input [WEIGHT_SIZE-1:0] Wgt_8_231;input [WEIGHT_SIZE-1:0] Wgt_8_232;input [WEIGHT_SIZE-1:0] Wgt_8_233;input [WEIGHT_SIZE-1:0] Wgt_8_234;input [WEIGHT_SIZE-1:0] Wgt_8_235;input [WEIGHT_SIZE-1:0] Wgt_8_236;input [WEIGHT_SIZE-1:0] Wgt_8_237;input [WEIGHT_SIZE-1:0] Wgt_8_238;input [WEIGHT_SIZE-1:0] Wgt_8_239;input [WEIGHT_SIZE-1:0] Wgt_8_240;input [WEIGHT_SIZE-1:0] Wgt_8_241;input [WEIGHT_SIZE-1:0] Wgt_8_242;input [WEIGHT_SIZE-1:0] Wgt_8_243;input [WEIGHT_SIZE-1:0] Wgt_8_244;input [WEIGHT_SIZE-1:0] Wgt_8_245;input [WEIGHT_SIZE-1:0] Wgt_8_246;input [WEIGHT_SIZE-1:0] Wgt_8_247;input [WEIGHT_SIZE-1:0] Wgt_8_248;input [WEIGHT_SIZE-1:0] Wgt_8_249;input [WEIGHT_SIZE-1:0] Wgt_8_250;input [WEIGHT_SIZE-1:0] Wgt_8_251;input [WEIGHT_SIZE-1:0] Wgt_8_252;input [WEIGHT_SIZE-1:0] Wgt_8_253;input [WEIGHT_SIZE-1:0] Wgt_8_254;input [WEIGHT_SIZE-1:0] Wgt_8_255;input [WEIGHT_SIZE-1:0] Wgt_8_256;input [WEIGHT_SIZE-1:0] Wgt_8_257;input [WEIGHT_SIZE-1:0] Wgt_8_258;input [WEIGHT_SIZE-1:0] Wgt_8_259;input [WEIGHT_SIZE-1:0] Wgt_8_260;input [WEIGHT_SIZE-1:0] Wgt_8_261;input [WEIGHT_SIZE-1:0] Wgt_8_262;input [WEIGHT_SIZE-1:0] Wgt_8_263;input [WEIGHT_SIZE-1:0] Wgt_8_264;input [WEIGHT_SIZE-1:0] Wgt_8_265;input [WEIGHT_SIZE-1:0] Wgt_8_266;input [WEIGHT_SIZE-1:0] Wgt_8_267;input [WEIGHT_SIZE-1:0] Wgt_8_268;input [WEIGHT_SIZE-1:0] Wgt_8_269;input [WEIGHT_SIZE-1:0] Wgt_8_270;input [WEIGHT_SIZE-1:0] Wgt_8_271;input [WEIGHT_SIZE-1:0] Wgt_8_272;input [WEIGHT_SIZE-1:0] Wgt_8_273;input [WEIGHT_SIZE-1:0] Wgt_8_274;input [WEIGHT_SIZE-1:0] Wgt_8_275;input [WEIGHT_SIZE-1:0] Wgt_8_276;input [WEIGHT_SIZE-1:0] Wgt_8_277;input [WEIGHT_SIZE-1:0] Wgt_8_278;input [WEIGHT_SIZE-1:0] Wgt_8_279;input [WEIGHT_SIZE-1:0] Wgt_8_280;input [WEIGHT_SIZE-1:0] Wgt_8_281;input [WEIGHT_SIZE-1:0] Wgt_8_282;input [WEIGHT_SIZE-1:0] Wgt_8_283;input [WEIGHT_SIZE-1:0] Wgt_8_284;input [WEIGHT_SIZE-1:0] Wgt_8_285;input [WEIGHT_SIZE-1:0] Wgt_8_286;input [WEIGHT_SIZE-1:0] Wgt_8_287;input [WEIGHT_SIZE-1:0] Wgt_8_288;input [WEIGHT_SIZE-1:0] Wgt_8_289;input [WEIGHT_SIZE-1:0] Wgt_8_290;input [WEIGHT_SIZE-1:0] Wgt_8_291;input [WEIGHT_SIZE-1:0] Wgt_8_292;input [WEIGHT_SIZE-1:0] Wgt_8_293;input [WEIGHT_SIZE-1:0] Wgt_8_294;input [WEIGHT_SIZE-1:0] Wgt_8_295;input [WEIGHT_SIZE-1:0] Wgt_8_296;input [WEIGHT_SIZE-1:0] Wgt_8_297;input [WEIGHT_SIZE-1:0] Wgt_8_298;input [WEIGHT_SIZE-1:0] Wgt_8_299;input [WEIGHT_SIZE-1:0] Wgt_8_300;input [WEIGHT_SIZE-1:0] Wgt_8_301;input [WEIGHT_SIZE-1:0] Wgt_8_302;input [WEIGHT_SIZE-1:0] Wgt_8_303;input [WEIGHT_SIZE-1:0] Wgt_8_304;input [WEIGHT_SIZE-1:0] Wgt_8_305;input [WEIGHT_SIZE-1:0] Wgt_8_306;input [WEIGHT_SIZE-1:0] Wgt_8_307;input [WEIGHT_SIZE-1:0] Wgt_8_308;input [WEIGHT_SIZE-1:0] Wgt_8_309;input [WEIGHT_SIZE-1:0] Wgt_8_310;input [WEIGHT_SIZE-1:0] Wgt_8_311;input [WEIGHT_SIZE-1:0] Wgt_8_312;input [WEIGHT_SIZE-1:0] Wgt_8_313;input [WEIGHT_SIZE-1:0] Wgt_8_314;input [WEIGHT_SIZE-1:0] Wgt_8_315;input [WEIGHT_SIZE-1:0] Wgt_8_316;input [WEIGHT_SIZE-1:0] Wgt_8_317;input [WEIGHT_SIZE-1:0] Wgt_8_318;input [WEIGHT_SIZE-1:0] Wgt_8_319;input [WEIGHT_SIZE-1:0] Wgt_8_320;input [WEIGHT_SIZE-1:0] Wgt_8_321;input [WEIGHT_SIZE-1:0] Wgt_8_322;input [WEIGHT_SIZE-1:0] Wgt_8_323;input [WEIGHT_SIZE-1:0] Wgt_8_324;input [WEIGHT_SIZE-1:0] Wgt_8_325;input [WEIGHT_SIZE-1:0] Wgt_8_326;input [WEIGHT_SIZE-1:0] Wgt_8_327;input [WEIGHT_SIZE-1:0] Wgt_8_328;input [WEIGHT_SIZE-1:0] Wgt_8_329;input [WEIGHT_SIZE-1:0] Wgt_8_330;input [WEIGHT_SIZE-1:0] Wgt_8_331;input [WEIGHT_SIZE-1:0] Wgt_8_332;input [WEIGHT_SIZE-1:0] Wgt_8_333;input [WEIGHT_SIZE-1:0] Wgt_8_334;input [WEIGHT_SIZE-1:0] Wgt_8_335;input [WEIGHT_SIZE-1:0] Wgt_8_336;input [WEIGHT_SIZE-1:0] Wgt_8_337;input [WEIGHT_SIZE-1:0] Wgt_8_338;input [WEIGHT_SIZE-1:0] Wgt_8_339;input [WEIGHT_SIZE-1:0] Wgt_8_340;input [WEIGHT_SIZE-1:0] Wgt_8_341;input [WEIGHT_SIZE-1:0] Wgt_8_342;input [WEIGHT_SIZE-1:0] Wgt_8_343;input [WEIGHT_SIZE-1:0] Wgt_8_344;input [WEIGHT_SIZE-1:0] Wgt_8_345;input [WEIGHT_SIZE-1:0] Wgt_8_346;input [WEIGHT_SIZE-1:0] Wgt_8_347;input [WEIGHT_SIZE-1:0] Wgt_8_348;input [WEIGHT_SIZE-1:0] Wgt_8_349;input [WEIGHT_SIZE-1:0] Wgt_8_350;input [WEIGHT_SIZE-1:0] Wgt_8_351;input [WEIGHT_SIZE-1:0] Wgt_8_352;input [WEIGHT_SIZE-1:0] Wgt_8_353;input [WEIGHT_SIZE-1:0] Wgt_8_354;input [WEIGHT_SIZE-1:0] Wgt_8_355;input [WEIGHT_SIZE-1:0] Wgt_8_356;input [WEIGHT_SIZE-1:0] Wgt_8_357;input [WEIGHT_SIZE-1:0] Wgt_8_358;input [WEIGHT_SIZE-1:0] Wgt_8_359;input [WEIGHT_SIZE-1:0] Wgt_8_360;input [WEIGHT_SIZE-1:0] Wgt_8_361;input [WEIGHT_SIZE-1:0] Wgt_8_362;input [WEIGHT_SIZE-1:0] Wgt_8_363;input [WEIGHT_SIZE-1:0] Wgt_8_364;input [WEIGHT_SIZE-1:0] Wgt_8_365;input [WEIGHT_SIZE-1:0] Wgt_8_366;input [WEIGHT_SIZE-1:0] Wgt_8_367;input [WEIGHT_SIZE-1:0] Wgt_8_368;input [WEIGHT_SIZE-1:0] Wgt_8_369;input [WEIGHT_SIZE-1:0] Wgt_8_370;input [WEIGHT_SIZE-1:0] Wgt_8_371;input [WEIGHT_SIZE-1:0] Wgt_8_372;input [WEIGHT_SIZE-1:0] Wgt_8_373;input [WEIGHT_SIZE-1:0] Wgt_8_374;input [WEIGHT_SIZE-1:0] Wgt_8_375;input [WEIGHT_SIZE-1:0] Wgt_8_376;input [WEIGHT_SIZE-1:0] Wgt_8_377;input [WEIGHT_SIZE-1:0] Wgt_8_378;input [WEIGHT_SIZE-1:0] Wgt_8_379;input [WEIGHT_SIZE-1:0] Wgt_8_380;input [WEIGHT_SIZE-1:0] Wgt_8_381;input [WEIGHT_SIZE-1:0] Wgt_8_382;input [WEIGHT_SIZE-1:0] Wgt_8_383;input [WEIGHT_SIZE-1:0] Wgt_8_384;input [WEIGHT_SIZE-1:0] Wgt_8_385;input [WEIGHT_SIZE-1:0] Wgt_8_386;input [WEIGHT_SIZE-1:0] Wgt_8_387;input [WEIGHT_SIZE-1:0] Wgt_8_388;input [WEIGHT_SIZE-1:0] Wgt_8_389;input [WEIGHT_SIZE-1:0] Wgt_8_390;input [WEIGHT_SIZE-1:0] Wgt_8_391;input [WEIGHT_SIZE-1:0] Wgt_8_392;input [WEIGHT_SIZE-1:0] Wgt_8_393;input [WEIGHT_SIZE-1:0] Wgt_8_394;input [WEIGHT_SIZE-1:0] Wgt_8_395;input [WEIGHT_SIZE-1:0] Wgt_8_396;input [WEIGHT_SIZE-1:0] Wgt_8_397;input [WEIGHT_SIZE-1:0] Wgt_8_398;input [WEIGHT_SIZE-1:0] Wgt_8_399;input [WEIGHT_SIZE-1:0] Wgt_8_400;input [WEIGHT_SIZE-1:0] Wgt_8_401;input [WEIGHT_SIZE-1:0] Wgt_8_402;input [WEIGHT_SIZE-1:0] Wgt_8_403;input [WEIGHT_SIZE-1:0] Wgt_8_404;input [WEIGHT_SIZE-1:0] Wgt_8_405;input [WEIGHT_SIZE-1:0] Wgt_8_406;input [WEIGHT_SIZE-1:0] Wgt_8_407;input [WEIGHT_SIZE-1:0] Wgt_8_408;input [WEIGHT_SIZE-1:0] Wgt_8_409;input [WEIGHT_SIZE-1:0] Wgt_8_410;input [WEIGHT_SIZE-1:0] Wgt_8_411;input [WEIGHT_SIZE-1:0] Wgt_8_412;input [WEIGHT_SIZE-1:0] Wgt_8_413;input [WEIGHT_SIZE-1:0] Wgt_8_414;input [WEIGHT_SIZE-1:0] Wgt_8_415;input [WEIGHT_SIZE-1:0] Wgt_8_416;input [WEIGHT_SIZE-1:0] Wgt_8_417;input [WEIGHT_SIZE-1:0] Wgt_8_418;input [WEIGHT_SIZE-1:0] Wgt_8_419;input [WEIGHT_SIZE-1:0] Wgt_8_420;input [WEIGHT_SIZE-1:0] Wgt_8_421;input [WEIGHT_SIZE-1:0] Wgt_8_422;input [WEIGHT_SIZE-1:0] Wgt_8_423;input [WEIGHT_SIZE-1:0] Wgt_8_424;input [WEIGHT_SIZE-1:0] Wgt_8_425;input [WEIGHT_SIZE-1:0] Wgt_8_426;input [WEIGHT_SIZE-1:0] Wgt_8_427;input [WEIGHT_SIZE-1:0] Wgt_8_428;input [WEIGHT_SIZE-1:0] Wgt_8_429;input [WEIGHT_SIZE-1:0] Wgt_8_430;input [WEIGHT_SIZE-1:0] Wgt_8_431;input [WEIGHT_SIZE-1:0] Wgt_8_432;input [WEIGHT_SIZE-1:0] Wgt_8_433;input [WEIGHT_SIZE-1:0] Wgt_8_434;input [WEIGHT_SIZE-1:0] Wgt_8_435;input [WEIGHT_SIZE-1:0] Wgt_8_436;input [WEIGHT_SIZE-1:0] Wgt_8_437;input [WEIGHT_SIZE-1:0] Wgt_8_438;input [WEIGHT_SIZE-1:0] Wgt_8_439;input [WEIGHT_SIZE-1:0] Wgt_8_440;input [WEIGHT_SIZE-1:0] Wgt_8_441;input [WEIGHT_SIZE-1:0] Wgt_8_442;input [WEIGHT_SIZE-1:0] Wgt_8_443;input [WEIGHT_SIZE-1:0] Wgt_8_444;input [WEIGHT_SIZE-1:0] Wgt_8_445;input [WEIGHT_SIZE-1:0] Wgt_8_446;input [WEIGHT_SIZE-1:0] Wgt_8_447;input [WEIGHT_SIZE-1:0] Wgt_8_448;input [WEIGHT_SIZE-1:0] Wgt_8_449;input [WEIGHT_SIZE-1:0] Wgt_8_450;input [WEIGHT_SIZE-1:0] Wgt_8_451;input [WEIGHT_SIZE-1:0] Wgt_8_452;input [WEIGHT_SIZE-1:0] Wgt_8_453;input [WEIGHT_SIZE-1:0] Wgt_8_454;input [WEIGHT_SIZE-1:0] Wgt_8_455;input [WEIGHT_SIZE-1:0] Wgt_8_456;input [WEIGHT_SIZE-1:0] Wgt_8_457;input [WEIGHT_SIZE-1:0] Wgt_8_458;input [WEIGHT_SIZE-1:0] Wgt_8_459;input [WEIGHT_SIZE-1:0] Wgt_8_460;input [WEIGHT_SIZE-1:0] Wgt_8_461;input [WEIGHT_SIZE-1:0] Wgt_8_462;input [WEIGHT_SIZE-1:0] Wgt_8_463;input [WEIGHT_SIZE-1:0] Wgt_8_464;input [WEIGHT_SIZE-1:0] Wgt_8_465;input [WEIGHT_SIZE-1:0] Wgt_8_466;input [WEIGHT_SIZE-1:0] Wgt_8_467;input [WEIGHT_SIZE-1:0] Wgt_8_468;input [WEIGHT_SIZE-1:0] Wgt_8_469;input [WEIGHT_SIZE-1:0] Wgt_8_470;input [WEIGHT_SIZE-1:0] Wgt_8_471;input [WEIGHT_SIZE-1:0] Wgt_8_472;input [WEIGHT_SIZE-1:0] Wgt_8_473;input [WEIGHT_SIZE-1:0] Wgt_8_474;input [WEIGHT_SIZE-1:0] Wgt_8_475;input [WEIGHT_SIZE-1:0] Wgt_8_476;input [WEIGHT_SIZE-1:0] Wgt_8_477;input [WEIGHT_SIZE-1:0] Wgt_8_478;input [WEIGHT_SIZE-1:0] Wgt_8_479;input [WEIGHT_SIZE-1:0] Wgt_8_480;input [WEIGHT_SIZE-1:0] Wgt_8_481;input [WEIGHT_SIZE-1:0] Wgt_8_482;input [WEIGHT_SIZE-1:0] Wgt_8_483;input [WEIGHT_SIZE-1:0] Wgt_8_484;input [WEIGHT_SIZE-1:0] Wgt_8_485;input [WEIGHT_SIZE-1:0] Wgt_8_486;input [WEIGHT_SIZE-1:0] Wgt_8_487;input [WEIGHT_SIZE-1:0] Wgt_8_488;input [WEIGHT_SIZE-1:0] Wgt_8_489;input [WEIGHT_SIZE-1:0] Wgt_8_490;input [WEIGHT_SIZE-1:0] Wgt_8_491;input [WEIGHT_SIZE-1:0] Wgt_8_492;input [WEIGHT_SIZE-1:0] Wgt_8_493;input [WEIGHT_SIZE-1:0] Wgt_8_494;input [WEIGHT_SIZE-1:0] Wgt_8_495;input [WEIGHT_SIZE-1:0] Wgt_8_496;input [WEIGHT_SIZE-1:0] Wgt_8_497;input [WEIGHT_SIZE-1:0] Wgt_8_498;input [WEIGHT_SIZE-1:0] Wgt_8_499;input [WEIGHT_SIZE-1:0] Wgt_8_500;input [WEIGHT_SIZE-1:0] Wgt_8_501;input [WEIGHT_SIZE-1:0] Wgt_8_502;input [WEIGHT_SIZE-1:0] Wgt_8_503;input [WEIGHT_SIZE-1:0] Wgt_8_504;input [WEIGHT_SIZE-1:0] Wgt_8_505;input [WEIGHT_SIZE-1:0] Wgt_8_506;input [WEIGHT_SIZE-1:0] Wgt_8_507;input [WEIGHT_SIZE-1:0] Wgt_8_508;input [WEIGHT_SIZE-1:0] Wgt_8_509;input [WEIGHT_SIZE-1:0] Wgt_8_510;input [WEIGHT_SIZE-1:0] Wgt_8_511;input [WEIGHT_SIZE-1:0] Wgt_8_512;input [WEIGHT_SIZE-1:0] Wgt_8_513;input [WEIGHT_SIZE-1:0] Wgt_8_514;input [WEIGHT_SIZE-1:0] Wgt_8_515;input [WEIGHT_SIZE-1:0] Wgt_8_516;input [WEIGHT_SIZE-1:0] Wgt_8_517;input [WEIGHT_SIZE-1:0] Wgt_8_518;input [WEIGHT_SIZE-1:0] Wgt_8_519;input [WEIGHT_SIZE-1:0] Wgt_8_520;input [WEIGHT_SIZE-1:0] Wgt_8_521;input [WEIGHT_SIZE-1:0] Wgt_8_522;input [WEIGHT_SIZE-1:0] Wgt_8_523;input [WEIGHT_SIZE-1:0] Wgt_8_524;input [WEIGHT_SIZE-1:0] Wgt_8_525;input [WEIGHT_SIZE-1:0] Wgt_8_526;input [WEIGHT_SIZE-1:0] Wgt_8_527;input [WEIGHT_SIZE-1:0] Wgt_8_528;input [WEIGHT_SIZE-1:0] Wgt_8_529;input [WEIGHT_SIZE-1:0] Wgt_8_530;input [WEIGHT_SIZE-1:0] Wgt_8_531;input [WEIGHT_SIZE-1:0] Wgt_8_532;input [WEIGHT_SIZE-1:0] Wgt_8_533;input [WEIGHT_SIZE-1:0] Wgt_8_534;input [WEIGHT_SIZE-1:0] Wgt_8_535;input [WEIGHT_SIZE-1:0] Wgt_8_536;input [WEIGHT_SIZE-1:0] Wgt_8_537;input [WEIGHT_SIZE-1:0] Wgt_8_538;input [WEIGHT_SIZE-1:0] Wgt_8_539;input [WEIGHT_SIZE-1:0] Wgt_8_540;input [WEIGHT_SIZE-1:0] Wgt_8_541;input [WEIGHT_SIZE-1:0] Wgt_8_542;input [WEIGHT_SIZE-1:0] Wgt_8_543;input [WEIGHT_SIZE-1:0] Wgt_8_544;input [WEIGHT_SIZE-1:0] Wgt_8_545;input [WEIGHT_SIZE-1:0] Wgt_8_546;input [WEIGHT_SIZE-1:0] Wgt_8_547;input [WEIGHT_SIZE-1:0] Wgt_8_548;input [WEIGHT_SIZE-1:0] Wgt_8_549;input [WEIGHT_SIZE-1:0] Wgt_8_550;input [WEIGHT_SIZE-1:0] Wgt_8_551;input [WEIGHT_SIZE-1:0] Wgt_8_552;input [WEIGHT_SIZE-1:0] Wgt_8_553;input [WEIGHT_SIZE-1:0] Wgt_8_554;input [WEIGHT_SIZE-1:0] Wgt_8_555;input [WEIGHT_SIZE-1:0] Wgt_8_556;input [WEIGHT_SIZE-1:0] Wgt_8_557;input [WEIGHT_SIZE-1:0] Wgt_8_558;input [WEIGHT_SIZE-1:0] Wgt_8_559;input [WEIGHT_SIZE-1:0] Wgt_8_560;input [WEIGHT_SIZE-1:0] Wgt_8_561;input [WEIGHT_SIZE-1:0] Wgt_8_562;input [WEIGHT_SIZE-1:0] Wgt_8_563;input [WEIGHT_SIZE-1:0] Wgt_8_564;input [WEIGHT_SIZE-1:0] Wgt_8_565;input [WEIGHT_SIZE-1:0] Wgt_8_566;input [WEIGHT_SIZE-1:0] Wgt_8_567;input [WEIGHT_SIZE-1:0] Wgt_8_568;input [WEIGHT_SIZE-1:0] Wgt_8_569;input [WEIGHT_SIZE-1:0] Wgt_8_570;input [WEIGHT_SIZE-1:0] Wgt_8_571;input [WEIGHT_SIZE-1:0] Wgt_8_572;input [WEIGHT_SIZE-1:0] Wgt_8_573;input [WEIGHT_SIZE-1:0] Wgt_8_574;input [WEIGHT_SIZE-1:0] Wgt_8_575;input [WEIGHT_SIZE-1:0] Wgt_8_576;input [WEIGHT_SIZE-1:0] Wgt_8_577;input [WEIGHT_SIZE-1:0] Wgt_8_578;input [WEIGHT_SIZE-1:0] Wgt_8_579;input [WEIGHT_SIZE-1:0] Wgt_8_580;input [WEIGHT_SIZE-1:0] Wgt_8_581;input [WEIGHT_SIZE-1:0] Wgt_8_582;input [WEIGHT_SIZE-1:0] Wgt_8_583;input [WEIGHT_SIZE-1:0] Wgt_8_584;input [WEIGHT_SIZE-1:0] Wgt_8_585;input [WEIGHT_SIZE-1:0] Wgt_8_586;input [WEIGHT_SIZE-1:0] Wgt_8_587;input [WEIGHT_SIZE-1:0] Wgt_8_588;input [WEIGHT_SIZE-1:0] Wgt_8_589;input [WEIGHT_SIZE-1:0] Wgt_8_590;input [WEIGHT_SIZE-1:0] Wgt_8_591;input [WEIGHT_SIZE-1:0] Wgt_8_592;input [WEIGHT_SIZE-1:0] Wgt_8_593;input [WEIGHT_SIZE-1:0] Wgt_8_594;input [WEIGHT_SIZE-1:0] Wgt_8_595;input [WEIGHT_SIZE-1:0] Wgt_8_596;input [WEIGHT_SIZE-1:0] Wgt_8_597;input [WEIGHT_SIZE-1:0] Wgt_8_598;input [WEIGHT_SIZE-1:0] Wgt_8_599;input [WEIGHT_SIZE-1:0] Wgt_8_600;input [WEIGHT_SIZE-1:0] Wgt_8_601;input [WEIGHT_SIZE-1:0] Wgt_8_602;input [WEIGHT_SIZE-1:0] Wgt_8_603;input [WEIGHT_SIZE-1:0] Wgt_8_604;input [WEIGHT_SIZE-1:0] Wgt_8_605;input [WEIGHT_SIZE-1:0] Wgt_8_606;input [WEIGHT_SIZE-1:0] Wgt_8_607;input [WEIGHT_SIZE-1:0] Wgt_8_608;input [WEIGHT_SIZE-1:0] Wgt_8_609;input [WEIGHT_SIZE-1:0] Wgt_8_610;input [WEIGHT_SIZE-1:0] Wgt_8_611;input [WEIGHT_SIZE-1:0] Wgt_8_612;input [WEIGHT_SIZE-1:0] Wgt_8_613;input [WEIGHT_SIZE-1:0] Wgt_8_614;input [WEIGHT_SIZE-1:0] Wgt_8_615;input [WEIGHT_SIZE-1:0] Wgt_8_616;input [WEIGHT_SIZE-1:0] Wgt_8_617;input [WEIGHT_SIZE-1:0] Wgt_8_618;input [WEIGHT_SIZE-1:0] Wgt_8_619;input [WEIGHT_SIZE-1:0] Wgt_8_620;input [WEIGHT_SIZE-1:0] Wgt_8_621;input [WEIGHT_SIZE-1:0] Wgt_8_622;input [WEIGHT_SIZE-1:0] Wgt_8_623;input [WEIGHT_SIZE-1:0] Wgt_8_624;input [WEIGHT_SIZE-1:0] Wgt_8_625;input [WEIGHT_SIZE-1:0] Wgt_8_626;input [WEIGHT_SIZE-1:0] Wgt_8_627;input [WEIGHT_SIZE-1:0] Wgt_8_628;input [WEIGHT_SIZE-1:0] Wgt_8_629;input [WEIGHT_SIZE-1:0] Wgt_8_630;input [WEIGHT_SIZE-1:0] Wgt_8_631;input [WEIGHT_SIZE-1:0] Wgt_8_632;input [WEIGHT_SIZE-1:0] Wgt_8_633;input [WEIGHT_SIZE-1:0] Wgt_8_634;input [WEIGHT_SIZE-1:0] Wgt_8_635;input [WEIGHT_SIZE-1:0] Wgt_8_636;input [WEIGHT_SIZE-1:0] Wgt_8_637;input [WEIGHT_SIZE-1:0] Wgt_8_638;input [WEIGHT_SIZE-1:0] Wgt_8_639;input [WEIGHT_SIZE-1:0] Wgt_8_640;input [WEIGHT_SIZE-1:0] Wgt_8_641;input [WEIGHT_SIZE-1:0] Wgt_8_642;input [WEIGHT_SIZE-1:0] Wgt_8_643;input [WEIGHT_SIZE-1:0] Wgt_8_644;input [WEIGHT_SIZE-1:0] Wgt_8_645;input [WEIGHT_SIZE-1:0] Wgt_8_646;input [WEIGHT_SIZE-1:0] Wgt_8_647;input [WEIGHT_SIZE-1:0] Wgt_8_648;input [WEIGHT_SIZE-1:0] Wgt_8_649;input [WEIGHT_SIZE-1:0] Wgt_8_650;input [WEIGHT_SIZE-1:0] Wgt_8_651;input [WEIGHT_SIZE-1:0] Wgt_8_652;input [WEIGHT_SIZE-1:0] Wgt_8_653;input [WEIGHT_SIZE-1:0] Wgt_8_654;input [WEIGHT_SIZE-1:0] Wgt_8_655;input [WEIGHT_SIZE-1:0] Wgt_8_656;input [WEIGHT_SIZE-1:0] Wgt_8_657;input [WEIGHT_SIZE-1:0] Wgt_8_658;input [WEIGHT_SIZE-1:0] Wgt_8_659;input [WEIGHT_SIZE-1:0] Wgt_8_660;input [WEIGHT_SIZE-1:0] Wgt_8_661;input [WEIGHT_SIZE-1:0] Wgt_8_662;input [WEIGHT_SIZE-1:0] Wgt_8_663;input [WEIGHT_SIZE-1:0] Wgt_8_664;input [WEIGHT_SIZE-1:0] Wgt_8_665;input [WEIGHT_SIZE-1:0] Wgt_8_666;input [WEIGHT_SIZE-1:0] Wgt_8_667;input [WEIGHT_SIZE-1:0] Wgt_8_668;input [WEIGHT_SIZE-1:0] Wgt_8_669;input [WEIGHT_SIZE-1:0] Wgt_8_670;input [WEIGHT_SIZE-1:0] Wgt_8_671;input [WEIGHT_SIZE-1:0] Wgt_8_672;input [WEIGHT_SIZE-1:0] Wgt_8_673;input [WEIGHT_SIZE-1:0] Wgt_8_674;input [WEIGHT_SIZE-1:0] Wgt_8_675;input [WEIGHT_SIZE-1:0] Wgt_8_676;input [WEIGHT_SIZE-1:0] Wgt_8_677;input [WEIGHT_SIZE-1:0] Wgt_8_678;input [WEIGHT_SIZE-1:0] Wgt_8_679;input [WEIGHT_SIZE-1:0] Wgt_8_680;input [WEIGHT_SIZE-1:0] Wgt_8_681;input [WEIGHT_SIZE-1:0] Wgt_8_682;input [WEIGHT_SIZE-1:0] Wgt_8_683;input [WEIGHT_SIZE-1:0] Wgt_8_684;input [WEIGHT_SIZE-1:0] Wgt_8_685;input [WEIGHT_SIZE-1:0] Wgt_8_686;input [WEIGHT_SIZE-1:0] Wgt_8_687;input [WEIGHT_SIZE-1:0] Wgt_8_688;input [WEIGHT_SIZE-1:0] Wgt_8_689;input [WEIGHT_SIZE-1:0] Wgt_8_690;input [WEIGHT_SIZE-1:0] Wgt_8_691;input [WEIGHT_SIZE-1:0] Wgt_8_692;input [WEIGHT_SIZE-1:0] Wgt_8_693;input [WEIGHT_SIZE-1:0] Wgt_8_694;input [WEIGHT_SIZE-1:0] Wgt_8_695;input [WEIGHT_SIZE-1:0] Wgt_8_696;input [WEIGHT_SIZE-1:0] Wgt_8_697;input [WEIGHT_SIZE-1:0] Wgt_8_698;input [WEIGHT_SIZE-1:0] Wgt_8_699;input [WEIGHT_SIZE-1:0] Wgt_8_700;input [WEIGHT_SIZE-1:0] Wgt_8_701;input [WEIGHT_SIZE-1:0] Wgt_8_702;input [WEIGHT_SIZE-1:0] Wgt_8_703;input [WEIGHT_SIZE-1:0] Wgt_8_704;input [WEIGHT_SIZE-1:0] Wgt_8_705;input [WEIGHT_SIZE-1:0] Wgt_8_706;input [WEIGHT_SIZE-1:0] Wgt_8_707;input [WEIGHT_SIZE-1:0] Wgt_8_708;input [WEIGHT_SIZE-1:0] Wgt_8_709;input [WEIGHT_SIZE-1:0] Wgt_8_710;input [WEIGHT_SIZE-1:0] Wgt_8_711;input [WEIGHT_SIZE-1:0] Wgt_8_712;input [WEIGHT_SIZE-1:0] Wgt_8_713;input [WEIGHT_SIZE-1:0] Wgt_8_714;input [WEIGHT_SIZE-1:0] Wgt_8_715;input [WEIGHT_SIZE-1:0] Wgt_8_716;input [WEIGHT_SIZE-1:0] Wgt_8_717;input [WEIGHT_SIZE-1:0] Wgt_8_718;input [WEIGHT_SIZE-1:0] Wgt_8_719;input [WEIGHT_SIZE-1:0] Wgt_8_720;input [WEIGHT_SIZE-1:0] Wgt_8_721;input [WEIGHT_SIZE-1:0] Wgt_8_722;input [WEIGHT_SIZE-1:0] Wgt_8_723;input [WEIGHT_SIZE-1:0] Wgt_8_724;input [WEIGHT_SIZE-1:0] Wgt_8_725;input [WEIGHT_SIZE-1:0] Wgt_8_726;input [WEIGHT_SIZE-1:0] Wgt_8_727;input [WEIGHT_SIZE-1:0] Wgt_8_728;input [WEIGHT_SIZE-1:0] Wgt_8_729;input [WEIGHT_SIZE-1:0] Wgt_8_730;input [WEIGHT_SIZE-1:0] Wgt_8_731;input [WEIGHT_SIZE-1:0] Wgt_8_732;input [WEIGHT_SIZE-1:0] Wgt_8_733;input [WEIGHT_SIZE-1:0] Wgt_8_734;input [WEIGHT_SIZE-1:0] Wgt_8_735;input [WEIGHT_SIZE-1:0] Wgt_8_736;input [WEIGHT_SIZE-1:0] Wgt_8_737;input [WEIGHT_SIZE-1:0] Wgt_8_738;input [WEIGHT_SIZE-1:0] Wgt_8_739;input [WEIGHT_SIZE-1:0] Wgt_8_740;input [WEIGHT_SIZE-1:0] Wgt_8_741;input [WEIGHT_SIZE-1:0] Wgt_8_742;input [WEIGHT_SIZE-1:0] Wgt_8_743;input [WEIGHT_SIZE-1:0] Wgt_8_744;input [WEIGHT_SIZE-1:0] Wgt_8_745;input [WEIGHT_SIZE-1:0] Wgt_8_746;input [WEIGHT_SIZE-1:0] Wgt_8_747;input [WEIGHT_SIZE-1:0] Wgt_8_748;input [WEIGHT_SIZE-1:0] Wgt_8_749;input [WEIGHT_SIZE-1:0] Wgt_8_750;input [WEIGHT_SIZE-1:0] Wgt_8_751;input [WEIGHT_SIZE-1:0] Wgt_8_752;input [WEIGHT_SIZE-1:0] Wgt_8_753;input [WEIGHT_SIZE-1:0] Wgt_8_754;input [WEIGHT_SIZE-1:0] Wgt_8_755;input [WEIGHT_SIZE-1:0] Wgt_8_756;input [WEIGHT_SIZE-1:0] Wgt_8_757;input [WEIGHT_SIZE-1:0] Wgt_8_758;input [WEIGHT_SIZE-1:0] Wgt_8_759;input [WEIGHT_SIZE-1:0] Wgt_8_760;input [WEIGHT_SIZE-1:0] Wgt_8_761;input [WEIGHT_SIZE-1:0] Wgt_8_762;input [WEIGHT_SIZE-1:0] Wgt_8_763;input [WEIGHT_SIZE-1:0] Wgt_8_764;input [WEIGHT_SIZE-1:0] Wgt_8_765;input [WEIGHT_SIZE-1:0] Wgt_8_766;input [WEIGHT_SIZE-1:0] Wgt_8_767;input [WEIGHT_SIZE-1:0] Wgt_8_768;input [WEIGHT_SIZE-1:0] Wgt_8_769;input [WEIGHT_SIZE-1:0] Wgt_8_770;input [WEIGHT_SIZE-1:0] Wgt_8_771;input [WEIGHT_SIZE-1:0] Wgt_8_772;input [WEIGHT_SIZE-1:0] Wgt_8_773;input [WEIGHT_SIZE-1:0] Wgt_8_774;input [WEIGHT_SIZE-1:0] Wgt_8_775;input [WEIGHT_SIZE-1:0] Wgt_8_776;input [WEIGHT_SIZE-1:0] Wgt_8_777;input [WEIGHT_SIZE-1:0] Wgt_8_778;input [WEIGHT_SIZE-1:0] Wgt_8_779;input [WEIGHT_SIZE-1:0] Wgt_8_780;input [WEIGHT_SIZE-1:0] Wgt_8_781;input [WEIGHT_SIZE-1:0] Wgt_8_782;input [WEIGHT_SIZE-1:0] Wgt_8_783;input [WEIGHT_SIZE-1:0] Wgt_8_784;input [WEIGHT_SIZE-1:0] Wgt_9_0;input [WEIGHT_SIZE-1:0] Wgt_9_1;input [WEIGHT_SIZE-1:0] Wgt_9_2;input [WEIGHT_SIZE-1:0] Wgt_9_3;input [WEIGHT_SIZE-1:0] Wgt_9_4;input [WEIGHT_SIZE-1:0] Wgt_9_5;input [WEIGHT_SIZE-1:0] Wgt_9_6;input [WEIGHT_SIZE-1:0] Wgt_9_7;input [WEIGHT_SIZE-1:0] Wgt_9_8;input [WEIGHT_SIZE-1:0] Wgt_9_9;input [WEIGHT_SIZE-1:0] Wgt_9_10;input [WEIGHT_SIZE-1:0] Wgt_9_11;input [WEIGHT_SIZE-1:0] Wgt_9_12;input [WEIGHT_SIZE-1:0] Wgt_9_13;input [WEIGHT_SIZE-1:0] Wgt_9_14;input [WEIGHT_SIZE-1:0] Wgt_9_15;input [WEIGHT_SIZE-1:0] Wgt_9_16;input [WEIGHT_SIZE-1:0] Wgt_9_17;input [WEIGHT_SIZE-1:0] Wgt_9_18;input [WEIGHT_SIZE-1:0] Wgt_9_19;input [WEIGHT_SIZE-1:0] Wgt_9_20;input [WEIGHT_SIZE-1:0] Wgt_9_21;input [WEIGHT_SIZE-1:0] Wgt_9_22;input [WEIGHT_SIZE-1:0] Wgt_9_23;input [WEIGHT_SIZE-1:0] Wgt_9_24;input [WEIGHT_SIZE-1:0] Wgt_9_25;input [WEIGHT_SIZE-1:0] Wgt_9_26;input [WEIGHT_SIZE-1:0] Wgt_9_27;input [WEIGHT_SIZE-1:0] Wgt_9_28;input [WEIGHT_SIZE-1:0] Wgt_9_29;input [WEIGHT_SIZE-1:0] Wgt_9_30;input [WEIGHT_SIZE-1:0] Wgt_9_31;input [WEIGHT_SIZE-1:0] Wgt_9_32;input [WEIGHT_SIZE-1:0] Wgt_9_33;input [WEIGHT_SIZE-1:0] Wgt_9_34;input [WEIGHT_SIZE-1:0] Wgt_9_35;input [WEIGHT_SIZE-1:0] Wgt_9_36;input [WEIGHT_SIZE-1:0] Wgt_9_37;input [WEIGHT_SIZE-1:0] Wgt_9_38;input [WEIGHT_SIZE-1:0] Wgt_9_39;input [WEIGHT_SIZE-1:0] Wgt_9_40;input [WEIGHT_SIZE-1:0] Wgt_9_41;input [WEIGHT_SIZE-1:0] Wgt_9_42;input [WEIGHT_SIZE-1:0] Wgt_9_43;input [WEIGHT_SIZE-1:0] Wgt_9_44;input [WEIGHT_SIZE-1:0] Wgt_9_45;input [WEIGHT_SIZE-1:0] Wgt_9_46;input [WEIGHT_SIZE-1:0] Wgt_9_47;input [WEIGHT_SIZE-1:0] Wgt_9_48;input [WEIGHT_SIZE-1:0] Wgt_9_49;input [WEIGHT_SIZE-1:0] Wgt_9_50;input [WEIGHT_SIZE-1:0] Wgt_9_51;input [WEIGHT_SIZE-1:0] Wgt_9_52;input [WEIGHT_SIZE-1:0] Wgt_9_53;input [WEIGHT_SIZE-1:0] Wgt_9_54;input [WEIGHT_SIZE-1:0] Wgt_9_55;input [WEIGHT_SIZE-1:0] Wgt_9_56;input [WEIGHT_SIZE-1:0] Wgt_9_57;input [WEIGHT_SIZE-1:0] Wgt_9_58;input [WEIGHT_SIZE-1:0] Wgt_9_59;input [WEIGHT_SIZE-1:0] Wgt_9_60;input [WEIGHT_SIZE-1:0] Wgt_9_61;input [WEIGHT_SIZE-1:0] Wgt_9_62;input [WEIGHT_SIZE-1:0] Wgt_9_63;input [WEIGHT_SIZE-1:0] Wgt_9_64;input [WEIGHT_SIZE-1:0] Wgt_9_65;input [WEIGHT_SIZE-1:0] Wgt_9_66;input [WEIGHT_SIZE-1:0] Wgt_9_67;input [WEIGHT_SIZE-1:0] Wgt_9_68;input [WEIGHT_SIZE-1:0] Wgt_9_69;input [WEIGHT_SIZE-1:0] Wgt_9_70;input [WEIGHT_SIZE-1:0] Wgt_9_71;input [WEIGHT_SIZE-1:0] Wgt_9_72;input [WEIGHT_SIZE-1:0] Wgt_9_73;input [WEIGHT_SIZE-1:0] Wgt_9_74;input [WEIGHT_SIZE-1:0] Wgt_9_75;input [WEIGHT_SIZE-1:0] Wgt_9_76;input [WEIGHT_SIZE-1:0] Wgt_9_77;input [WEIGHT_SIZE-1:0] Wgt_9_78;input [WEIGHT_SIZE-1:0] Wgt_9_79;input [WEIGHT_SIZE-1:0] Wgt_9_80;input [WEIGHT_SIZE-1:0] Wgt_9_81;input [WEIGHT_SIZE-1:0] Wgt_9_82;input [WEIGHT_SIZE-1:0] Wgt_9_83;input [WEIGHT_SIZE-1:0] Wgt_9_84;input [WEIGHT_SIZE-1:0] Wgt_9_85;input [WEIGHT_SIZE-1:0] Wgt_9_86;input [WEIGHT_SIZE-1:0] Wgt_9_87;input [WEIGHT_SIZE-1:0] Wgt_9_88;input [WEIGHT_SIZE-1:0] Wgt_9_89;input [WEIGHT_SIZE-1:0] Wgt_9_90;input [WEIGHT_SIZE-1:0] Wgt_9_91;input [WEIGHT_SIZE-1:0] Wgt_9_92;input [WEIGHT_SIZE-1:0] Wgt_9_93;input [WEIGHT_SIZE-1:0] Wgt_9_94;input [WEIGHT_SIZE-1:0] Wgt_9_95;input [WEIGHT_SIZE-1:0] Wgt_9_96;input [WEIGHT_SIZE-1:0] Wgt_9_97;input [WEIGHT_SIZE-1:0] Wgt_9_98;input [WEIGHT_SIZE-1:0] Wgt_9_99;input [WEIGHT_SIZE-1:0] Wgt_9_100;input [WEIGHT_SIZE-1:0] Wgt_9_101;input [WEIGHT_SIZE-1:0] Wgt_9_102;input [WEIGHT_SIZE-1:0] Wgt_9_103;input [WEIGHT_SIZE-1:0] Wgt_9_104;input [WEIGHT_SIZE-1:0] Wgt_9_105;input [WEIGHT_SIZE-1:0] Wgt_9_106;input [WEIGHT_SIZE-1:0] Wgt_9_107;input [WEIGHT_SIZE-1:0] Wgt_9_108;input [WEIGHT_SIZE-1:0] Wgt_9_109;input [WEIGHT_SIZE-1:0] Wgt_9_110;input [WEIGHT_SIZE-1:0] Wgt_9_111;input [WEIGHT_SIZE-1:0] Wgt_9_112;input [WEIGHT_SIZE-1:0] Wgt_9_113;input [WEIGHT_SIZE-1:0] Wgt_9_114;input [WEIGHT_SIZE-1:0] Wgt_9_115;input [WEIGHT_SIZE-1:0] Wgt_9_116;input [WEIGHT_SIZE-1:0] Wgt_9_117;input [WEIGHT_SIZE-1:0] Wgt_9_118;input [WEIGHT_SIZE-1:0] Wgt_9_119;input [WEIGHT_SIZE-1:0] Wgt_9_120;input [WEIGHT_SIZE-1:0] Wgt_9_121;input [WEIGHT_SIZE-1:0] Wgt_9_122;input [WEIGHT_SIZE-1:0] Wgt_9_123;input [WEIGHT_SIZE-1:0] Wgt_9_124;input [WEIGHT_SIZE-1:0] Wgt_9_125;input [WEIGHT_SIZE-1:0] Wgt_9_126;input [WEIGHT_SIZE-1:0] Wgt_9_127;input [WEIGHT_SIZE-1:0] Wgt_9_128;input [WEIGHT_SIZE-1:0] Wgt_9_129;input [WEIGHT_SIZE-1:0] Wgt_9_130;input [WEIGHT_SIZE-1:0] Wgt_9_131;input [WEIGHT_SIZE-1:0] Wgt_9_132;input [WEIGHT_SIZE-1:0] Wgt_9_133;input [WEIGHT_SIZE-1:0] Wgt_9_134;input [WEIGHT_SIZE-1:0] Wgt_9_135;input [WEIGHT_SIZE-1:0] Wgt_9_136;input [WEIGHT_SIZE-1:0] Wgt_9_137;input [WEIGHT_SIZE-1:0] Wgt_9_138;input [WEIGHT_SIZE-1:0] Wgt_9_139;input [WEIGHT_SIZE-1:0] Wgt_9_140;input [WEIGHT_SIZE-1:0] Wgt_9_141;input [WEIGHT_SIZE-1:0] Wgt_9_142;input [WEIGHT_SIZE-1:0] Wgt_9_143;input [WEIGHT_SIZE-1:0] Wgt_9_144;input [WEIGHT_SIZE-1:0] Wgt_9_145;input [WEIGHT_SIZE-1:0] Wgt_9_146;input [WEIGHT_SIZE-1:0] Wgt_9_147;input [WEIGHT_SIZE-1:0] Wgt_9_148;input [WEIGHT_SIZE-1:0] Wgt_9_149;input [WEIGHT_SIZE-1:0] Wgt_9_150;input [WEIGHT_SIZE-1:0] Wgt_9_151;input [WEIGHT_SIZE-1:0] Wgt_9_152;input [WEIGHT_SIZE-1:0] Wgt_9_153;input [WEIGHT_SIZE-1:0] Wgt_9_154;input [WEIGHT_SIZE-1:0] Wgt_9_155;input [WEIGHT_SIZE-1:0] Wgt_9_156;input [WEIGHT_SIZE-1:0] Wgt_9_157;input [WEIGHT_SIZE-1:0] Wgt_9_158;input [WEIGHT_SIZE-1:0] Wgt_9_159;input [WEIGHT_SIZE-1:0] Wgt_9_160;input [WEIGHT_SIZE-1:0] Wgt_9_161;input [WEIGHT_SIZE-1:0] Wgt_9_162;input [WEIGHT_SIZE-1:0] Wgt_9_163;input [WEIGHT_SIZE-1:0] Wgt_9_164;input [WEIGHT_SIZE-1:0] Wgt_9_165;input [WEIGHT_SIZE-1:0] Wgt_9_166;input [WEIGHT_SIZE-1:0] Wgt_9_167;input [WEIGHT_SIZE-1:0] Wgt_9_168;input [WEIGHT_SIZE-1:0] Wgt_9_169;input [WEIGHT_SIZE-1:0] Wgt_9_170;input [WEIGHT_SIZE-1:0] Wgt_9_171;input [WEIGHT_SIZE-1:0] Wgt_9_172;input [WEIGHT_SIZE-1:0] Wgt_9_173;input [WEIGHT_SIZE-1:0] Wgt_9_174;input [WEIGHT_SIZE-1:0] Wgt_9_175;input [WEIGHT_SIZE-1:0] Wgt_9_176;input [WEIGHT_SIZE-1:0] Wgt_9_177;input [WEIGHT_SIZE-1:0] Wgt_9_178;input [WEIGHT_SIZE-1:0] Wgt_9_179;input [WEIGHT_SIZE-1:0] Wgt_9_180;input [WEIGHT_SIZE-1:0] Wgt_9_181;input [WEIGHT_SIZE-1:0] Wgt_9_182;input [WEIGHT_SIZE-1:0] Wgt_9_183;input [WEIGHT_SIZE-1:0] Wgt_9_184;input [WEIGHT_SIZE-1:0] Wgt_9_185;input [WEIGHT_SIZE-1:0] Wgt_9_186;input [WEIGHT_SIZE-1:0] Wgt_9_187;input [WEIGHT_SIZE-1:0] Wgt_9_188;input [WEIGHT_SIZE-1:0] Wgt_9_189;input [WEIGHT_SIZE-1:0] Wgt_9_190;input [WEIGHT_SIZE-1:0] Wgt_9_191;input [WEIGHT_SIZE-1:0] Wgt_9_192;input [WEIGHT_SIZE-1:0] Wgt_9_193;input [WEIGHT_SIZE-1:0] Wgt_9_194;input [WEIGHT_SIZE-1:0] Wgt_9_195;input [WEIGHT_SIZE-1:0] Wgt_9_196;input [WEIGHT_SIZE-1:0] Wgt_9_197;input [WEIGHT_SIZE-1:0] Wgt_9_198;input [WEIGHT_SIZE-1:0] Wgt_9_199;input [WEIGHT_SIZE-1:0] Wgt_9_200;input [WEIGHT_SIZE-1:0] Wgt_9_201;input [WEIGHT_SIZE-1:0] Wgt_9_202;input [WEIGHT_SIZE-1:0] Wgt_9_203;input [WEIGHT_SIZE-1:0] Wgt_9_204;input [WEIGHT_SIZE-1:0] Wgt_9_205;input [WEIGHT_SIZE-1:0] Wgt_9_206;input [WEIGHT_SIZE-1:0] Wgt_9_207;input [WEIGHT_SIZE-1:0] Wgt_9_208;input [WEIGHT_SIZE-1:0] Wgt_9_209;input [WEIGHT_SIZE-1:0] Wgt_9_210;input [WEIGHT_SIZE-1:0] Wgt_9_211;input [WEIGHT_SIZE-1:0] Wgt_9_212;input [WEIGHT_SIZE-1:0] Wgt_9_213;input [WEIGHT_SIZE-1:0] Wgt_9_214;input [WEIGHT_SIZE-1:0] Wgt_9_215;input [WEIGHT_SIZE-1:0] Wgt_9_216;input [WEIGHT_SIZE-1:0] Wgt_9_217;input [WEIGHT_SIZE-1:0] Wgt_9_218;input [WEIGHT_SIZE-1:0] Wgt_9_219;input [WEIGHT_SIZE-1:0] Wgt_9_220;input [WEIGHT_SIZE-1:0] Wgt_9_221;input [WEIGHT_SIZE-1:0] Wgt_9_222;input [WEIGHT_SIZE-1:0] Wgt_9_223;input [WEIGHT_SIZE-1:0] Wgt_9_224;input [WEIGHT_SIZE-1:0] Wgt_9_225;input [WEIGHT_SIZE-1:0] Wgt_9_226;input [WEIGHT_SIZE-1:0] Wgt_9_227;input [WEIGHT_SIZE-1:0] Wgt_9_228;input [WEIGHT_SIZE-1:0] Wgt_9_229;input [WEIGHT_SIZE-1:0] Wgt_9_230;input [WEIGHT_SIZE-1:0] Wgt_9_231;input [WEIGHT_SIZE-1:0] Wgt_9_232;input [WEIGHT_SIZE-1:0] Wgt_9_233;input [WEIGHT_SIZE-1:0] Wgt_9_234;input [WEIGHT_SIZE-1:0] Wgt_9_235;input [WEIGHT_SIZE-1:0] Wgt_9_236;input [WEIGHT_SIZE-1:0] Wgt_9_237;input [WEIGHT_SIZE-1:0] Wgt_9_238;input [WEIGHT_SIZE-1:0] Wgt_9_239;input [WEIGHT_SIZE-1:0] Wgt_9_240;input [WEIGHT_SIZE-1:0] Wgt_9_241;input [WEIGHT_SIZE-1:0] Wgt_9_242;input [WEIGHT_SIZE-1:0] Wgt_9_243;input [WEIGHT_SIZE-1:0] Wgt_9_244;input [WEIGHT_SIZE-1:0] Wgt_9_245;input [WEIGHT_SIZE-1:0] Wgt_9_246;input [WEIGHT_SIZE-1:0] Wgt_9_247;input [WEIGHT_SIZE-1:0] Wgt_9_248;input [WEIGHT_SIZE-1:0] Wgt_9_249;input [WEIGHT_SIZE-1:0] Wgt_9_250;input [WEIGHT_SIZE-1:0] Wgt_9_251;input [WEIGHT_SIZE-1:0] Wgt_9_252;input [WEIGHT_SIZE-1:0] Wgt_9_253;input [WEIGHT_SIZE-1:0] Wgt_9_254;input [WEIGHT_SIZE-1:0] Wgt_9_255;input [WEIGHT_SIZE-1:0] Wgt_9_256;input [WEIGHT_SIZE-1:0] Wgt_9_257;input [WEIGHT_SIZE-1:0] Wgt_9_258;input [WEIGHT_SIZE-1:0] Wgt_9_259;input [WEIGHT_SIZE-1:0] Wgt_9_260;input [WEIGHT_SIZE-1:0] Wgt_9_261;input [WEIGHT_SIZE-1:0] Wgt_9_262;input [WEIGHT_SIZE-1:0] Wgt_9_263;input [WEIGHT_SIZE-1:0] Wgt_9_264;input [WEIGHT_SIZE-1:0] Wgt_9_265;input [WEIGHT_SIZE-1:0] Wgt_9_266;input [WEIGHT_SIZE-1:0] Wgt_9_267;input [WEIGHT_SIZE-1:0] Wgt_9_268;input [WEIGHT_SIZE-1:0] Wgt_9_269;input [WEIGHT_SIZE-1:0] Wgt_9_270;input [WEIGHT_SIZE-1:0] Wgt_9_271;input [WEIGHT_SIZE-1:0] Wgt_9_272;input [WEIGHT_SIZE-1:0] Wgt_9_273;input [WEIGHT_SIZE-1:0] Wgt_9_274;input [WEIGHT_SIZE-1:0] Wgt_9_275;input [WEIGHT_SIZE-1:0] Wgt_9_276;input [WEIGHT_SIZE-1:0] Wgt_9_277;input [WEIGHT_SIZE-1:0] Wgt_9_278;input [WEIGHT_SIZE-1:0] Wgt_9_279;input [WEIGHT_SIZE-1:0] Wgt_9_280;input [WEIGHT_SIZE-1:0] Wgt_9_281;input [WEIGHT_SIZE-1:0] Wgt_9_282;input [WEIGHT_SIZE-1:0] Wgt_9_283;input [WEIGHT_SIZE-1:0] Wgt_9_284;input [WEIGHT_SIZE-1:0] Wgt_9_285;input [WEIGHT_SIZE-1:0] Wgt_9_286;input [WEIGHT_SIZE-1:0] Wgt_9_287;input [WEIGHT_SIZE-1:0] Wgt_9_288;input [WEIGHT_SIZE-1:0] Wgt_9_289;input [WEIGHT_SIZE-1:0] Wgt_9_290;input [WEIGHT_SIZE-1:0] Wgt_9_291;input [WEIGHT_SIZE-1:0] Wgt_9_292;input [WEIGHT_SIZE-1:0] Wgt_9_293;input [WEIGHT_SIZE-1:0] Wgt_9_294;input [WEIGHT_SIZE-1:0] Wgt_9_295;input [WEIGHT_SIZE-1:0] Wgt_9_296;input [WEIGHT_SIZE-1:0] Wgt_9_297;input [WEIGHT_SIZE-1:0] Wgt_9_298;input [WEIGHT_SIZE-1:0] Wgt_9_299;input [WEIGHT_SIZE-1:0] Wgt_9_300;input [WEIGHT_SIZE-1:0] Wgt_9_301;input [WEIGHT_SIZE-1:0] Wgt_9_302;input [WEIGHT_SIZE-1:0] Wgt_9_303;input [WEIGHT_SIZE-1:0] Wgt_9_304;input [WEIGHT_SIZE-1:0] Wgt_9_305;input [WEIGHT_SIZE-1:0] Wgt_9_306;input [WEIGHT_SIZE-1:0] Wgt_9_307;input [WEIGHT_SIZE-1:0] Wgt_9_308;input [WEIGHT_SIZE-1:0] Wgt_9_309;input [WEIGHT_SIZE-1:0] Wgt_9_310;input [WEIGHT_SIZE-1:0] Wgt_9_311;input [WEIGHT_SIZE-1:0] Wgt_9_312;input [WEIGHT_SIZE-1:0] Wgt_9_313;input [WEIGHT_SIZE-1:0] Wgt_9_314;input [WEIGHT_SIZE-1:0] Wgt_9_315;input [WEIGHT_SIZE-1:0] Wgt_9_316;input [WEIGHT_SIZE-1:0] Wgt_9_317;input [WEIGHT_SIZE-1:0] Wgt_9_318;input [WEIGHT_SIZE-1:0] Wgt_9_319;input [WEIGHT_SIZE-1:0] Wgt_9_320;input [WEIGHT_SIZE-1:0] Wgt_9_321;input [WEIGHT_SIZE-1:0] Wgt_9_322;input [WEIGHT_SIZE-1:0] Wgt_9_323;input [WEIGHT_SIZE-1:0] Wgt_9_324;input [WEIGHT_SIZE-1:0] Wgt_9_325;input [WEIGHT_SIZE-1:0] Wgt_9_326;input [WEIGHT_SIZE-1:0] Wgt_9_327;input [WEIGHT_SIZE-1:0] Wgt_9_328;input [WEIGHT_SIZE-1:0] Wgt_9_329;input [WEIGHT_SIZE-1:0] Wgt_9_330;input [WEIGHT_SIZE-1:0] Wgt_9_331;input [WEIGHT_SIZE-1:0] Wgt_9_332;input [WEIGHT_SIZE-1:0] Wgt_9_333;input [WEIGHT_SIZE-1:0] Wgt_9_334;input [WEIGHT_SIZE-1:0] Wgt_9_335;input [WEIGHT_SIZE-1:0] Wgt_9_336;input [WEIGHT_SIZE-1:0] Wgt_9_337;input [WEIGHT_SIZE-1:0] Wgt_9_338;input [WEIGHT_SIZE-1:0] Wgt_9_339;input [WEIGHT_SIZE-1:0] Wgt_9_340;input [WEIGHT_SIZE-1:0] Wgt_9_341;input [WEIGHT_SIZE-1:0] Wgt_9_342;input [WEIGHT_SIZE-1:0] Wgt_9_343;input [WEIGHT_SIZE-1:0] Wgt_9_344;input [WEIGHT_SIZE-1:0] Wgt_9_345;input [WEIGHT_SIZE-1:0] Wgt_9_346;input [WEIGHT_SIZE-1:0] Wgt_9_347;input [WEIGHT_SIZE-1:0] Wgt_9_348;input [WEIGHT_SIZE-1:0] Wgt_9_349;input [WEIGHT_SIZE-1:0] Wgt_9_350;input [WEIGHT_SIZE-1:0] Wgt_9_351;input [WEIGHT_SIZE-1:0] Wgt_9_352;input [WEIGHT_SIZE-1:0] Wgt_9_353;input [WEIGHT_SIZE-1:0] Wgt_9_354;input [WEIGHT_SIZE-1:0] Wgt_9_355;input [WEIGHT_SIZE-1:0] Wgt_9_356;input [WEIGHT_SIZE-1:0] Wgt_9_357;input [WEIGHT_SIZE-1:0] Wgt_9_358;input [WEIGHT_SIZE-1:0] Wgt_9_359;input [WEIGHT_SIZE-1:0] Wgt_9_360;input [WEIGHT_SIZE-1:0] Wgt_9_361;input [WEIGHT_SIZE-1:0] Wgt_9_362;input [WEIGHT_SIZE-1:0] Wgt_9_363;input [WEIGHT_SIZE-1:0] Wgt_9_364;input [WEIGHT_SIZE-1:0] Wgt_9_365;input [WEIGHT_SIZE-1:0] Wgt_9_366;input [WEIGHT_SIZE-1:0] Wgt_9_367;input [WEIGHT_SIZE-1:0] Wgt_9_368;input [WEIGHT_SIZE-1:0] Wgt_9_369;input [WEIGHT_SIZE-1:0] Wgt_9_370;input [WEIGHT_SIZE-1:0] Wgt_9_371;input [WEIGHT_SIZE-1:0] Wgt_9_372;input [WEIGHT_SIZE-1:0] Wgt_9_373;input [WEIGHT_SIZE-1:0] Wgt_9_374;input [WEIGHT_SIZE-1:0] Wgt_9_375;input [WEIGHT_SIZE-1:0] Wgt_9_376;input [WEIGHT_SIZE-1:0] Wgt_9_377;input [WEIGHT_SIZE-1:0] Wgt_9_378;input [WEIGHT_SIZE-1:0] Wgt_9_379;input [WEIGHT_SIZE-1:0] Wgt_9_380;input [WEIGHT_SIZE-1:0] Wgt_9_381;input [WEIGHT_SIZE-1:0] Wgt_9_382;input [WEIGHT_SIZE-1:0] Wgt_9_383;input [WEIGHT_SIZE-1:0] Wgt_9_384;input [WEIGHT_SIZE-1:0] Wgt_9_385;input [WEIGHT_SIZE-1:0] Wgt_9_386;input [WEIGHT_SIZE-1:0] Wgt_9_387;input [WEIGHT_SIZE-1:0] Wgt_9_388;input [WEIGHT_SIZE-1:0] Wgt_9_389;input [WEIGHT_SIZE-1:0] Wgt_9_390;input [WEIGHT_SIZE-1:0] Wgt_9_391;input [WEIGHT_SIZE-1:0] Wgt_9_392;input [WEIGHT_SIZE-1:0] Wgt_9_393;input [WEIGHT_SIZE-1:0] Wgt_9_394;input [WEIGHT_SIZE-1:0] Wgt_9_395;input [WEIGHT_SIZE-1:0] Wgt_9_396;input [WEIGHT_SIZE-1:0] Wgt_9_397;input [WEIGHT_SIZE-1:0] Wgt_9_398;input [WEIGHT_SIZE-1:0] Wgt_9_399;input [WEIGHT_SIZE-1:0] Wgt_9_400;input [WEIGHT_SIZE-1:0] Wgt_9_401;input [WEIGHT_SIZE-1:0] Wgt_9_402;input [WEIGHT_SIZE-1:0] Wgt_9_403;input [WEIGHT_SIZE-1:0] Wgt_9_404;input [WEIGHT_SIZE-1:0] Wgt_9_405;input [WEIGHT_SIZE-1:0] Wgt_9_406;input [WEIGHT_SIZE-1:0] Wgt_9_407;input [WEIGHT_SIZE-1:0] Wgt_9_408;input [WEIGHT_SIZE-1:0] Wgt_9_409;input [WEIGHT_SIZE-1:0] Wgt_9_410;input [WEIGHT_SIZE-1:0] Wgt_9_411;input [WEIGHT_SIZE-1:0] Wgt_9_412;input [WEIGHT_SIZE-1:0] Wgt_9_413;input [WEIGHT_SIZE-1:0] Wgt_9_414;input [WEIGHT_SIZE-1:0] Wgt_9_415;input [WEIGHT_SIZE-1:0] Wgt_9_416;input [WEIGHT_SIZE-1:0] Wgt_9_417;input [WEIGHT_SIZE-1:0] Wgt_9_418;input [WEIGHT_SIZE-1:0] Wgt_9_419;input [WEIGHT_SIZE-1:0] Wgt_9_420;input [WEIGHT_SIZE-1:0] Wgt_9_421;input [WEIGHT_SIZE-1:0] Wgt_9_422;input [WEIGHT_SIZE-1:0] Wgt_9_423;input [WEIGHT_SIZE-1:0] Wgt_9_424;input [WEIGHT_SIZE-1:0] Wgt_9_425;input [WEIGHT_SIZE-1:0] Wgt_9_426;input [WEIGHT_SIZE-1:0] Wgt_9_427;input [WEIGHT_SIZE-1:0] Wgt_9_428;input [WEIGHT_SIZE-1:0] Wgt_9_429;input [WEIGHT_SIZE-1:0] Wgt_9_430;input [WEIGHT_SIZE-1:0] Wgt_9_431;input [WEIGHT_SIZE-1:0] Wgt_9_432;input [WEIGHT_SIZE-1:0] Wgt_9_433;input [WEIGHT_SIZE-1:0] Wgt_9_434;input [WEIGHT_SIZE-1:0] Wgt_9_435;input [WEIGHT_SIZE-1:0] Wgt_9_436;input [WEIGHT_SIZE-1:0] Wgt_9_437;input [WEIGHT_SIZE-1:0] Wgt_9_438;input [WEIGHT_SIZE-1:0] Wgt_9_439;input [WEIGHT_SIZE-1:0] Wgt_9_440;input [WEIGHT_SIZE-1:0] Wgt_9_441;input [WEIGHT_SIZE-1:0] Wgt_9_442;input [WEIGHT_SIZE-1:0] Wgt_9_443;input [WEIGHT_SIZE-1:0] Wgt_9_444;input [WEIGHT_SIZE-1:0] Wgt_9_445;input [WEIGHT_SIZE-1:0] Wgt_9_446;input [WEIGHT_SIZE-1:0] Wgt_9_447;input [WEIGHT_SIZE-1:0] Wgt_9_448;input [WEIGHT_SIZE-1:0] Wgt_9_449;input [WEIGHT_SIZE-1:0] Wgt_9_450;input [WEIGHT_SIZE-1:0] Wgt_9_451;input [WEIGHT_SIZE-1:0] Wgt_9_452;input [WEIGHT_SIZE-1:0] Wgt_9_453;input [WEIGHT_SIZE-1:0] Wgt_9_454;input [WEIGHT_SIZE-1:0] Wgt_9_455;input [WEIGHT_SIZE-1:0] Wgt_9_456;input [WEIGHT_SIZE-1:0] Wgt_9_457;input [WEIGHT_SIZE-1:0] Wgt_9_458;input [WEIGHT_SIZE-1:0] Wgt_9_459;input [WEIGHT_SIZE-1:0] Wgt_9_460;input [WEIGHT_SIZE-1:0] Wgt_9_461;input [WEIGHT_SIZE-1:0] Wgt_9_462;input [WEIGHT_SIZE-1:0] Wgt_9_463;input [WEIGHT_SIZE-1:0] Wgt_9_464;input [WEIGHT_SIZE-1:0] Wgt_9_465;input [WEIGHT_SIZE-1:0] Wgt_9_466;input [WEIGHT_SIZE-1:0] Wgt_9_467;input [WEIGHT_SIZE-1:0] Wgt_9_468;input [WEIGHT_SIZE-1:0] Wgt_9_469;input [WEIGHT_SIZE-1:0] Wgt_9_470;input [WEIGHT_SIZE-1:0] Wgt_9_471;input [WEIGHT_SIZE-1:0] Wgt_9_472;input [WEIGHT_SIZE-1:0] Wgt_9_473;input [WEIGHT_SIZE-1:0] Wgt_9_474;input [WEIGHT_SIZE-1:0] Wgt_9_475;input [WEIGHT_SIZE-1:0] Wgt_9_476;input [WEIGHT_SIZE-1:0] Wgt_9_477;input [WEIGHT_SIZE-1:0] Wgt_9_478;input [WEIGHT_SIZE-1:0] Wgt_9_479;input [WEIGHT_SIZE-1:0] Wgt_9_480;input [WEIGHT_SIZE-1:0] Wgt_9_481;input [WEIGHT_SIZE-1:0] Wgt_9_482;input [WEIGHT_SIZE-1:0] Wgt_9_483;input [WEIGHT_SIZE-1:0] Wgt_9_484;input [WEIGHT_SIZE-1:0] Wgt_9_485;input [WEIGHT_SIZE-1:0] Wgt_9_486;input [WEIGHT_SIZE-1:0] Wgt_9_487;input [WEIGHT_SIZE-1:0] Wgt_9_488;input [WEIGHT_SIZE-1:0] Wgt_9_489;input [WEIGHT_SIZE-1:0] Wgt_9_490;input [WEIGHT_SIZE-1:0] Wgt_9_491;input [WEIGHT_SIZE-1:0] Wgt_9_492;input [WEIGHT_SIZE-1:0] Wgt_9_493;input [WEIGHT_SIZE-1:0] Wgt_9_494;input [WEIGHT_SIZE-1:0] Wgt_9_495;input [WEIGHT_SIZE-1:0] Wgt_9_496;input [WEIGHT_SIZE-1:0] Wgt_9_497;input [WEIGHT_SIZE-1:0] Wgt_9_498;input [WEIGHT_SIZE-1:0] Wgt_9_499;input [WEIGHT_SIZE-1:0] Wgt_9_500;input [WEIGHT_SIZE-1:0] Wgt_9_501;input [WEIGHT_SIZE-1:0] Wgt_9_502;input [WEIGHT_SIZE-1:0] Wgt_9_503;input [WEIGHT_SIZE-1:0] Wgt_9_504;input [WEIGHT_SIZE-1:0] Wgt_9_505;input [WEIGHT_SIZE-1:0] Wgt_9_506;input [WEIGHT_SIZE-1:0] Wgt_9_507;input [WEIGHT_SIZE-1:0] Wgt_9_508;input [WEIGHT_SIZE-1:0] Wgt_9_509;input [WEIGHT_SIZE-1:0] Wgt_9_510;input [WEIGHT_SIZE-1:0] Wgt_9_511;input [WEIGHT_SIZE-1:0] Wgt_9_512;input [WEIGHT_SIZE-1:0] Wgt_9_513;input [WEIGHT_SIZE-1:0] Wgt_9_514;input [WEIGHT_SIZE-1:0] Wgt_9_515;input [WEIGHT_SIZE-1:0] Wgt_9_516;input [WEIGHT_SIZE-1:0] Wgt_9_517;input [WEIGHT_SIZE-1:0] Wgt_9_518;input [WEIGHT_SIZE-1:0] Wgt_9_519;input [WEIGHT_SIZE-1:0] Wgt_9_520;input [WEIGHT_SIZE-1:0] Wgt_9_521;input [WEIGHT_SIZE-1:0] Wgt_9_522;input [WEIGHT_SIZE-1:0] Wgt_9_523;input [WEIGHT_SIZE-1:0] Wgt_9_524;input [WEIGHT_SIZE-1:0] Wgt_9_525;input [WEIGHT_SIZE-1:0] Wgt_9_526;input [WEIGHT_SIZE-1:0] Wgt_9_527;input [WEIGHT_SIZE-1:0] Wgt_9_528;input [WEIGHT_SIZE-1:0] Wgt_9_529;input [WEIGHT_SIZE-1:0] Wgt_9_530;input [WEIGHT_SIZE-1:0] Wgt_9_531;input [WEIGHT_SIZE-1:0] Wgt_9_532;input [WEIGHT_SIZE-1:0] Wgt_9_533;input [WEIGHT_SIZE-1:0] Wgt_9_534;input [WEIGHT_SIZE-1:0] Wgt_9_535;input [WEIGHT_SIZE-1:0] Wgt_9_536;input [WEIGHT_SIZE-1:0] Wgt_9_537;input [WEIGHT_SIZE-1:0] Wgt_9_538;input [WEIGHT_SIZE-1:0] Wgt_9_539;input [WEIGHT_SIZE-1:0] Wgt_9_540;input [WEIGHT_SIZE-1:0] Wgt_9_541;input [WEIGHT_SIZE-1:0] Wgt_9_542;input [WEIGHT_SIZE-1:0] Wgt_9_543;input [WEIGHT_SIZE-1:0] Wgt_9_544;input [WEIGHT_SIZE-1:0] Wgt_9_545;input [WEIGHT_SIZE-1:0] Wgt_9_546;input [WEIGHT_SIZE-1:0] Wgt_9_547;input [WEIGHT_SIZE-1:0] Wgt_9_548;input [WEIGHT_SIZE-1:0] Wgt_9_549;input [WEIGHT_SIZE-1:0] Wgt_9_550;input [WEIGHT_SIZE-1:0] Wgt_9_551;input [WEIGHT_SIZE-1:0] Wgt_9_552;input [WEIGHT_SIZE-1:0] Wgt_9_553;input [WEIGHT_SIZE-1:0] Wgt_9_554;input [WEIGHT_SIZE-1:0] Wgt_9_555;input [WEIGHT_SIZE-1:0] Wgt_9_556;input [WEIGHT_SIZE-1:0] Wgt_9_557;input [WEIGHT_SIZE-1:0] Wgt_9_558;input [WEIGHT_SIZE-1:0] Wgt_9_559;input [WEIGHT_SIZE-1:0] Wgt_9_560;input [WEIGHT_SIZE-1:0] Wgt_9_561;input [WEIGHT_SIZE-1:0] Wgt_9_562;input [WEIGHT_SIZE-1:0] Wgt_9_563;input [WEIGHT_SIZE-1:0] Wgt_9_564;input [WEIGHT_SIZE-1:0] Wgt_9_565;input [WEIGHT_SIZE-1:0] Wgt_9_566;input [WEIGHT_SIZE-1:0] Wgt_9_567;input [WEIGHT_SIZE-1:0] Wgt_9_568;input [WEIGHT_SIZE-1:0] Wgt_9_569;input [WEIGHT_SIZE-1:0] Wgt_9_570;input [WEIGHT_SIZE-1:0] Wgt_9_571;input [WEIGHT_SIZE-1:0] Wgt_9_572;input [WEIGHT_SIZE-1:0] Wgt_9_573;input [WEIGHT_SIZE-1:0] Wgt_9_574;input [WEIGHT_SIZE-1:0] Wgt_9_575;input [WEIGHT_SIZE-1:0] Wgt_9_576;input [WEIGHT_SIZE-1:0] Wgt_9_577;input [WEIGHT_SIZE-1:0] Wgt_9_578;input [WEIGHT_SIZE-1:0] Wgt_9_579;input [WEIGHT_SIZE-1:0] Wgt_9_580;input [WEIGHT_SIZE-1:0] Wgt_9_581;input [WEIGHT_SIZE-1:0] Wgt_9_582;input [WEIGHT_SIZE-1:0] Wgt_9_583;input [WEIGHT_SIZE-1:0] Wgt_9_584;input [WEIGHT_SIZE-1:0] Wgt_9_585;input [WEIGHT_SIZE-1:0] Wgt_9_586;input [WEIGHT_SIZE-1:0] Wgt_9_587;input [WEIGHT_SIZE-1:0] Wgt_9_588;input [WEIGHT_SIZE-1:0] Wgt_9_589;input [WEIGHT_SIZE-1:0] Wgt_9_590;input [WEIGHT_SIZE-1:0] Wgt_9_591;input [WEIGHT_SIZE-1:0] Wgt_9_592;input [WEIGHT_SIZE-1:0] Wgt_9_593;input [WEIGHT_SIZE-1:0] Wgt_9_594;input [WEIGHT_SIZE-1:0] Wgt_9_595;input [WEIGHT_SIZE-1:0] Wgt_9_596;input [WEIGHT_SIZE-1:0] Wgt_9_597;input [WEIGHT_SIZE-1:0] Wgt_9_598;input [WEIGHT_SIZE-1:0] Wgt_9_599;input [WEIGHT_SIZE-1:0] Wgt_9_600;input [WEIGHT_SIZE-1:0] Wgt_9_601;input [WEIGHT_SIZE-1:0] Wgt_9_602;input [WEIGHT_SIZE-1:0] Wgt_9_603;input [WEIGHT_SIZE-1:0] Wgt_9_604;input [WEIGHT_SIZE-1:0] Wgt_9_605;input [WEIGHT_SIZE-1:0] Wgt_9_606;input [WEIGHT_SIZE-1:0] Wgt_9_607;input [WEIGHT_SIZE-1:0] Wgt_9_608;input [WEIGHT_SIZE-1:0] Wgt_9_609;input [WEIGHT_SIZE-1:0] Wgt_9_610;input [WEIGHT_SIZE-1:0] Wgt_9_611;input [WEIGHT_SIZE-1:0] Wgt_9_612;input [WEIGHT_SIZE-1:0] Wgt_9_613;input [WEIGHT_SIZE-1:0] Wgt_9_614;input [WEIGHT_SIZE-1:0] Wgt_9_615;input [WEIGHT_SIZE-1:0] Wgt_9_616;input [WEIGHT_SIZE-1:0] Wgt_9_617;input [WEIGHT_SIZE-1:0] Wgt_9_618;input [WEIGHT_SIZE-1:0] Wgt_9_619;input [WEIGHT_SIZE-1:0] Wgt_9_620;input [WEIGHT_SIZE-1:0] Wgt_9_621;input [WEIGHT_SIZE-1:0] Wgt_9_622;input [WEIGHT_SIZE-1:0] Wgt_9_623;input [WEIGHT_SIZE-1:0] Wgt_9_624;input [WEIGHT_SIZE-1:0] Wgt_9_625;input [WEIGHT_SIZE-1:0] Wgt_9_626;input [WEIGHT_SIZE-1:0] Wgt_9_627;input [WEIGHT_SIZE-1:0] Wgt_9_628;input [WEIGHT_SIZE-1:0] Wgt_9_629;input [WEIGHT_SIZE-1:0] Wgt_9_630;input [WEIGHT_SIZE-1:0] Wgt_9_631;input [WEIGHT_SIZE-1:0] Wgt_9_632;input [WEIGHT_SIZE-1:0] Wgt_9_633;input [WEIGHT_SIZE-1:0] Wgt_9_634;input [WEIGHT_SIZE-1:0] Wgt_9_635;input [WEIGHT_SIZE-1:0] Wgt_9_636;input [WEIGHT_SIZE-1:0] Wgt_9_637;input [WEIGHT_SIZE-1:0] Wgt_9_638;input [WEIGHT_SIZE-1:0] Wgt_9_639;input [WEIGHT_SIZE-1:0] Wgt_9_640;input [WEIGHT_SIZE-1:0] Wgt_9_641;input [WEIGHT_SIZE-1:0] Wgt_9_642;input [WEIGHT_SIZE-1:0] Wgt_9_643;input [WEIGHT_SIZE-1:0] Wgt_9_644;input [WEIGHT_SIZE-1:0] Wgt_9_645;input [WEIGHT_SIZE-1:0] Wgt_9_646;input [WEIGHT_SIZE-1:0] Wgt_9_647;input [WEIGHT_SIZE-1:0] Wgt_9_648;input [WEIGHT_SIZE-1:0] Wgt_9_649;input [WEIGHT_SIZE-1:0] Wgt_9_650;input [WEIGHT_SIZE-1:0] Wgt_9_651;input [WEIGHT_SIZE-1:0] Wgt_9_652;input [WEIGHT_SIZE-1:0] Wgt_9_653;input [WEIGHT_SIZE-1:0] Wgt_9_654;input [WEIGHT_SIZE-1:0] Wgt_9_655;input [WEIGHT_SIZE-1:0] Wgt_9_656;input [WEIGHT_SIZE-1:0] Wgt_9_657;input [WEIGHT_SIZE-1:0] Wgt_9_658;input [WEIGHT_SIZE-1:0] Wgt_9_659;input [WEIGHT_SIZE-1:0] Wgt_9_660;input [WEIGHT_SIZE-1:0] Wgt_9_661;input [WEIGHT_SIZE-1:0] Wgt_9_662;input [WEIGHT_SIZE-1:0] Wgt_9_663;input [WEIGHT_SIZE-1:0] Wgt_9_664;input [WEIGHT_SIZE-1:0] Wgt_9_665;input [WEIGHT_SIZE-1:0] Wgt_9_666;input [WEIGHT_SIZE-1:0] Wgt_9_667;input [WEIGHT_SIZE-1:0] Wgt_9_668;input [WEIGHT_SIZE-1:0] Wgt_9_669;input [WEIGHT_SIZE-1:0] Wgt_9_670;input [WEIGHT_SIZE-1:0] Wgt_9_671;input [WEIGHT_SIZE-1:0] Wgt_9_672;input [WEIGHT_SIZE-1:0] Wgt_9_673;input [WEIGHT_SIZE-1:0] Wgt_9_674;input [WEIGHT_SIZE-1:0] Wgt_9_675;input [WEIGHT_SIZE-1:0] Wgt_9_676;input [WEIGHT_SIZE-1:0] Wgt_9_677;input [WEIGHT_SIZE-1:0] Wgt_9_678;input [WEIGHT_SIZE-1:0] Wgt_9_679;input [WEIGHT_SIZE-1:0] Wgt_9_680;input [WEIGHT_SIZE-1:0] Wgt_9_681;input [WEIGHT_SIZE-1:0] Wgt_9_682;input [WEIGHT_SIZE-1:0] Wgt_9_683;input [WEIGHT_SIZE-1:0] Wgt_9_684;input [WEIGHT_SIZE-1:0] Wgt_9_685;input [WEIGHT_SIZE-1:0] Wgt_9_686;input [WEIGHT_SIZE-1:0] Wgt_9_687;input [WEIGHT_SIZE-1:0] Wgt_9_688;input [WEIGHT_SIZE-1:0] Wgt_9_689;input [WEIGHT_SIZE-1:0] Wgt_9_690;input [WEIGHT_SIZE-1:0] Wgt_9_691;input [WEIGHT_SIZE-1:0] Wgt_9_692;input [WEIGHT_SIZE-1:0] Wgt_9_693;input [WEIGHT_SIZE-1:0] Wgt_9_694;input [WEIGHT_SIZE-1:0] Wgt_9_695;input [WEIGHT_SIZE-1:0] Wgt_9_696;input [WEIGHT_SIZE-1:0] Wgt_9_697;input [WEIGHT_SIZE-1:0] Wgt_9_698;input [WEIGHT_SIZE-1:0] Wgt_9_699;input [WEIGHT_SIZE-1:0] Wgt_9_700;input [WEIGHT_SIZE-1:0] Wgt_9_701;input [WEIGHT_SIZE-1:0] Wgt_9_702;input [WEIGHT_SIZE-1:0] Wgt_9_703;input [WEIGHT_SIZE-1:0] Wgt_9_704;input [WEIGHT_SIZE-1:0] Wgt_9_705;input [WEIGHT_SIZE-1:0] Wgt_9_706;input [WEIGHT_SIZE-1:0] Wgt_9_707;input [WEIGHT_SIZE-1:0] Wgt_9_708;input [WEIGHT_SIZE-1:0] Wgt_9_709;input [WEIGHT_SIZE-1:0] Wgt_9_710;input [WEIGHT_SIZE-1:0] Wgt_9_711;input [WEIGHT_SIZE-1:0] Wgt_9_712;input [WEIGHT_SIZE-1:0] Wgt_9_713;input [WEIGHT_SIZE-1:0] Wgt_9_714;input [WEIGHT_SIZE-1:0] Wgt_9_715;input [WEIGHT_SIZE-1:0] Wgt_9_716;input [WEIGHT_SIZE-1:0] Wgt_9_717;input [WEIGHT_SIZE-1:0] Wgt_9_718;input [WEIGHT_SIZE-1:0] Wgt_9_719;input [WEIGHT_SIZE-1:0] Wgt_9_720;input [WEIGHT_SIZE-1:0] Wgt_9_721;input [WEIGHT_SIZE-1:0] Wgt_9_722;input [WEIGHT_SIZE-1:0] Wgt_9_723;input [WEIGHT_SIZE-1:0] Wgt_9_724;input [WEIGHT_SIZE-1:0] Wgt_9_725;input [WEIGHT_SIZE-1:0] Wgt_9_726;input [WEIGHT_SIZE-1:0] Wgt_9_727;input [WEIGHT_SIZE-1:0] Wgt_9_728;input [WEIGHT_SIZE-1:0] Wgt_9_729;input [WEIGHT_SIZE-1:0] Wgt_9_730;input [WEIGHT_SIZE-1:0] Wgt_9_731;input [WEIGHT_SIZE-1:0] Wgt_9_732;input [WEIGHT_SIZE-1:0] Wgt_9_733;input [WEIGHT_SIZE-1:0] Wgt_9_734;input [WEIGHT_SIZE-1:0] Wgt_9_735;input [WEIGHT_SIZE-1:0] Wgt_9_736;input [WEIGHT_SIZE-1:0] Wgt_9_737;input [WEIGHT_SIZE-1:0] Wgt_9_738;input [WEIGHT_SIZE-1:0] Wgt_9_739;input [WEIGHT_SIZE-1:0] Wgt_9_740;input [WEIGHT_SIZE-1:0] Wgt_9_741;input [WEIGHT_SIZE-1:0] Wgt_9_742;input [WEIGHT_SIZE-1:0] Wgt_9_743;input [WEIGHT_SIZE-1:0] Wgt_9_744;input [WEIGHT_SIZE-1:0] Wgt_9_745;input [WEIGHT_SIZE-1:0] Wgt_9_746;input [WEIGHT_SIZE-1:0] Wgt_9_747;input [WEIGHT_SIZE-1:0] Wgt_9_748;input [WEIGHT_SIZE-1:0] Wgt_9_749;input [WEIGHT_SIZE-1:0] Wgt_9_750;input [WEIGHT_SIZE-1:0] Wgt_9_751;input [WEIGHT_SIZE-1:0] Wgt_9_752;input [WEIGHT_SIZE-1:0] Wgt_9_753;input [WEIGHT_SIZE-1:0] Wgt_9_754;input [WEIGHT_SIZE-1:0] Wgt_9_755;input [WEIGHT_SIZE-1:0] Wgt_9_756;input [WEIGHT_SIZE-1:0] Wgt_9_757;input [WEIGHT_SIZE-1:0] Wgt_9_758;input [WEIGHT_SIZE-1:0] Wgt_9_759;input [WEIGHT_SIZE-1:0] Wgt_9_760;input [WEIGHT_SIZE-1:0] Wgt_9_761;input [WEIGHT_SIZE-1:0] Wgt_9_762;input [WEIGHT_SIZE-1:0] Wgt_9_763;input [WEIGHT_SIZE-1:0] Wgt_9_764;input [WEIGHT_SIZE-1:0] Wgt_9_765;input [WEIGHT_SIZE-1:0] Wgt_9_766;input [WEIGHT_SIZE-1:0] Wgt_9_767;input [WEIGHT_SIZE-1:0] Wgt_9_768;input [WEIGHT_SIZE-1:0] Wgt_9_769;input [WEIGHT_SIZE-1:0] Wgt_9_770;input [WEIGHT_SIZE-1:0] Wgt_9_771;input [WEIGHT_SIZE-1:0] Wgt_9_772;input [WEIGHT_SIZE-1:0] Wgt_9_773;input [WEIGHT_SIZE-1:0] Wgt_9_774;input [WEIGHT_SIZE-1:0] Wgt_9_775;input [WEIGHT_SIZE-1:0] Wgt_9_776;input [WEIGHT_SIZE-1:0] Wgt_9_777;input [WEIGHT_SIZE-1:0] Wgt_9_778;input [WEIGHT_SIZE-1:0] Wgt_9_779;input [WEIGHT_SIZE-1:0] Wgt_9_780;input [WEIGHT_SIZE-1:0] Wgt_9_781;input [WEIGHT_SIZE-1:0] Wgt_9_782;input [WEIGHT_SIZE-1:0] Wgt_9_783;input [WEIGHT_SIZE-1:0] Wgt_9_784;
input [PIXEL_SIZE-1:0] Pix_0;input [PIXEL_SIZE-1:0] Pix_1;input [PIXEL_SIZE-1:0] Pix_2;input [PIXEL_SIZE-1:0] Pix_3;input [PIXEL_SIZE-1:0] Pix_4;input [PIXEL_SIZE-1:0] Pix_5;input [PIXEL_SIZE-1:0] Pix_6;input [PIXEL_SIZE-1:0] Pix_7;input [PIXEL_SIZE-1:0] Pix_8;input [PIXEL_SIZE-1:0] Pix_9;input [PIXEL_SIZE-1:0] Pix_10;input [PIXEL_SIZE-1:0] Pix_11;input [PIXEL_SIZE-1:0] Pix_12;input [PIXEL_SIZE-1:0] Pix_13;input [PIXEL_SIZE-1:0] Pix_14;input [PIXEL_SIZE-1:0] Pix_15;input [PIXEL_SIZE-1:0] Pix_16;input [PIXEL_SIZE-1:0] Pix_17;input [PIXEL_SIZE-1:0] Pix_18;input [PIXEL_SIZE-1:0] Pix_19;input [PIXEL_SIZE-1:0] Pix_20;input [PIXEL_SIZE-1:0] Pix_21;input [PIXEL_SIZE-1:0] Pix_22;input [PIXEL_SIZE-1:0] Pix_23;input [PIXEL_SIZE-1:0] Pix_24;input [PIXEL_SIZE-1:0] Pix_25;input [PIXEL_SIZE-1:0] Pix_26;input [PIXEL_SIZE-1:0] Pix_27;input [PIXEL_SIZE-1:0] Pix_28;input [PIXEL_SIZE-1:0] Pix_29;input [PIXEL_SIZE-1:0] Pix_30;input [PIXEL_SIZE-1:0] Pix_31;input [PIXEL_SIZE-1:0] Pix_32;input [PIXEL_SIZE-1:0] Pix_33;input [PIXEL_SIZE-1:0] Pix_34;input [PIXEL_SIZE-1:0] Pix_35;input [PIXEL_SIZE-1:0] Pix_36;input [PIXEL_SIZE-1:0] Pix_37;input [PIXEL_SIZE-1:0] Pix_38;input [PIXEL_SIZE-1:0] Pix_39;input [PIXEL_SIZE-1:0] Pix_40;input [PIXEL_SIZE-1:0] Pix_41;input [PIXEL_SIZE-1:0] Pix_42;input [PIXEL_SIZE-1:0] Pix_43;input [PIXEL_SIZE-1:0] Pix_44;input [PIXEL_SIZE-1:0] Pix_45;input [PIXEL_SIZE-1:0] Pix_46;input [PIXEL_SIZE-1:0] Pix_47;input [PIXEL_SIZE-1:0] Pix_48;input [PIXEL_SIZE-1:0] Pix_49;input [PIXEL_SIZE-1:0] Pix_50;input [PIXEL_SIZE-1:0] Pix_51;input [PIXEL_SIZE-1:0] Pix_52;input [PIXEL_SIZE-1:0] Pix_53;input [PIXEL_SIZE-1:0] Pix_54;input [PIXEL_SIZE-1:0] Pix_55;input [PIXEL_SIZE-1:0] Pix_56;input [PIXEL_SIZE-1:0] Pix_57;input [PIXEL_SIZE-1:0] Pix_58;input [PIXEL_SIZE-1:0] Pix_59;input [PIXEL_SIZE-1:0] Pix_60;input [PIXEL_SIZE-1:0] Pix_61;input [PIXEL_SIZE-1:0] Pix_62;input [PIXEL_SIZE-1:0] Pix_63;input [PIXEL_SIZE-1:0] Pix_64;input [PIXEL_SIZE-1:0] Pix_65;input [PIXEL_SIZE-1:0] Pix_66;input [PIXEL_SIZE-1:0] Pix_67;input [PIXEL_SIZE-1:0] Pix_68;input [PIXEL_SIZE-1:0] Pix_69;input [PIXEL_SIZE-1:0] Pix_70;input [PIXEL_SIZE-1:0] Pix_71;input [PIXEL_SIZE-1:0] Pix_72;input [PIXEL_SIZE-1:0] Pix_73;input [PIXEL_SIZE-1:0] Pix_74;input [PIXEL_SIZE-1:0] Pix_75;input [PIXEL_SIZE-1:0] Pix_76;input [PIXEL_SIZE-1:0] Pix_77;input [PIXEL_SIZE-1:0] Pix_78;input [PIXEL_SIZE-1:0] Pix_79;input [PIXEL_SIZE-1:0] Pix_80;input [PIXEL_SIZE-1:0] Pix_81;input [PIXEL_SIZE-1:0] Pix_82;input [PIXEL_SIZE-1:0] Pix_83;input [PIXEL_SIZE-1:0] Pix_84;input [PIXEL_SIZE-1:0] Pix_85;input [PIXEL_SIZE-1:0] Pix_86;input [PIXEL_SIZE-1:0] Pix_87;input [PIXEL_SIZE-1:0] Pix_88;input [PIXEL_SIZE-1:0] Pix_89;input [PIXEL_SIZE-1:0] Pix_90;input [PIXEL_SIZE-1:0] Pix_91;input [PIXEL_SIZE-1:0] Pix_92;input [PIXEL_SIZE-1:0] Pix_93;input [PIXEL_SIZE-1:0] Pix_94;input [PIXEL_SIZE-1:0] Pix_95;input [PIXEL_SIZE-1:0] Pix_96;input [PIXEL_SIZE-1:0] Pix_97;input [PIXEL_SIZE-1:0] Pix_98;input [PIXEL_SIZE-1:0] Pix_99;input [PIXEL_SIZE-1:0] Pix_100;input [PIXEL_SIZE-1:0] Pix_101;input [PIXEL_SIZE-1:0] Pix_102;input [PIXEL_SIZE-1:0] Pix_103;input [PIXEL_SIZE-1:0] Pix_104;input [PIXEL_SIZE-1:0] Pix_105;input [PIXEL_SIZE-1:0] Pix_106;input [PIXEL_SIZE-1:0] Pix_107;input [PIXEL_SIZE-1:0] Pix_108;input [PIXEL_SIZE-1:0] Pix_109;input [PIXEL_SIZE-1:0] Pix_110;input [PIXEL_SIZE-1:0] Pix_111;input [PIXEL_SIZE-1:0] Pix_112;input [PIXEL_SIZE-1:0] Pix_113;input [PIXEL_SIZE-1:0] Pix_114;input [PIXEL_SIZE-1:0] Pix_115;input [PIXEL_SIZE-1:0] Pix_116;input [PIXEL_SIZE-1:0] Pix_117;input [PIXEL_SIZE-1:0] Pix_118;input [PIXEL_SIZE-1:0] Pix_119;input [PIXEL_SIZE-1:0] Pix_120;input [PIXEL_SIZE-1:0] Pix_121;input [PIXEL_SIZE-1:0] Pix_122;input [PIXEL_SIZE-1:0] Pix_123;input [PIXEL_SIZE-1:0] Pix_124;input [PIXEL_SIZE-1:0] Pix_125;input [PIXEL_SIZE-1:0] Pix_126;input [PIXEL_SIZE-1:0] Pix_127;input [PIXEL_SIZE-1:0] Pix_128;input [PIXEL_SIZE-1:0] Pix_129;input [PIXEL_SIZE-1:0] Pix_130;input [PIXEL_SIZE-1:0] Pix_131;input [PIXEL_SIZE-1:0] Pix_132;input [PIXEL_SIZE-1:0] Pix_133;input [PIXEL_SIZE-1:0] Pix_134;input [PIXEL_SIZE-1:0] Pix_135;input [PIXEL_SIZE-1:0] Pix_136;input [PIXEL_SIZE-1:0] Pix_137;input [PIXEL_SIZE-1:0] Pix_138;input [PIXEL_SIZE-1:0] Pix_139;input [PIXEL_SIZE-1:0] Pix_140;input [PIXEL_SIZE-1:0] Pix_141;input [PIXEL_SIZE-1:0] Pix_142;input [PIXEL_SIZE-1:0] Pix_143;input [PIXEL_SIZE-1:0] Pix_144;input [PIXEL_SIZE-1:0] Pix_145;input [PIXEL_SIZE-1:0] Pix_146;input [PIXEL_SIZE-1:0] Pix_147;input [PIXEL_SIZE-1:0] Pix_148;input [PIXEL_SIZE-1:0] Pix_149;input [PIXEL_SIZE-1:0] Pix_150;input [PIXEL_SIZE-1:0] Pix_151;input [PIXEL_SIZE-1:0] Pix_152;input [PIXEL_SIZE-1:0] Pix_153;input [PIXEL_SIZE-1:0] Pix_154;input [PIXEL_SIZE-1:0] Pix_155;input [PIXEL_SIZE-1:0] Pix_156;input [PIXEL_SIZE-1:0] Pix_157;input [PIXEL_SIZE-1:0] Pix_158;input [PIXEL_SIZE-1:0] Pix_159;input [PIXEL_SIZE-1:0] Pix_160;input [PIXEL_SIZE-1:0] Pix_161;input [PIXEL_SIZE-1:0] Pix_162;input [PIXEL_SIZE-1:0] Pix_163;input [PIXEL_SIZE-1:0] Pix_164;input [PIXEL_SIZE-1:0] Pix_165;input [PIXEL_SIZE-1:0] Pix_166;input [PIXEL_SIZE-1:0] Pix_167;input [PIXEL_SIZE-1:0] Pix_168;input [PIXEL_SIZE-1:0] Pix_169;input [PIXEL_SIZE-1:0] Pix_170;input [PIXEL_SIZE-1:0] Pix_171;input [PIXEL_SIZE-1:0] Pix_172;input [PIXEL_SIZE-1:0] Pix_173;input [PIXEL_SIZE-1:0] Pix_174;input [PIXEL_SIZE-1:0] Pix_175;input [PIXEL_SIZE-1:0] Pix_176;input [PIXEL_SIZE-1:0] Pix_177;input [PIXEL_SIZE-1:0] Pix_178;input [PIXEL_SIZE-1:0] Pix_179;input [PIXEL_SIZE-1:0] Pix_180;input [PIXEL_SIZE-1:0] Pix_181;input [PIXEL_SIZE-1:0] Pix_182;input [PIXEL_SIZE-1:0] Pix_183;input [PIXEL_SIZE-1:0] Pix_184;input [PIXEL_SIZE-1:0] Pix_185;input [PIXEL_SIZE-1:0] Pix_186;input [PIXEL_SIZE-1:0] Pix_187;input [PIXEL_SIZE-1:0] Pix_188;input [PIXEL_SIZE-1:0] Pix_189;input [PIXEL_SIZE-1:0] Pix_190;input [PIXEL_SIZE-1:0] Pix_191;input [PIXEL_SIZE-1:0] Pix_192;input [PIXEL_SIZE-1:0] Pix_193;input [PIXEL_SIZE-1:0] Pix_194;input [PIXEL_SIZE-1:0] Pix_195;input [PIXEL_SIZE-1:0] Pix_196;input [PIXEL_SIZE-1:0] Pix_197;input [PIXEL_SIZE-1:0] Pix_198;input [PIXEL_SIZE-1:0] Pix_199;input [PIXEL_SIZE-1:0] Pix_200;input [PIXEL_SIZE-1:0] Pix_201;input [PIXEL_SIZE-1:0] Pix_202;input [PIXEL_SIZE-1:0] Pix_203;input [PIXEL_SIZE-1:0] Pix_204;input [PIXEL_SIZE-1:0] Pix_205;input [PIXEL_SIZE-1:0] Pix_206;input [PIXEL_SIZE-1:0] Pix_207;input [PIXEL_SIZE-1:0] Pix_208;input [PIXEL_SIZE-1:0] Pix_209;input [PIXEL_SIZE-1:0] Pix_210;input [PIXEL_SIZE-1:0] Pix_211;input [PIXEL_SIZE-1:0] Pix_212;input [PIXEL_SIZE-1:0] Pix_213;input [PIXEL_SIZE-1:0] Pix_214;input [PIXEL_SIZE-1:0] Pix_215;input [PIXEL_SIZE-1:0] Pix_216;input [PIXEL_SIZE-1:0] Pix_217;input [PIXEL_SIZE-1:0] Pix_218;input [PIXEL_SIZE-1:0] Pix_219;input [PIXEL_SIZE-1:0] Pix_220;input [PIXEL_SIZE-1:0] Pix_221;input [PIXEL_SIZE-1:0] Pix_222;input [PIXEL_SIZE-1:0] Pix_223;input [PIXEL_SIZE-1:0] Pix_224;input [PIXEL_SIZE-1:0] Pix_225;input [PIXEL_SIZE-1:0] Pix_226;input [PIXEL_SIZE-1:0] Pix_227;input [PIXEL_SIZE-1:0] Pix_228;input [PIXEL_SIZE-1:0] Pix_229;input [PIXEL_SIZE-1:0] Pix_230;input [PIXEL_SIZE-1:0] Pix_231;input [PIXEL_SIZE-1:0] Pix_232;input [PIXEL_SIZE-1:0] Pix_233;input [PIXEL_SIZE-1:0] Pix_234;input [PIXEL_SIZE-1:0] Pix_235;input [PIXEL_SIZE-1:0] Pix_236;input [PIXEL_SIZE-1:0] Pix_237;input [PIXEL_SIZE-1:0] Pix_238;input [PIXEL_SIZE-1:0] Pix_239;input [PIXEL_SIZE-1:0] Pix_240;input [PIXEL_SIZE-1:0] Pix_241;input [PIXEL_SIZE-1:0] Pix_242;input [PIXEL_SIZE-1:0] Pix_243;input [PIXEL_SIZE-1:0] Pix_244;input [PIXEL_SIZE-1:0] Pix_245;input [PIXEL_SIZE-1:0] Pix_246;input [PIXEL_SIZE-1:0] Pix_247;input [PIXEL_SIZE-1:0] Pix_248;input [PIXEL_SIZE-1:0] Pix_249;input [PIXEL_SIZE-1:0] Pix_250;input [PIXEL_SIZE-1:0] Pix_251;input [PIXEL_SIZE-1:0] Pix_252;input [PIXEL_SIZE-1:0] Pix_253;input [PIXEL_SIZE-1:0] Pix_254;input [PIXEL_SIZE-1:0] Pix_255;input [PIXEL_SIZE-1:0] Pix_256;input [PIXEL_SIZE-1:0] Pix_257;input [PIXEL_SIZE-1:0] Pix_258;input [PIXEL_SIZE-1:0] Pix_259;input [PIXEL_SIZE-1:0] Pix_260;input [PIXEL_SIZE-1:0] Pix_261;input [PIXEL_SIZE-1:0] Pix_262;input [PIXEL_SIZE-1:0] Pix_263;input [PIXEL_SIZE-1:0] Pix_264;input [PIXEL_SIZE-1:0] Pix_265;input [PIXEL_SIZE-1:0] Pix_266;input [PIXEL_SIZE-1:0] Pix_267;input [PIXEL_SIZE-1:0] Pix_268;input [PIXEL_SIZE-1:0] Pix_269;input [PIXEL_SIZE-1:0] Pix_270;input [PIXEL_SIZE-1:0] Pix_271;input [PIXEL_SIZE-1:0] Pix_272;input [PIXEL_SIZE-1:0] Pix_273;input [PIXEL_SIZE-1:0] Pix_274;input [PIXEL_SIZE-1:0] Pix_275;input [PIXEL_SIZE-1:0] Pix_276;input [PIXEL_SIZE-1:0] Pix_277;input [PIXEL_SIZE-1:0] Pix_278;input [PIXEL_SIZE-1:0] Pix_279;input [PIXEL_SIZE-1:0] Pix_280;input [PIXEL_SIZE-1:0] Pix_281;input [PIXEL_SIZE-1:0] Pix_282;input [PIXEL_SIZE-1:0] Pix_283;input [PIXEL_SIZE-1:0] Pix_284;input [PIXEL_SIZE-1:0] Pix_285;input [PIXEL_SIZE-1:0] Pix_286;input [PIXEL_SIZE-1:0] Pix_287;input [PIXEL_SIZE-1:0] Pix_288;input [PIXEL_SIZE-1:0] Pix_289;input [PIXEL_SIZE-1:0] Pix_290;input [PIXEL_SIZE-1:0] Pix_291;input [PIXEL_SIZE-1:0] Pix_292;input [PIXEL_SIZE-1:0] Pix_293;input [PIXEL_SIZE-1:0] Pix_294;input [PIXEL_SIZE-1:0] Pix_295;input [PIXEL_SIZE-1:0] Pix_296;input [PIXEL_SIZE-1:0] Pix_297;input [PIXEL_SIZE-1:0] Pix_298;input [PIXEL_SIZE-1:0] Pix_299;input [PIXEL_SIZE-1:0] Pix_300;input [PIXEL_SIZE-1:0] Pix_301;input [PIXEL_SIZE-1:0] Pix_302;input [PIXEL_SIZE-1:0] Pix_303;input [PIXEL_SIZE-1:0] Pix_304;input [PIXEL_SIZE-1:0] Pix_305;input [PIXEL_SIZE-1:0] Pix_306;input [PIXEL_SIZE-1:0] Pix_307;input [PIXEL_SIZE-1:0] Pix_308;input [PIXEL_SIZE-1:0] Pix_309;input [PIXEL_SIZE-1:0] Pix_310;input [PIXEL_SIZE-1:0] Pix_311;input [PIXEL_SIZE-1:0] Pix_312;input [PIXEL_SIZE-1:0] Pix_313;input [PIXEL_SIZE-1:0] Pix_314;input [PIXEL_SIZE-1:0] Pix_315;input [PIXEL_SIZE-1:0] Pix_316;input [PIXEL_SIZE-1:0] Pix_317;input [PIXEL_SIZE-1:0] Pix_318;input [PIXEL_SIZE-1:0] Pix_319;input [PIXEL_SIZE-1:0] Pix_320;input [PIXEL_SIZE-1:0] Pix_321;input [PIXEL_SIZE-1:0] Pix_322;input [PIXEL_SIZE-1:0] Pix_323;input [PIXEL_SIZE-1:0] Pix_324;input [PIXEL_SIZE-1:0] Pix_325;input [PIXEL_SIZE-1:0] Pix_326;input [PIXEL_SIZE-1:0] Pix_327;input [PIXEL_SIZE-1:0] Pix_328;input [PIXEL_SIZE-1:0] Pix_329;input [PIXEL_SIZE-1:0] Pix_330;input [PIXEL_SIZE-1:0] Pix_331;input [PIXEL_SIZE-1:0] Pix_332;input [PIXEL_SIZE-1:0] Pix_333;input [PIXEL_SIZE-1:0] Pix_334;input [PIXEL_SIZE-1:0] Pix_335;input [PIXEL_SIZE-1:0] Pix_336;input [PIXEL_SIZE-1:0] Pix_337;input [PIXEL_SIZE-1:0] Pix_338;input [PIXEL_SIZE-1:0] Pix_339;input [PIXEL_SIZE-1:0] Pix_340;input [PIXEL_SIZE-1:0] Pix_341;input [PIXEL_SIZE-1:0] Pix_342;input [PIXEL_SIZE-1:0] Pix_343;input [PIXEL_SIZE-1:0] Pix_344;input [PIXEL_SIZE-1:0] Pix_345;input [PIXEL_SIZE-1:0] Pix_346;input [PIXEL_SIZE-1:0] Pix_347;input [PIXEL_SIZE-1:0] Pix_348;input [PIXEL_SIZE-1:0] Pix_349;input [PIXEL_SIZE-1:0] Pix_350;input [PIXEL_SIZE-1:0] Pix_351;input [PIXEL_SIZE-1:0] Pix_352;input [PIXEL_SIZE-1:0] Pix_353;input [PIXEL_SIZE-1:0] Pix_354;input [PIXEL_SIZE-1:0] Pix_355;input [PIXEL_SIZE-1:0] Pix_356;input [PIXEL_SIZE-1:0] Pix_357;input [PIXEL_SIZE-1:0] Pix_358;input [PIXEL_SIZE-1:0] Pix_359;input [PIXEL_SIZE-1:0] Pix_360;input [PIXEL_SIZE-1:0] Pix_361;input [PIXEL_SIZE-1:0] Pix_362;input [PIXEL_SIZE-1:0] Pix_363;input [PIXEL_SIZE-1:0] Pix_364;input [PIXEL_SIZE-1:0] Pix_365;input [PIXEL_SIZE-1:0] Pix_366;input [PIXEL_SIZE-1:0] Pix_367;input [PIXEL_SIZE-1:0] Pix_368;input [PIXEL_SIZE-1:0] Pix_369;input [PIXEL_SIZE-1:0] Pix_370;input [PIXEL_SIZE-1:0] Pix_371;input [PIXEL_SIZE-1:0] Pix_372;input [PIXEL_SIZE-1:0] Pix_373;input [PIXEL_SIZE-1:0] Pix_374;input [PIXEL_SIZE-1:0] Pix_375;input [PIXEL_SIZE-1:0] Pix_376;input [PIXEL_SIZE-1:0] Pix_377;input [PIXEL_SIZE-1:0] Pix_378;input [PIXEL_SIZE-1:0] Pix_379;input [PIXEL_SIZE-1:0] Pix_380;input [PIXEL_SIZE-1:0] Pix_381;input [PIXEL_SIZE-1:0] Pix_382;input [PIXEL_SIZE-1:0] Pix_383;input [PIXEL_SIZE-1:0] Pix_384;input [PIXEL_SIZE-1:0] Pix_385;input [PIXEL_SIZE-1:0] Pix_386;input [PIXEL_SIZE-1:0] Pix_387;input [PIXEL_SIZE-1:0] Pix_388;input [PIXEL_SIZE-1:0] Pix_389;input [PIXEL_SIZE-1:0] Pix_390;input [PIXEL_SIZE-1:0] Pix_391;input [PIXEL_SIZE-1:0] Pix_392;input [PIXEL_SIZE-1:0] Pix_393;input [PIXEL_SIZE-1:0] Pix_394;input [PIXEL_SIZE-1:0] Pix_395;input [PIXEL_SIZE-1:0] Pix_396;input [PIXEL_SIZE-1:0] Pix_397;input [PIXEL_SIZE-1:0] Pix_398;input [PIXEL_SIZE-1:0] Pix_399;input [PIXEL_SIZE-1:0] Pix_400;input [PIXEL_SIZE-1:0] Pix_401;input [PIXEL_SIZE-1:0] Pix_402;input [PIXEL_SIZE-1:0] Pix_403;input [PIXEL_SIZE-1:0] Pix_404;input [PIXEL_SIZE-1:0] Pix_405;input [PIXEL_SIZE-1:0] Pix_406;input [PIXEL_SIZE-1:0] Pix_407;input [PIXEL_SIZE-1:0] Pix_408;input [PIXEL_SIZE-1:0] Pix_409;input [PIXEL_SIZE-1:0] Pix_410;input [PIXEL_SIZE-1:0] Pix_411;input [PIXEL_SIZE-1:0] Pix_412;input [PIXEL_SIZE-1:0] Pix_413;input [PIXEL_SIZE-1:0] Pix_414;input [PIXEL_SIZE-1:0] Pix_415;input [PIXEL_SIZE-1:0] Pix_416;input [PIXEL_SIZE-1:0] Pix_417;input [PIXEL_SIZE-1:0] Pix_418;input [PIXEL_SIZE-1:0] Pix_419;input [PIXEL_SIZE-1:0] Pix_420;input [PIXEL_SIZE-1:0] Pix_421;input [PIXEL_SIZE-1:0] Pix_422;input [PIXEL_SIZE-1:0] Pix_423;input [PIXEL_SIZE-1:0] Pix_424;input [PIXEL_SIZE-1:0] Pix_425;input [PIXEL_SIZE-1:0] Pix_426;input [PIXEL_SIZE-1:0] Pix_427;input [PIXEL_SIZE-1:0] Pix_428;input [PIXEL_SIZE-1:0] Pix_429;input [PIXEL_SIZE-1:0] Pix_430;input [PIXEL_SIZE-1:0] Pix_431;input [PIXEL_SIZE-1:0] Pix_432;input [PIXEL_SIZE-1:0] Pix_433;input [PIXEL_SIZE-1:0] Pix_434;input [PIXEL_SIZE-1:0] Pix_435;input [PIXEL_SIZE-1:0] Pix_436;input [PIXEL_SIZE-1:0] Pix_437;input [PIXEL_SIZE-1:0] Pix_438;input [PIXEL_SIZE-1:0] Pix_439;input [PIXEL_SIZE-1:0] Pix_440;input [PIXEL_SIZE-1:0] Pix_441;input [PIXEL_SIZE-1:0] Pix_442;input [PIXEL_SIZE-1:0] Pix_443;input [PIXEL_SIZE-1:0] Pix_444;input [PIXEL_SIZE-1:0] Pix_445;input [PIXEL_SIZE-1:0] Pix_446;input [PIXEL_SIZE-1:0] Pix_447;input [PIXEL_SIZE-1:0] Pix_448;input [PIXEL_SIZE-1:0] Pix_449;input [PIXEL_SIZE-1:0] Pix_450;input [PIXEL_SIZE-1:0] Pix_451;input [PIXEL_SIZE-1:0] Pix_452;input [PIXEL_SIZE-1:0] Pix_453;input [PIXEL_SIZE-1:0] Pix_454;input [PIXEL_SIZE-1:0] Pix_455;input [PIXEL_SIZE-1:0] Pix_456;input [PIXEL_SIZE-1:0] Pix_457;input [PIXEL_SIZE-1:0] Pix_458;input [PIXEL_SIZE-1:0] Pix_459;input [PIXEL_SIZE-1:0] Pix_460;input [PIXEL_SIZE-1:0] Pix_461;input [PIXEL_SIZE-1:0] Pix_462;input [PIXEL_SIZE-1:0] Pix_463;input [PIXEL_SIZE-1:0] Pix_464;input [PIXEL_SIZE-1:0] Pix_465;input [PIXEL_SIZE-1:0] Pix_466;input [PIXEL_SIZE-1:0] Pix_467;input [PIXEL_SIZE-1:0] Pix_468;input [PIXEL_SIZE-1:0] Pix_469;input [PIXEL_SIZE-1:0] Pix_470;input [PIXEL_SIZE-1:0] Pix_471;input [PIXEL_SIZE-1:0] Pix_472;input [PIXEL_SIZE-1:0] Pix_473;input [PIXEL_SIZE-1:0] Pix_474;input [PIXEL_SIZE-1:0] Pix_475;input [PIXEL_SIZE-1:0] Pix_476;input [PIXEL_SIZE-1:0] Pix_477;input [PIXEL_SIZE-1:0] Pix_478;input [PIXEL_SIZE-1:0] Pix_479;input [PIXEL_SIZE-1:0] Pix_480;input [PIXEL_SIZE-1:0] Pix_481;input [PIXEL_SIZE-1:0] Pix_482;input [PIXEL_SIZE-1:0] Pix_483;input [PIXEL_SIZE-1:0] Pix_484;input [PIXEL_SIZE-1:0] Pix_485;input [PIXEL_SIZE-1:0] Pix_486;input [PIXEL_SIZE-1:0] Pix_487;input [PIXEL_SIZE-1:0] Pix_488;input [PIXEL_SIZE-1:0] Pix_489;input [PIXEL_SIZE-1:0] Pix_490;input [PIXEL_SIZE-1:0] Pix_491;input [PIXEL_SIZE-1:0] Pix_492;input [PIXEL_SIZE-1:0] Pix_493;input [PIXEL_SIZE-1:0] Pix_494;input [PIXEL_SIZE-1:0] Pix_495;input [PIXEL_SIZE-1:0] Pix_496;input [PIXEL_SIZE-1:0] Pix_497;input [PIXEL_SIZE-1:0] Pix_498;input [PIXEL_SIZE-1:0] Pix_499;input [PIXEL_SIZE-1:0] Pix_500;input [PIXEL_SIZE-1:0] Pix_501;input [PIXEL_SIZE-1:0] Pix_502;input [PIXEL_SIZE-1:0] Pix_503;input [PIXEL_SIZE-1:0] Pix_504;input [PIXEL_SIZE-1:0] Pix_505;input [PIXEL_SIZE-1:0] Pix_506;input [PIXEL_SIZE-1:0] Pix_507;input [PIXEL_SIZE-1:0] Pix_508;input [PIXEL_SIZE-1:0] Pix_509;input [PIXEL_SIZE-1:0] Pix_510;input [PIXEL_SIZE-1:0] Pix_511;input [PIXEL_SIZE-1:0] Pix_512;input [PIXEL_SIZE-1:0] Pix_513;input [PIXEL_SIZE-1:0] Pix_514;input [PIXEL_SIZE-1:0] Pix_515;input [PIXEL_SIZE-1:0] Pix_516;input [PIXEL_SIZE-1:0] Pix_517;input [PIXEL_SIZE-1:0] Pix_518;input [PIXEL_SIZE-1:0] Pix_519;input [PIXEL_SIZE-1:0] Pix_520;input [PIXEL_SIZE-1:0] Pix_521;input [PIXEL_SIZE-1:0] Pix_522;input [PIXEL_SIZE-1:0] Pix_523;input [PIXEL_SIZE-1:0] Pix_524;input [PIXEL_SIZE-1:0] Pix_525;input [PIXEL_SIZE-1:0] Pix_526;input [PIXEL_SIZE-1:0] Pix_527;input [PIXEL_SIZE-1:0] Pix_528;input [PIXEL_SIZE-1:0] Pix_529;input [PIXEL_SIZE-1:0] Pix_530;input [PIXEL_SIZE-1:0] Pix_531;input [PIXEL_SIZE-1:0] Pix_532;input [PIXEL_SIZE-1:0] Pix_533;input [PIXEL_SIZE-1:0] Pix_534;input [PIXEL_SIZE-1:0] Pix_535;input [PIXEL_SIZE-1:0] Pix_536;input [PIXEL_SIZE-1:0] Pix_537;input [PIXEL_SIZE-1:0] Pix_538;input [PIXEL_SIZE-1:0] Pix_539;input [PIXEL_SIZE-1:0] Pix_540;input [PIXEL_SIZE-1:0] Pix_541;input [PIXEL_SIZE-1:0] Pix_542;input [PIXEL_SIZE-1:0] Pix_543;input [PIXEL_SIZE-1:0] Pix_544;input [PIXEL_SIZE-1:0] Pix_545;input [PIXEL_SIZE-1:0] Pix_546;input [PIXEL_SIZE-1:0] Pix_547;input [PIXEL_SIZE-1:0] Pix_548;input [PIXEL_SIZE-1:0] Pix_549;input [PIXEL_SIZE-1:0] Pix_550;input [PIXEL_SIZE-1:0] Pix_551;input [PIXEL_SIZE-1:0] Pix_552;input [PIXEL_SIZE-1:0] Pix_553;input [PIXEL_SIZE-1:0] Pix_554;input [PIXEL_SIZE-1:0] Pix_555;input [PIXEL_SIZE-1:0] Pix_556;input [PIXEL_SIZE-1:0] Pix_557;input [PIXEL_SIZE-1:0] Pix_558;input [PIXEL_SIZE-1:0] Pix_559;input [PIXEL_SIZE-1:0] Pix_560;input [PIXEL_SIZE-1:0] Pix_561;input [PIXEL_SIZE-1:0] Pix_562;input [PIXEL_SIZE-1:0] Pix_563;input [PIXEL_SIZE-1:0] Pix_564;input [PIXEL_SIZE-1:0] Pix_565;input [PIXEL_SIZE-1:0] Pix_566;input [PIXEL_SIZE-1:0] Pix_567;input [PIXEL_SIZE-1:0] Pix_568;input [PIXEL_SIZE-1:0] Pix_569;input [PIXEL_SIZE-1:0] Pix_570;input [PIXEL_SIZE-1:0] Pix_571;input [PIXEL_SIZE-1:0] Pix_572;input [PIXEL_SIZE-1:0] Pix_573;input [PIXEL_SIZE-1:0] Pix_574;input [PIXEL_SIZE-1:0] Pix_575;input [PIXEL_SIZE-1:0] Pix_576;input [PIXEL_SIZE-1:0] Pix_577;input [PIXEL_SIZE-1:0] Pix_578;input [PIXEL_SIZE-1:0] Pix_579;input [PIXEL_SIZE-1:0] Pix_580;input [PIXEL_SIZE-1:0] Pix_581;input [PIXEL_SIZE-1:0] Pix_582;input [PIXEL_SIZE-1:0] Pix_583;input [PIXEL_SIZE-1:0] Pix_584;input [PIXEL_SIZE-1:0] Pix_585;input [PIXEL_SIZE-1:0] Pix_586;input [PIXEL_SIZE-1:0] Pix_587;input [PIXEL_SIZE-1:0] Pix_588;input [PIXEL_SIZE-1:0] Pix_589;input [PIXEL_SIZE-1:0] Pix_590;input [PIXEL_SIZE-1:0] Pix_591;input [PIXEL_SIZE-1:0] Pix_592;input [PIXEL_SIZE-1:0] Pix_593;input [PIXEL_SIZE-1:0] Pix_594;input [PIXEL_SIZE-1:0] Pix_595;input [PIXEL_SIZE-1:0] Pix_596;input [PIXEL_SIZE-1:0] Pix_597;input [PIXEL_SIZE-1:0] Pix_598;input [PIXEL_SIZE-1:0] Pix_599;input [PIXEL_SIZE-1:0] Pix_600;input [PIXEL_SIZE-1:0] Pix_601;input [PIXEL_SIZE-1:0] Pix_602;input [PIXEL_SIZE-1:0] Pix_603;input [PIXEL_SIZE-1:0] Pix_604;input [PIXEL_SIZE-1:0] Pix_605;input [PIXEL_SIZE-1:0] Pix_606;input [PIXEL_SIZE-1:0] Pix_607;input [PIXEL_SIZE-1:0] Pix_608;input [PIXEL_SIZE-1:0] Pix_609;input [PIXEL_SIZE-1:0] Pix_610;input [PIXEL_SIZE-1:0] Pix_611;input [PIXEL_SIZE-1:0] Pix_612;input [PIXEL_SIZE-1:0] Pix_613;input [PIXEL_SIZE-1:0] Pix_614;input [PIXEL_SIZE-1:0] Pix_615;input [PIXEL_SIZE-1:0] Pix_616;input [PIXEL_SIZE-1:0] Pix_617;input [PIXEL_SIZE-1:0] Pix_618;input [PIXEL_SIZE-1:0] Pix_619;input [PIXEL_SIZE-1:0] Pix_620;input [PIXEL_SIZE-1:0] Pix_621;input [PIXEL_SIZE-1:0] Pix_622;input [PIXEL_SIZE-1:0] Pix_623;input [PIXEL_SIZE-1:0] Pix_624;input [PIXEL_SIZE-1:0] Pix_625;input [PIXEL_SIZE-1:0] Pix_626;input [PIXEL_SIZE-1:0] Pix_627;input [PIXEL_SIZE-1:0] Pix_628;input [PIXEL_SIZE-1:0] Pix_629;input [PIXEL_SIZE-1:0] Pix_630;input [PIXEL_SIZE-1:0] Pix_631;input [PIXEL_SIZE-1:0] Pix_632;input [PIXEL_SIZE-1:0] Pix_633;input [PIXEL_SIZE-1:0] Pix_634;input [PIXEL_SIZE-1:0] Pix_635;input [PIXEL_SIZE-1:0] Pix_636;input [PIXEL_SIZE-1:0] Pix_637;input [PIXEL_SIZE-1:0] Pix_638;input [PIXEL_SIZE-1:0] Pix_639;input [PIXEL_SIZE-1:0] Pix_640;input [PIXEL_SIZE-1:0] Pix_641;input [PIXEL_SIZE-1:0] Pix_642;input [PIXEL_SIZE-1:0] Pix_643;input [PIXEL_SIZE-1:0] Pix_644;input [PIXEL_SIZE-1:0] Pix_645;input [PIXEL_SIZE-1:0] Pix_646;input [PIXEL_SIZE-1:0] Pix_647;input [PIXEL_SIZE-1:0] Pix_648;input [PIXEL_SIZE-1:0] Pix_649;input [PIXEL_SIZE-1:0] Pix_650;input [PIXEL_SIZE-1:0] Pix_651;input [PIXEL_SIZE-1:0] Pix_652;input [PIXEL_SIZE-1:0] Pix_653;input [PIXEL_SIZE-1:0] Pix_654;input [PIXEL_SIZE-1:0] Pix_655;input [PIXEL_SIZE-1:0] Pix_656;input [PIXEL_SIZE-1:0] Pix_657;input [PIXEL_SIZE-1:0] Pix_658;input [PIXEL_SIZE-1:0] Pix_659;input [PIXEL_SIZE-1:0] Pix_660;input [PIXEL_SIZE-1:0] Pix_661;input [PIXEL_SIZE-1:0] Pix_662;input [PIXEL_SIZE-1:0] Pix_663;input [PIXEL_SIZE-1:0] Pix_664;input [PIXEL_SIZE-1:0] Pix_665;input [PIXEL_SIZE-1:0] Pix_666;input [PIXEL_SIZE-1:0] Pix_667;input [PIXEL_SIZE-1:0] Pix_668;input [PIXEL_SIZE-1:0] Pix_669;input [PIXEL_SIZE-1:0] Pix_670;input [PIXEL_SIZE-1:0] Pix_671;input [PIXEL_SIZE-1:0] Pix_672;input [PIXEL_SIZE-1:0] Pix_673;input [PIXEL_SIZE-1:0] Pix_674;input [PIXEL_SIZE-1:0] Pix_675;input [PIXEL_SIZE-1:0] Pix_676;input [PIXEL_SIZE-1:0] Pix_677;input [PIXEL_SIZE-1:0] Pix_678;input [PIXEL_SIZE-1:0] Pix_679;input [PIXEL_SIZE-1:0] Pix_680;input [PIXEL_SIZE-1:0] Pix_681;input [PIXEL_SIZE-1:0] Pix_682;input [PIXEL_SIZE-1:0] Pix_683;input [PIXEL_SIZE-1:0] Pix_684;input [PIXEL_SIZE-1:0] Pix_685;input [PIXEL_SIZE-1:0] Pix_686;input [PIXEL_SIZE-1:0] Pix_687;input [PIXEL_SIZE-1:0] Pix_688;input [PIXEL_SIZE-1:0] Pix_689;input [PIXEL_SIZE-1:0] Pix_690;input [PIXEL_SIZE-1:0] Pix_691;input [PIXEL_SIZE-1:0] Pix_692;input [PIXEL_SIZE-1:0] Pix_693;input [PIXEL_SIZE-1:0] Pix_694;input [PIXEL_SIZE-1:0] Pix_695;input [PIXEL_SIZE-1:0] Pix_696;input [PIXEL_SIZE-1:0] Pix_697;input [PIXEL_SIZE-1:0] Pix_698;input [PIXEL_SIZE-1:0] Pix_699;input [PIXEL_SIZE-1:0] Pix_700;input [PIXEL_SIZE-1:0] Pix_701;input [PIXEL_SIZE-1:0] Pix_702;input [PIXEL_SIZE-1:0] Pix_703;input [PIXEL_SIZE-1:0] Pix_704;input [PIXEL_SIZE-1:0] Pix_705;input [PIXEL_SIZE-1:0] Pix_706;input [PIXEL_SIZE-1:0] Pix_707;input [PIXEL_SIZE-1:0] Pix_708;input [PIXEL_SIZE-1:0] Pix_709;input [PIXEL_SIZE-1:0] Pix_710;input [PIXEL_SIZE-1:0] Pix_711;input [PIXEL_SIZE-1:0] Pix_712;input [PIXEL_SIZE-1:0] Pix_713;input [PIXEL_SIZE-1:0] Pix_714;input [PIXEL_SIZE-1:0] Pix_715;input [PIXEL_SIZE-1:0] Pix_716;input [PIXEL_SIZE-1:0] Pix_717;input [PIXEL_SIZE-1:0] Pix_718;input [PIXEL_SIZE-1:0] Pix_719;input [PIXEL_SIZE-1:0] Pix_720;input [PIXEL_SIZE-1:0] Pix_721;input [PIXEL_SIZE-1:0] Pix_722;input [PIXEL_SIZE-1:0] Pix_723;input [PIXEL_SIZE-1:0] Pix_724;input [PIXEL_SIZE-1:0] Pix_725;input [PIXEL_SIZE-1:0] Pix_726;input [PIXEL_SIZE-1:0] Pix_727;input [PIXEL_SIZE-1:0] Pix_728;input [PIXEL_SIZE-1:0] Pix_729;input [PIXEL_SIZE-1:0] Pix_730;input [PIXEL_SIZE-1:0] Pix_731;input [PIXEL_SIZE-1:0] Pix_732;input [PIXEL_SIZE-1:0] Pix_733;input [PIXEL_SIZE-1:0] Pix_734;input [PIXEL_SIZE-1:0] Pix_735;input [PIXEL_SIZE-1:0] Pix_736;input [PIXEL_SIZE-1:0] Pix_737;input [PIXEL_SIZE-1:0] Pix_738;input [PIXEL_SIZE-1:0] Pix_739;input [PIXEL_SIZE-1:0] Pix_740;input [PIXEL_SIZE-1:0] Pix_741;input [PIXEL_SIZE-1:0] Pix_742;input [PIXEL_SIZE-1:0] Pix_743;input [PIXEL_SIZE-1:0] Pix_744;input [PIXEL_SIZE-1:0] Pix_745;input [PIXEL_SIZE-1:0] Pix_746;input [PIXEL_SIZE-1:0] Pix_747;input [PIXEL_SIZE-1:0] Pix_748;input [PIXEL_SIZE-1:0] Pix_749;input [PIXEL_SIZE-1:0] Pix_750;input [PIXEL_SIZE-1:0] Pix_751;input [PIXEL_SIZE-1:0] Pix_752;input [PIXEL_SIZE-1:0] Pix_753;input [PIXEL_SIZE-1:0] Pix_754;input [PIXEL_SIZE-1:0] Pix_755;input [PIXEL_SIZE-1:0] Pix_756;input [PIXEL_SIZE-1:0] Pix_757;input [PIXEL_SIZE-1:0] Pix_758;input [PIXEL_SIZE-1:0] Pix_759;input [PIXEL_SIZE-1:0] Pix_760;input [PIXEL_SIZE-1:0] Pix_761;input [PIXEL_SIZE-1:0] Pix_762;input [PIXEL_SIZE-1:0] Pix_763;input [PIXEL_SIZE-1:0] Pix_764;input [PIXEL_SIZE-1:0] Pix_765;input [PIXEL_SIZE-1:0] Pix_766;input [PIXEL_SIZE-1:0] Pix_767;input [PIXEL_SIZE-1:0] Pix_768;input [PIXEL_SIZE-1:0] Pix_769;input [PIXEL_SIZE-1:0] Pix_770;input [PIXEL_SIZE-1:0] Pix_771;input [PIXEL_SIZE-1:0] Pix_772;input [PIXEL_SIZE-1:0] Pix_773;input [PIXEL_SIZE-1:0] Pix_774;input [PIXEL_SIZE-1:0] Pix_775;input [PIXEL_SIZE-1:0] Pix_776;input [PIXEL_SIZE-1:0] Pix_777;input [PIXEL_SIZE-1:0] Pix_778;input [PIXEL_SIZE-1:0] Pix_779;input [PIXEL_SIZE-1:0] Pix_780;input [PIXEL_SIZE-1:0] Pix_781;input [PIXEL_SIZE-1:0] Pix_782;input [PIXEL_SIZE-1:0] Pix_783;input [PIXEL_SIZE-1:0] Pix_784;
output [3:0] Image_Number;
output Output_Valid;

reg[PIXEL_SIZE*PIXEL_N-1:0] PixelsStore;
reg[WEIGHT_SIZE*PIXEL_N-1:0] WeightsStore[0:NEURONS-1];
reg[31:0] switchCounter;
reg[`CLOG2(BUS_WIDTH)-1:0] busCounter;
reg[`CLOG2(PIXEL_N/BUS_WIDTH/PARALLEL)-1:0] shiftCounter;
reg ready;
reg internalReset;
wire[VAL_SIZE*NEURONS-1:0] value;
reg flag;

assign Output_Valid = ready;

genvar k;
genvar j;
generate
	for(k=0; k<NEURONS; k=k+1) begin:neurgen
        for(j=0; j<PARALLEL; j=j+1) begin:pargen
    		DotProductSt DP(.clk(clk),
    			.GlobalReset(internalReset),
    			.Pixels(PixelInput[j*PIXEL_N/PARALLEL*PIXEL_SIZE +: PIXEL_N/PARALLEL*PIXEL_SIZE]),
    			.Weights(WeightInput[k][j*PIXEL_N/PARALLEL*WEIGHT_SIZE +: PIXEL_N/PARALLEL*WEIGHT_SIZE]),
    			.value(value[VAL_SIZE*k +: VAL_SIZE]));
        end
	end
endgenerate

Max MX(.GlobalReset(internalReset),
	.Num(value),
	.Index(Image_Number));

always@(posedge clk) begin
	if(GlobalReset == 1'b0) begin
		switchCounter <= 0;
		busCounter <= 0;
		shiftCounter <= 0;
		ready <= 1'b0;
		internalReset <= 1'b1;
		WeightInput[0]<=0;WeightInput[1]<=0;WeightInput[2]<=0;WeightInput[3]<=0;WeightInput[4]<=0;WeightInput[5]<=0;WeightInput[6]<=0;WeightInput[7]<=0;WeightInput[8]<=0;WeightInput[9]<=0;
		PixelsStore<=0;
		WeightsStore[0]<=0;WeightsStore[1]<=0;WeightsStore[2]<=0;WeightsStore[3]<=0;WeightsStore[4]<=0;WeightsStore[5]<=0;WeightsStore[6]<=0;WeightsStore[7]<=0;WeightsStore[8]<=0;WeightsStore[9]<=0;
		flag <= 0;
	end
	else if(Input_Valid == 1'b1) begin
		switchCounter <= 0;
		busCounter <= 0;
		shiftCounter <= 0;
		ready <= 1'b0;
		internalReset <= 1'b1;
		PixelsStore[0*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_0;PixelsStore[1*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_1;PixelsStore[2*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_2;PixelsStore[3*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_3;PixelsStore[4*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_4;PixelsStore[5*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_5;PixelsStore[6*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_6;PixelsStore[7*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_7;PixelsStore[8*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_8;PixelsStore[9*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_9;PixelsStore[10*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_10;PixelsStore[11*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_11;PixelsStore[12*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_12;PixelsStore[13*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_13;PixelsStore[14*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_14;PixelsStore[15*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_15;PixelsStore[16*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_16;PixelsStore[17*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_17;PixelsStore[18*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_18;PixelsStore[19*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_19;PixelsStore[20*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_20;PixelsStore[21*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_21;PixelsStore[22*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_22;PixelsStore[23*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_23;PixelsStore[24*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_24;PixelsStore[25*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_25;PixelsStore[26*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_26;PixelsStore[27*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_27;PixelsStore[28*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_28;PixelsStore[29*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_29;PixelsStore[30*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_30;PixelsStore[31*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_31;PixelsStore[32*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_32;PixelsStore[33*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_33;PixelsStore[34*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_34;PixelsStore[35*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_35;PixelsStore[36*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_36;PixelsStore[37*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_37;PixelsStore[38*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_38;PixelsStore[39*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_39;PixelsStore[40*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_40;PixelsStore[41*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_41;PixelsStore[42*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_42;PixelsStore[43*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_43;PixelsStore[44*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_44;PixelsStore[45*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_45;PixelsStore[46*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_46;PixelsStore[47*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_47;PixelsStore[48*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_48;PixelsStore[49*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_49;PixelsStore[50*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_50;PixelsStore[51*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_51;PixelsStore[52*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_52;PixelsStore[53*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_53;PixelsStore[54*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_54;PixelsStore[55*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_55;PixelsStore[56*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_56;PixelsStore[57*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_57;PixelsStore[58*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_58;PixelsStore[59*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_59;PixelsStore[60*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_60;PixelsStore[61*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_61;PixelsStore[62*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_62;PixelsStore[63*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_63;PixelsStore[64*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_64;PixelsStore[65*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_65;PixelsStore[66*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_66;PixelsStore[67*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_67;PixelsStore[68*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_68;PixelsStore[69*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_69;PixelsStore[70*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_70;PixelsStore[71*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_71;PixelsStore[72*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_72;PixelsStore[73*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_73;PixelsStore[74*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_74;PixelsStore[75*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_75;PixelsStore[76*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_76;PixelsStore[77*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_77;PixelsStore[78*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_78;PixelsStore[79*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_79;PixelsStore[80*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_80;PixelsStore[81*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_81;PixelsStore[82*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_82;PixelsStore[83*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_83;PixelsStore[84*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_84;PixelsStore[85*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_85;PixelsStore[86*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_86;PixelsStore[87*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_87;PixelsStore[88*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_88;PixelsStore[89*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_89;PixelsStore[90*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_90;PixelsStore[91*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_91;PixelsStore[92*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_92;PixelsStore[93*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_93;PixelsStore[94*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_94;PixelsStore[95*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_95;PixelsStore[96*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_96;PixelsStore[97*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_97;PixelsStore[98*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_98;PixelsStore[99*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_99;PixelsStore[100*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_100;PixelsStore[101*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_101;PixelsStore[102*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_102;PixelsStore[103*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_103;PixelsStore[104*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_104;PixelsStore[105*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_105;PixelsStore[106*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_106;PixelsStore[107*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_107;PixelsStore[108*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_108;PixelsStore[109*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_109;PixelsStore[110*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_110;PixelsStore[111*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_111;PixelsStore[112*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_112;PixelsStore[113*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_113;PixelsStore[114*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_114;PixelsStore[115*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_115;PixelsStore[116*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_116;PixelsStore[117*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_117;PixelsStore[118*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_118;PixelsStore[119*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_119;PixelsStore[120*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_120;PixelsStore[121*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_121;PixelsStore[122*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_122;PixelsStore[123*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_123;PixelsStore[124*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_124;PixelsStore[125*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_125;PixelsStore[126*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_126;PixelsStore[127*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_127;PixelsStore[128*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_128;PixelsStore[129*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_129;PixelsStore[130*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_130;PixelsStore[131*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_131;PixelsStore[132*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_132;PixelsStore[133*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_133;PixelsStore[134*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_134;PixelsStore[135*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_135;PixelsStore[136*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_136;PixelsStore[137*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_137;PixelsStore[138*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_138;PixelsStore[139*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_139;PixelsStore[140*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_140;PixelsStore[141*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_141;PixelsStore[142*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_142;PixelsStore[143*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_143;PixelsStore[144*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_144;PixelsStore[145*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_145;PixelsStore[146*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_146;PixelsStore[147*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_147;PixelsStore[148*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_148;PixelsStore[149*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_149;PixelsStore[150*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_150;PixelsStore[151*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_151;PixelsStore[152*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_152;PixelsStore[153*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_153;PixelsStore[154*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_154;PixelsStore[155*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_155;PixelsStore[156*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_156;PixelsStore[157*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_157;PixelsStore[158*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_158;PixelsStore[159*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_159;PixelsStore[160*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_160;PixelsStore[161*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_161;PixelsStore[162*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_162;PixelsStore[163*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_163;PixelsStore[164*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_164;PixelsStore[165*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_165;PixelsStore[166*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_166;PixelsStore[167*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_167;PixelsStore[168*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_168;PixelsStore[169*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_169;PixelsStore[170*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_170;PixelsStore[171*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_171;PixelsStore[172*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_172;PixelsStore[173*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_173;PixelsStore[174*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_174;PixelsStore[175*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_175;PixelsStore[176*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_176;PixelsStore[177*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_177;PixelsStore[178*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_178;PixelsStore[179*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_179;PixelsStore[180*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_180;PixelsStore[181*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_181;PixelsStore[182*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_182;PixelsStore[183*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_183;PixelsStore[184*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_184;PixelsStore[185*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_185;PixelsStore[186*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_186;PixelsStore[187*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_187;PixelsStore[188*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_188;PixelsStore[189*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_189;PixelsStore[190*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_190;PixelsStore[191*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_191;PixelsStore[192*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_192;PixelsStore[193*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_193;PixelsStore[194*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_194;PixelsStore[195*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_195;PixelsStore[196*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_196;PixelsStore[197*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_197;PixelsStore[198*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_198;PixelsStore[199*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_199;PixelsStore[200*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_200;PixelsStore[201*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_201;PixelsStore[202*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_202;PixelsStore[203*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_203;PixelsStore[204*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_204;PixelsStore[205*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_205;PixelsStore[206*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_206;PixelsStore[207*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_207;PixelsStore[208*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_208;PixelsStore[209*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_209;PixelsStore[210*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_210;PixelsStore[211*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_211;PixelsStore[212*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_212;PixelsStore[213*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_213;PixelsStore[214*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_214;PixelsStore[215*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_215;PixelsStore[216*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_216;PixelsStore[217*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_217;PixelsStore[218*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_218;PixelsStore[219*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_219;PixelsStore[220*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_220;PixelsStore[221*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_221;PixelsStore[222*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_222;PixelsStore[223*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_223;PixelsStore[224*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_224;PixelsStore[225*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_225;PixelsStore[226*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_226;PixelsStore[227*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_227;PixelsStore[228*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_228;PixelsStore[229*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_229;PixelsStore[230*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_230;PixelsStore[231*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_231;PixelsStore[232*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_232;PixelsStore[233*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_233;PixelsStore[234*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_234;PixelsStore[235*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_235;PixelsStore[236*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_236;PixelsStore[237*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_237;PixelsStore[238*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_238;PixelsStore[239*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_239;PixelsStore[240*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_240;PixelsStore[241*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_241;PixelsStore[242*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_242;PixelsStore[243*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_243;PixelsStore[244*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_244;PixelsStore[245*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_245;PixelsStore[246*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_246;PixelsStore[247*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_247;PixelsStore[248*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_248;PixelsStore[249*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_249;PixelsStore[250*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_250;PixelsStore[251*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_251;PixelsStore[252*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_252;PixelsStore[253*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_253;PixelsStore[254*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_254;PixelsStore[255*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_255;PixelsStore[256*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_256;PixelsStore[257*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_257;PixelsStore[258*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_258;PixelsStore[259*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_259;PixelsStore[260*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_260;PixelsStore[261*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_261;PixelsStore[262*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_262;PixelsStore[263*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_263;PixelsStore[264*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_264;PixelsStore[265*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_265;PixelsStore[266*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_266;PixelsStore[267*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_267;PixelsStore[268*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_268;PixelsStore[269*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_269;PixelsStore[270*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_270;PixelsStore[271*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_271;PixelsStore[272*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_272;PixelsStore[273*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_273;PixelsStore[274*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_274;PixelsStore[275*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_275;PixelsStore[276*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_276;PixelsStore[277*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_277;PixelsStore[278*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_278;PixelsStore[279*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_279;PixelsStore[280*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_280;PixelsStore[281*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_281;PixelsStore[282*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_282;PixelsStore[283*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_283;PixelsStore[284*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_284;PixelsStore[285*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_285;PixelsStore[286*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_286;PixelsStore[287*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_287;PixelsStore[288*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_288;PixelsStore[289*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_289;PixelsStore[290*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_290;PixelsStore[291*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_291;PixelsStore[292*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_292;PixelsStore[293*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_293;PixelsStore[294*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_294;PixelsStore[295*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_295;PixelsStore[296*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_296;PixelsStore[297*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_297;PixelsStore[298*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_298;PixelsStore[299*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_299;PixelsStore[300*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_300;PixelsStore[301*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_301;PixelsStore[302*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_302;PixelsStore[303*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_303;PixelsStore[304*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_304;PixelsStore[305*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_305;PixelsStore[306*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_306;PixelsStore[307*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_307;PixelsStore[308*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_308;PixelsStore[309*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_309;PixelsStore[310*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_310;PixelsStore[311*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_311;PixelsStore[312*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_312;PixelsStore[313*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_313;PixelsStore[314*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_314;PixelsStore[315*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_315;PixelsStore[316*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_316;PixelsStore[317*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_317;PixelsStore[318*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_318;PixelsStore[319*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_319;PixelsStore[320*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_320;PixelsStore[321*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_321;PixelsStore[322*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_322;PixelsStore[323*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_323;PixelsStore[324*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_324;PixelsStore[325*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_325;PixelsStore[326*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_326;PixelsStore[327*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_327;PixelsStore[328*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_328;PixelsStore[329*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_329;PixelsStore[330*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_330;PixelsStore[331*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_331;PixelsStore[332*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_332;PixelsStore[333*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_333;PixelsStore[334*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_334;PixelsStore[335*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_335;PixelsStore[336*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_336;PixelsStore[337*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_337;PixelsStore[338*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_338;PixelsStore[339*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_339;PixelsStore[340*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_340;PixelsStore[341*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_341;PixelsStore[342*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_342;PixelsStore[343*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_343;PixelsStore[344*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_344;PixelsStore[345*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_345;PixelsStore[346*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_346;PixelsStore[347*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_347;PixelsStore[348*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_348;PixelsStore[349*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_349;PixelsStore[350*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_350;PixelsStore[351*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_351;PixelsStore[352*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_352;PixelsStore[353*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_353;PixelsStore[354*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_354;PixelsStore[355*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_355;PixelsStore[356*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_356;PixelsStore[357*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_357;PixelsStore[358*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_358;PixelsStore[359*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_359;PixelsStore[360*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_360;PixelsStore[361*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_361;PixelsStore[362*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_362;PixelsStore[363*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_363;PixelsStore[364*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_364;PixelsStore[365*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_365;PixelsStore[366*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_366;PixelsStore[367*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_367;PixelsStore[368*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_368;PixelsStore[369*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_369;PixelsStore[370*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_370;PixelsStore[371*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_371;PixelsStore[372*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_372;PixelsStore[373*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_373;PixelsStore[374*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_374;PixelsStore[375*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_375;PixelsStore[376*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_376;PixelsStore[377*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_377;PixelsStore[378*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_378;PixelsStore[379*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_379;PixelsStore[380*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_380;PixelsStore[381*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_381;PixelsStore[382*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_382;PixelsStore[383*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_383;PixelsStore[384*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_384;PixelsStore[385*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_385;PixelsStore[386*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_386;PixelsStore[387*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_387;PixelsStore[388*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_388;PixelsStore[389*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_389;PixelsStore[390*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_390;PixelsStore[391*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_391;PixelsStore[392*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_392;PixelsStore[393*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_393;PixelsStore[394*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_394;PixelsStore[395*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_395;PixelsStore[396*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_396;PixelsStore[397*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_397;PixelsStore[398*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_398;PixelsStore[399*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_399;PixelsStore[400*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_400;PixelsStore[401*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_401;PixelsStore[402*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_402;PixelsStore[403*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_403;PixelsStore[404*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_404;PixelsStore[405*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_405;PixelsStore[406*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_406;PixelsStore[407*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_407;PixelsStore[408*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_408;PixelsStore[409*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_409;PixelsStore[410*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_410;PixelsStore[411*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_411;PixelsStore[412*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_412;PixelsStore[413*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_413;PixelsStore[414*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_414;PixelsStore[415*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_415;PixelsStore[416*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_416;PixelsStore[417*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_417;PixelsStore[418*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_418;PixelsStore[419*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_419;PixelsStore[420*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_420;PixelsStore[421*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_421;PixelsStore[422*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_422;PixelsStore[423*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_423;PixelsStore[424*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_424;PixelsStore[425*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_425;PixelsStore[426*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_426;PixelsStore[427*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_427;PixelsStore[428*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_428;PixelsStore[429*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_429;PixelsStore[430*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_430;PixelsStore[431*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_431;PixelsStore[432*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_432;PixelsStore[433*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_433;PixelsStore[434*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_434;PixelsStore[435*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_435;PixelsStore[436*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_436;PixelsStore[437*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_437;PixelsStore[438*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_438;PixelsStore[439*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_439;PixelsStore[440*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_440;PixelsStore[441*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_441;PixelsStore[442*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_442;PixelsStore[443*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_443;PixelsStore[444*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_444;PixelsStore[445*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_445;PixelsStore[446*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_446;PixelsStore[447*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_447;PixelsStore[448*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_448;PixelsStore[449*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_449;PixelsStore[450*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_450;PixelsStore[451*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_451;PixelsStore[452*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_452;PixelsStore[453*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_453;PixelsStore[454*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_454;PixelsStore[455*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_455;PixelsStore[456*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_456;PixelsStore[457*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_457;PixelsStore[458*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_458;PixelsStore[459*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_459;PixelsStore[460*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_460;PixelsStore[461*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_461;PixelsStore[462*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_462;PixelsStore[463*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_463;PixelsStore[464*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_464;PixelsStore[465*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_465;PixelsStore[466*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_466;PixelsStore[467*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_467;PixelsStore[468*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_468;PixelsStore[469*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_469;PixelsStore[470*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_470;PixelsStore[471*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_471;PixelsStore[472*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_472;PixelsStore[473*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_473;PixelsStore[474*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_474;PixelsStore[475*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_475;PixelsStore[476*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_476;PixelsStore[477*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_477;PixelsStore[478*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_478;PixelsStore[479*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_479;PixelsStore[480*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_480;PixelsStore[481*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_481;PixelsStore[482*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_482;PixelsStore[483*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_483;PixelsStore[484*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_484;PixelsStore[485*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_485;PixelsStore[486*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_486;PixelsStore[487*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_487;PixelsStore[488*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_488;PixelsStore[489*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_489;PixelsStore[490*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_490;PixelsStore[491*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_491;PixelsStore[492*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_492;PixelsStore[493*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_493;PixelsStore[494*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_494;PixelsStore[495*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_495;PixelsStore[496*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_496;PixelsStore[497*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_497;PixelsStore[498*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_498;PixelsStore[499*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_499;PixelsStore[500*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_500;PixelsStore[501*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_501;PixelsStore[502*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_502;PixelsStore[503*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_503;PixelsStore[504*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_504;PixelsStore[505*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_505;PixelsStore[506*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_506;PixelsStore[507*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_507;PixelsStore[508*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_508;PixelsStore[509*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_509;PixelsStore[510*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_510;PixelsStore[511*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_511;PixelsStore[512*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_512;PixelsStore[513*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_513;PixelsStore[514*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_514;PixelsStore[515*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_515;PixelsStore[516*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_516;PixelsStore[517*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_517;PixelsStore[518*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_518;PixelsStore[519*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_519;PixelsStore[520*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_520;PixelsStore[521*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_521;PixelsStore[522*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_522;PixelsStore[523*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_523;PixelsStore[524*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_524;PixelsStore[525*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_525;PixelsStore[526*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_526;PixelsStore[527*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_527;PixelsStore[528*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_528;PixelsStore[529*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_529;PixelsStore[530*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_530;PixelsStore[531*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_531;PixelsStore[532*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_532;PixelsStore[533*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_533;PixelsStore[534*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_534;PixelsStore[535*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_535;PixelsStore[536*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_536;PixelsStore[537*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_537;PixelsStore[538*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_538;PixelsStore[539*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_539;PixelsStore[540*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_540;PixelsStore[541*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_541;PixelsStore[542*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_542;PixelsStore[543*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_543;PixelsStore[544*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_544;PixelsStore[545*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_545;PixelsStore[546*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_546;PixelsStore[547*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_547;PixelsStore[548*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_548;PixelsStore[549*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_549;PixelsStore[550*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_550;PixelsStore[551*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_551;PixelsStore[552*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_552;PixelsStore[553*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_553;PixelsStore[554*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_554;PixelsStore[555*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_555;PixelsStore[556*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_556;PixelsStore[557*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_557;PixelsStore[558*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_558;PixelsStore[559*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_559;PixelsStore[560*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_560;PixelsStore[561*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_561;PixelsStore[562*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_562;PixelsStore[563*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_563;PixelsStore[564*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_564;PixelsStore[565*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_565;PixelsStore[566*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_566;PixelsStore[567*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_567;PixelsStore[568*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_568;PixelsStore[569*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_569;PixelsStore[570*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_570;PixelsStore[571*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_571;PixelsStore[572*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_572;PixelsStore[573*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_573;PixelsStore[574*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_574;PixelsStore[575*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_575;PixelsStore[576*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_576;PixelsStore[577*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_577;PixelsStore[578*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_578;PixelsStore[579*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_579;PixelsStore[580*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_580;PixelsStore[581*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_581;PixelsStore[582*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_582;PixelsStore[583*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_583;PixelsStore[584*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_584;PixelsStore[585*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_585;PixelsStore[586*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_586;PixelsStore[587*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_587;PixelsStore[588*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_588;PixelsStore[589*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_589;PixelsStore[590*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_590;PixelsStore[591*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_591;PixelsStore[592*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_592;PixelsStore[593*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_593;PixelsStore[594*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_594;PixelsStore[595*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_595;PixelsStore[596*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_596;PixelsStore[597*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_597;PixelsStore[598*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_598;PixelsStore[599*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_599;PixelsStore[600*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_600;PixelsStore[601*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_601;PixelsStore[602*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_602;PixelsStore[603*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_603;PixelsStore[604*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_604;PixelsStore[605*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_605;PixelsStore[606*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_606;PixelsStore[607*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_607;PixelsStore[608*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_608;PixelsStore[609*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_609;PixelsStore[610*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_610;PixelsStore[611*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_611;PixelsStore[612*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_612;PixelsStore[613*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_613;PixelsStore[614*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_614;PixelsStore[615*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_615;PixelsStore[616*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_616;PixelsStore[617*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_617;PixelsStore[618*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_618;PixelsStore[619*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_619;PixelsStore[620*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_620;PixelsStore[621*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_621;PixelsStore[622*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_622;PixelsStore[623*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_623;PixelsStore[624*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_624;PixelsStore[625*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_625;PixelsStore[626*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_626;PixelsStore[627*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_627;PixelsStore[628*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_628;PixelsStore[629*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_629;PixelsStore[630*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_630;PixelsStore[631*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_631;PixelsStore[632*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_632;PixelsStore[633*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_633;PixelsStore[634*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_634;PixelsStore[635*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_635;PixelsStore[636*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_636;PixelsStore[637*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_637;PixelsStore[638*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_638;PixelsStore[639*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_639;PixelsStore[640*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_640;PixelsStore[641*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_641;PixelsStore[642*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_642;PixelsStore[643*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_643;PixelsStore[644*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_644;PixelsStore[645*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_645;PixelsStore[646*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_646;PixelsStore[647*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_647;PixelsStore[648*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_648;PixelsStore[649*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_649;PixelsStore[650*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_650;PixelsStore[651*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_651;PixelsStore[652*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_652;PixelsStore[653*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_653;PixelsStore[654*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_654;PixelsStore[655*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_655;PixelsStore[656*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_656;PixelsStore[657*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_657;PixelsStore[658*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_658;PixelsStore[659*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_659;PixelsStore[660*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_660;PixelsStore[661*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_661;PixelsStore[662*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_662;PixelsStore[663*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_663;PixelsStore[664*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_664;PixelsStore[665*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_665;PixelsStore[666*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_666;PixelsStore[667*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_667;PixelsStore[668*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_668;PixelsStore[669*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_669;PixelsStore[670*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_670;PixelsStore[671*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_671;PixelsStore[672*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_672;PixelsStore[673*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_673;PixelsStore[674*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_674;PixelsStore[675*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_675;PixelsStore[676*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_676;PixelsStore[677*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_677;PixelsStore[678*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_678;PixelsStore[679*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_679;PixelsStore[680*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_680;PixelsStore[681*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_681;PixelsStore[682*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_682;PixelsStore[683*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_683;PixelsStore[684*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_684;PixelsStore[685*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_685;PixelsStore[686*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_686;PixelsStore[687*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_687;PixelsStore[688*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_688;PixelsStore[689*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_689;PixelsStore[690*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_690;PixelsStore[691*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_691;PixelsStore[692*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_692;PixelsStore[693*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_693;PixelsStore[694*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_694;PixelsStore[695*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_695;PixelsStore[696*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_696;PixelsStore[697*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_697;PixelsStore[698*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_698;PixelsStore[699*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_699;PixelsStore[700*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_700;PixelsStore[701*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_701;PixelsStore[702*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_702;PixelsStore[703*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_703;PixelsStore[704*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_704;PixelsStore[705*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_705;PixelsStore[706*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_706;PixelsStore[707*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_707;PixelsStore[708*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_708;PixelsStore[709*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_709;PixelsStore[710*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_710;PixelsStore[711*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_711;PixelsStore[712*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_712;PixelsStore[713*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_713;PixelsStore[714*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_714;PixelsStore[715*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_715;PixelsStore[716*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_716;PixelsStore[717*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_717;PixelsStore[718*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_718;PixelsStore[719*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_719;PixelsStore[720*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_720;PixelsStore[721*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_721;PixelsStore[722*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_722;PixelsStore[723*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_723;PixelsStore[724*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_724;PixelsStore[725*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_725;PixelsStore[726*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_726;PixelsStore[727*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_727;PixelsStore[728*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_728;PixelsStore[729*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_729;PixelsStore[730*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_730;PixelsStore[731*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_731;PixelsStore[732*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_732;PixelsStore[733*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_733;PixelsStore[734*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_734;PixelsStore[735*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_735;PixelsStore[736*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_736;PixelsStore[737*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_737;PixelsStore[738*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_738;PixelsStore[739*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_739;PixelsStore[740*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_740;PixelsStore[741*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_741;PixelsStore[742*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_742;PixelsStore[743*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_743;PixelsStore[744*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_744;PixelsStore[745*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_745;PixelsStore[746*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_746;PixelsStore[747*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_747;PixelsStore[748*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_748;PixelsStore[749*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_749;PixelsStore[750*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_750;PixelsStore[751*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_751;PixelsStore[752*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_752;PixelsStore[753*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_753;PixelsStore[754*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_754;PixelsStore[755*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_755;PixelsStore[756*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_756;PixelsStore[757*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_757;PixelsStore[758*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_758;PixelsStore[759*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_759;PixelsStore[760*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_760;PixelsStore[761*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_761;PixelsStore[762*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_762;PixelsStore[763*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_763;PixelsStore[764*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_764;PixelsStore[765*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_765;PixelsStore[766*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_766;PixelsStore[767*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_767;PixelsStore[768*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_768;PixelsStore[769*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_769;PixelsStore[770*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_770;PixelsStore[771*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_771;PixelsStore[772*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_772;PixelsStore[773*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_773;PixelsStore[774*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_774;PixelsStore[775*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_775;PixelsStore[776*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_776;PixelsStore[777*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_777;PixelsStore[778*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_778;PixelsStore[779*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_779;PixelsStore[780*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_780;PixelsStore[781*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_781;PixelsStore[782*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_782;PixelsStore[783*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_783;PixelsStore[784*PIXEL_SIZE+:PIXEL_SIZE]<=Pix_784;
		WeightsStore[0][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_0;WeightsStore[0][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_1;WeightsStore[0][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_2;WeightsStore[0][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_3;WeightsStore[0][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_4;WeightsStore[0][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_5;WeightsStore[0][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_6;WeightsStore[0][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_7;WeightsStore[0][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_8;WeightsStore[0][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_9;WeightsStore[0][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_10;WeightsStore[0][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_11;WeightsStore[0][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_12;WeightsStore[0][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_13;WeightsStore[0][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_14;WeightsStore[0][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_15;WeightsStore[0][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_16;WeightsStore[0][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_17;WeightsStore[0][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_18;WeightsStore[0][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_19;WeightsStore[0][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_20;WeightsStore[0][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_21;WeightsStore[0][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_22;WeightsStore[0][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_23;WeightsStore[0][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_24;WeightsStore[0][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_25;WeightsStore[0][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_26;WeightsStore[0][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_27;WeightsStore[0][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_28;WeightsStore[0][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_29;WeightsStore[0][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_30;WeightsStore[0][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_31;WeightsStore[0][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_32;WeightsStore[0][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_33;WeightsStore[0][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_34;WeightsStore[0][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_35;WeightsStore[0][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_36;WeightsStore[0][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_37;WeightsStore[0][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_38;WeightsStore[0][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_39;WeightsStore[0][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_40;WeightsStore[0][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_41;WeightsStore[0][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_42;WeightsStore[0][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_43;WeightsStore[0][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_44;WeightsStore[0][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_45;WeightsStore[0][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_46;WeightsStore[0][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_47;WeightsStore[0][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_48;WeightsStore[0][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_49;WeightsStore[0][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_50;WeightsStore[0][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_51;WeightsStore[0][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_52;WeightsStore[0][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_53;WeightsStore[0][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_54;WeightsStore[0][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_55;WeightsStore[0][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_56;WeightsStore[0][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_57;WeightsStore[0][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_58;WeightsStore[0][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_59;WeightsStore[0][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_60;WeightsStore[0][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_61;WeightsStore[0][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_62;WeightsStore[0][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_63;WeightsStore[0][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_64;WeightsStore[0][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_65;WeightsStore[0][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_66;WeightsStore[0][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_67;WeightsStore[0][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_68;WeightsStore[0][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_69;WeightsStore[0][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_70;WeightsStore[0][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_71;WeightsStore[0][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_72;WeightsStore[0][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_73;WeightsStore[0][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_74;WeightsStore[0][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_75;WeightsStore[0][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_76;WeightsStore[0][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_77;WeightsStore[0][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_78;WeightsStore[0][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_79;WeightsStore[0][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_80;WeightsStore[0][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_81;WeightsStore[0][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_82;WeightsStore[0][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_83;WeightsStore[0][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_84;WeightsStore[0][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_85;WeightsStore[0][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_86;WeightsStore[0][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_87;WeightsStore[0][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_88;WeightsStore[0][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_89;WeightsStore[0][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_90;WeightsStore[0][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_91;WeightsStore[0][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_92;WeightsStore[0][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_93;WeightsStore[0][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_94;WeightsStore[0][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_95;WeightsStore[0][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_96;WeightsStore[0][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_97;WeightsStore[0][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_98;WeightsStore[0][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_99;WeightsStore[0][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_100;WeightsStore[0][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_101;WeightsStore[0][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_102;WeightsStore[0][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_103;WeightsStore[0][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_104;WeightsStore[0][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_105;WeightsStore[0][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_106;WeightsStore[0][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_107;WeightsStore[0][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_108;WeightsStore[0][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_109;WeightsStore[0][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_110;WeightsStore[0][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_111;WeightsStore[0][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_112;WeightsStore[0][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_113;WeightsStore[0][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_114;WeightsStore[0][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_115;WeightsStore[0][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_116;WeightsStore[0][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_117;WeightsStore[0][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_118;WeightsStore[0][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_119;WeightsStore[0][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_120;WeightsStore[0][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_121;WeightsStore[0][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_122;WeightsStore[0][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_123;WeightsStore[0][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_124;WeightsStore[0][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_125;WeightsStore[0][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_126;WeightsStore[0][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_127;WeightsStore[0][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_128;WeightsStore[0][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_129;WeightsStore[0][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_130;WeightsStore[0][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_131;WeightsStore[0][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_132;WeightsStore[0][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_133;WeightsStore[0][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_134;WeightsStore[0][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_135;WeightsStore[0][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_136;WeightsStore[0][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_137;WeightsStore[0][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_138;WeightsStore[0][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_139;WeightsStore[0][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_140;WeightsStore[0][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_141;WeightsStore[0][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_142;WeightsStore[0][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_143;WeightsStore[0][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_144;WeightsStore[0][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_145;WeightsStore[0][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_146;WeightsStore[0][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_147;WeightsStore[0][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_148;WeightsStore[0][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_149;WeightsStore[0][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_150;WeightsStore[0][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_151;WeightsStore[0][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_152;WeightsStore[0][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_153;WeightsStore[0][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_154;WeightsStore[0][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_155;WeightsStore[0][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_156;WeightsStore[0][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_157;WeightsStore[0][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_158;WeightsStore[0][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_159;WeightsStore[0][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_160;WeightsStore[0][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_161;WeightsStore[0][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_162;WeightsStore[0][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_163;WeightsStore[0][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_164;WeightsStore[0][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_165;WeightsStore[0][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_166;WeightsStore[0][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_167;WeightsStore[0][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_168;WeightsStore[0][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_169;WeightsStore[0][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_170;WeightsStore[0][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_171;WeightsStore[0][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_172;WeightsStore[0][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_173;WeightsStore[0][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_174;WeightsStore[0][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_175;WeightsStore[0][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_176;WeightsStore[0][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_177;WeightsStore[0][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_178;WeightsStore[0][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_179;WeightsStore[0][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_180;WeightsStore[0][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_181;WeightsStore[0][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_182;WeightsStore[0][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_183;WeightsStore[0][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_184;WeightsStore[0][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_185;WeightsStore[0][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_186;WeightsStore[0][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_187;WeightsStore[0][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_188;WeightsStore[0][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_189;WeightsStore[0][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_190;WeightsStore[0][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_191;WeightsStore[0][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_192;WeightsStore[0][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_193;WeightsStore[0][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_194;WeightsStore[0][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_195;WeightsStore[0][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_196;WeightsStore[0][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_197;WeightsStore[0][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_198;WeightsStore[0][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_199;WeightsStore[0][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_200;WeightsStore[0][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_201;WeightsStore[0][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_202;WeightsStore[0][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_203;WeightsStore[0][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_204;WeightsStore[0][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_205;WeightsStore[0][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_206;WeightsStore[0][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_207;WeightsStore[0][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_208;WeightsStore[0][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_209;WeightsStore[0][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_210;WeightsStore[0][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_211;WeightsStore[0][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_212;WeightsStore[0][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_213;WeightsStore[0][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_214;WeightsStore[0][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_215;WeightsStore[0][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_216;WeightsStore[0][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_217;WeightsStore[0][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_218;WeightsStore[0][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_219;WeightsStore[0][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_220;WeightsStore[0][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_221;WeightsStore[0][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_222;WeightsStore[0][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_223;WeightsStore[0][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_224;WeightsStore[0][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_225;WeightsStore[0][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_226;WeightsStore[0][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_227;WeightsStore[0][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_228;WeightsStore[0][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_229;WeightsStore[0][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_230;WeightsStore[0][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_231;WeightsStore[0][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_232;WeightsStore[0][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_233;WeightsStore[0][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_234;WeightsStore[0][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_235;WeightsStore[0][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_236;WeightsStore[0][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_237;WeightsStore[0][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_238;WeightsStore[0][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_239;WeightsStore[0][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_240;WeightsStore[0][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_241;WeightsStore[0][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_242;WeightsStore[0][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_243;WeightsStore[0][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_244;WeightsStore[0][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_245;WeightsStore[0][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_246;WeightsStore[0][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_247;WeightsStore[0][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_248;WeightsStore[0][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_249;WeightsStore[0][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_250;WeightsStore[0][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_251;WeightsStore[0][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_252;WeightsStore[0][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_253;WeightsStore[0][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_254;WeightsStore[0][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_255;WeightsStore[0][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_256;WeightsStore[0][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_257;WeightsStore[0][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_258;WeightsStore[0][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_259;WeightsStore[0][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_260;WeightsStore[0][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_261;WeightsStore[0][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_262;WeightsStore[0][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_263;WeightsStore[0][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_264;WeightsStore[0][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_265;WeightsStore[0][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_266;WeightsStore[0][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_267;WeightsStore[0][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_268;WeightsStore[0][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_269;WeightsStore[0][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_270;WeightsStore[0][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_271;WeightsStore[0][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_272;WeightsStore[0][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_273;WeightsStore[0][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_274;WeightsStore[0][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_275;WeightsStore[0][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_276;WeightsStore[0][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_277;WeightsStore[0][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_278;WeightsStore[0][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_279;WeightsStore[0][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_280;WeightsStore[0][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_281;WeightsStore[0][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_282;WeightsStore[0][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_283;WeightsStore[0][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_284;WeightsStore[0][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_285;WeightsStore[0][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_286;WeightsStore[0][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_287;WeightsStore[0][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_288;WeightsStore[0][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_289;WeightsStore[0][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_290;WeightsStore[0][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_291;WeightsStore[0][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_292;WeightsStore[0][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_293;WeightsStore[0][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_294;WeightsStore[0][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_295;WeightsStore[0][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_296;WeightsStore[0][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_297;WeightsStore[0][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_298;WeightsStore[0][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_299;WeightsStore[0][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_300;WeightsStore[0][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_301;WeightsStore[0][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_302;WeightsStore[0][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_303;WeightsStore[0][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_304;WeightsStore[0][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_305;WeightsStore[0][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_306;WeightsStore[0][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_307;WeightsStore[0][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_308;WeightsStore[0][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_309;WeightsStore[0][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_310;WeightsStore[0][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_311;WeightsStore[0][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_312;WeightsStore[0][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_313;WeightsStore[0][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_314;WeightsStore[0][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_315;WeightsStore[0][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_316;WeightsStore[0][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_317;WeightsStore[0][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_318;WeightsStore[0][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_319;WeightsStore[0][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_320;WeightsStore[0][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_321;WeightsStore[0][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_322;WeightsStore[0][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_323;WeightsStore[0][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_324;WeightsStore[0][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_325;WeightsStore[0][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_326;WeightsStore[0][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_327;WeightsStore[0][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_328;WeightsStore[0][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_329;WeightsStore[0][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_330;WeightsStore[0][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_331;WeightsStore[0][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_332;WeightsStore[0][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_333;WeightsStore[0][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_334;WeightsStore[0][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_335;WeightsStore[0][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_336;WeightsStore[0][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_337;WeightsStore[0][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_338;WeightsStore[0][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_339;WeightsStore[0][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_340;WeightsStore[0][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_341;WeightsStore[0][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_342;WeightsStore[0][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_343;WeightsStore[0][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_344;WeightsStore[0][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_345;WeightsStore[0][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_346;WeightsStore[0][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_347;WeightsStore[0][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_348;WeightsStore[0][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_349;WeightsStore[0][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_350;WeightsStore[0][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_351;WeightsStore[0][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_352;WeightsStore[0][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_353;WeightsStore[0][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_354;WeightsStore[0][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_355;WeightsStore[0][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_356;WeightsStore[0][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_357;WeightsStore[0][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_358;WeightsStore[0][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_359;WeightsStore[0][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_360;WeightsStore[0][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_361;WeightsStore[0][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_362;WeightsStore[0][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_363;WeightsStore[0][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_364;WeightsStore[0][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_365;WeightsStore[0][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_366;WeightsStore[0][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_367;WeightsStore[0][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_368;WeightsStore[0][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_369;WeightsStore[0][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_370;WeightsStore[0][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_371;WeightsStore[0][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_372;WeightsStore[0][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_373;WeightsStore[0][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_374;WeightsStore[0][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_375;WeightsStore[0][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_376;WeightsStore[0][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_377;WeightsStore[0][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_378;WeightsStore[0][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_379;WeightsStore[0][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_380;WeightsStore[0][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_381;WeightsStore[0][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_382;WeightsStore[0][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_383;WeightsStore[0][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_384;WeightsStore[0][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_385;WeightsStore[0][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_386;WeightsStore[0][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_387;WeightsStore[0][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_388;WeightsStore[0][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_389;WeightsStore[0][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_390;WeightsStore[0][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_391;WeightsStore[0][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_392;WeightsStore[0][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_393;WeightsStore[0][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_394;WeightsStore[0][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_395;WeightsStore[0][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_396;WeightsStore[0][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_397;WeightsStore[0][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_398;WeightsStore[0][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_399;WeightsStore[0][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_400;WeightsStore[0][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_401;WeightsStore[0][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_402;WeightsStore[0][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_403;WeightsStore[0][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_404;WeightsStore[0][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_405;WeightsStore[0][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_406;WeightsStore[0][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_407;WeightsStore[0][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_408;WeightsStore[0][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_409;WeightsStore[0][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_410;WeightsStore[0][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_411;WeightsStore[0][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_412;WeightsStore[0][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_413;WeightsStore[0][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_414;WeightsStore[0][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_415;WeightsStore[0][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_416;WeightsStore[0][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_417;WeightsStore[0][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_418;WeightsStore[0][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_419;WeightsStore[0][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_420;WeightsStore[0][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_421;WeightsStore[0][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_422;WeightsStore[0][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_423;WeightsStore[0][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_424;WeightsStore[0][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_425;WeightsStore[0][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_426;WeightsStore[0][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_427;WeightsStore[0][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_428;WeightsStore[0][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_429;WeightsStore[0][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_430;WeightsStore[0][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_431;WeightsStore[0][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_432;WeightsStore[0][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_433;WeightsStore[0][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_434;WeightsStore[0][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_435;WeightsStore[0][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_436;WeightsStore[0][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_437;WeightsStore[0][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_438;WeightsStore[0][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_439;WeightsStore[0][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_440;WeightsStore[0][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_441;WeightsStore[0][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_442;WeightsStore[0][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_443;WeightsStore[0][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_444;WeightsStore[0][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_445;WeightsStore[0][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_446;WeightsStore[0][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_447;WeightsStore[0][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_448;WeightsStore[0][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_449;WeightsStore[0][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_450;WeightsStore[0][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_451;WeightsStore[0][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_452;WeightsStore[0][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_453;WeightsStore[0][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_454;WeightsStore[0][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_455;WeightsStore[0][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_456;WeightsStore[0][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_457;WeightsStore[0][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_458;WeightsStore[0][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_459;WeightsStore[0][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_460;WeightsStore[0][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_461;WeightsStore[0][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_462;WeightsStore[0][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_463;WeightsStore[0][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_464;WeightsStore[0][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_465;WeightsStore[0][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_466;WeightsStore[0][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_467;WeightsStore[0][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_468;WeightsStore[0][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_469;WeightsStore[0][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_470;WeightsStore[0][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_471;WeightsStore[0][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_472;WeightsStore[0][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_473;WeightsStore[0][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_474;WeightsStore[0][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_475;WeightsStore[0][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_476;WeightsStore[0][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_477;WeightsStore[0][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_478;WeightsStore[0][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_479;WeightsStore[0][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_480;WeightsStore[0][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_481;WeightsStore[0][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_482;WeightsStore[0][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_483;WeightsStore[0][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_484;WeightsStore[0][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_485;WeightsStore[0][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_486;WeightsStore[0][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_487;WeightsStore[0][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_488;WeightsStore[0][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_489;WeightsStore[0][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_490;WeightsStore[0][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_491;WeightsStore[0][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_492;WeightsStore[0][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_493;WeightsStore[0][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_494;WeightsStore[0][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_495;WeightsStore[0][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_496;WeightsStore[0][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_497;WeightsStore[0][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_498;WeightsStore[0][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_499;WeightsStore[0][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_500;WeightsStore[0][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_501;WeightsStore[0][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_502;WeightsStore[0][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_503;WeightsStore[0][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_504;WeightsStore[0][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_505;WeightsStore[0][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_506;WeightsStore[0][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_507;WeightsStore[0][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_508;WeightsStore[0][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_509;WeightsStore[0][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_510;WeightsStore[0][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_511;WeightsStore[0][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_512;WeightsStore[0][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_513;WeightsStore[0][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_514;WeightsStore[0][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_515;WeightsStore[0][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_516;WeightsStore[0][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_517;WeightsStore[0][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_518;WeightsStore[0][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_519;WeightsStore[0][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_520;WeightsStore[0][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_521;WeightsStore[0][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_522;WeightsStore[0][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_523;WeightsStore[0][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_524;WeightsStore[0][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_525;WeightsStore[0][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_526;WeightsStore[0][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_527;WeightsStore[0][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_528;WeightsStore[0][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_529;WeightsStore[0][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_530;WeightsStore[0][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_531;WeightsStore[0][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_532;WeightsStore[0][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_533;WeightsStore[0][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_534;WeightsStore[0][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_535;WeightsStore[0][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_536;WeightsStore[0][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_537;WeightsStore[0][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_538;WeightsStore[0][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_539;WeightsStore[0][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_540;WeightsStore[0][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_541;WeightsStore[0][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_542;WeightsStore[0][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_543;WeightsStore[0][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_544;WeightsStore[0][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_545;WeightsStore[0][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_546;WeightsStore[0][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_547;WeightsStore[0][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_548;WeightsStore[0][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_549;WeightsStore[0][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_550;WeightsStore[0][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_551;WeightsStore[0][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_552;WeightsStore[0][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_553;WeightsStore[0][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_554;WeightsStore[0][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_555;WeightsStore[0][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_556;WeightsStore[0][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_557;WeightsStore[0][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_558;WeightsStore[0][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_559;WeightsStore[0][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_560;WeightsStore[0][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_561;WeightsStore[0][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_562;WeightsStore[0][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_563;WeightsStore[0][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_564;WeightsStore[0][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_565;WeightsStore[0][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_566;WeightsStore[0][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_567;WeightsStore[0][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_568;WeightsStore[0][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_569;WeightsStore[0][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_570;WeightsStore[0][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_571;WeightsStore[0][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_572;WeightsStore[0][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_573;WeightsStore[0][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_574;WeightsStore[0][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_575;WeightsStore[0][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_576;WeightsStore[0][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_577;WeightsStore[0][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_578;WeightsStore[0][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_579;WeightsStore[0][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_580;WeightsStore[0][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_581;WeightsStore[0][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_582;WeightsStore[0][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_583;WeightsStore[0][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_584;WeightsStore[0][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_585;WeightsStore[0][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_586;WeightsStore[0][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_587;WeightsStore[0][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_588;WeightsStore[0][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_589;WeightsStore[0][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_590;WeightsStore[0][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_591;WeightsStore[0][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_592;WeightsStore[0][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_593;WeightsStore[0][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_594;WeightsStore[0][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_595;WeightsStore[0][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_596;WeightsStore[0][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_597;WeightsStore[0][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_598;WeightsStore[0][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_599;WeightsStore[0][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_600;WeightsStore[0][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_601;WeightsStore[0][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_602;WeightsStore[0][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_603;WeightsStore[0][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_604;WeightsStore[0][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_605;WeightsStore[0][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_606;WeightsStore[0][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_607;WeightsStore[0][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_608;WeightsStore[0][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_609;WeightsStore[0][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_610;WeightsStore[0][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_611;WeightsStore[0][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_612;WeightsStore[0][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_613;WeightsStore[0][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_614;WeightsStore[0][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_615;WeightsStore[0][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_616;WeightsStore[0][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_617;WeightsStore[0][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_618;WeightsStore[0][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_619;WeightsStore[0][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_620;WeightsStore[0][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_621;WeightsStore[0][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_622;WeightsStore[0][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_623;WeightsStore[0][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_624;WeightsStore[0][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_625;WeightsStore[0][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_626;WeightsStore[0][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_627;WeightsStore[0][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_628;WeightsStore[0][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_629;WeightsStore[0][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_630;WeightsStore[0][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_631;WeightsStore[0][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_632;WeightsStore[0][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_633;WeightsStore[0][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_634;WeightsStore[0][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_635;WeightsStore[0][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_636;WeightsStore[0][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_637;WeightsStore[0][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_638;WeightsStore[0][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_639;WeightsStore[0][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_640;WeightsStore[0][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_641;WeightsStore[0][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_642;WeightsStore[0][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_643;WeightsStore[0][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_644;WeightsStore[0][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_645;WeightsStore[0][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_646;WeightsStore[0][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_647;WeightsStore[0][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_648;WeightsStore[0][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_649;WeightsStore[0][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_650;WeightsStore[0][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_651;WeightsStore[0][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_652;WeightsStore[0][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_653;WeightsStore[0][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_654;WeightsStore[0][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_655;WeightsStore[0][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_656;WeightsStore[0][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_657;WeightsStore[0][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_658;WeightsStore[0][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_659;WeightsStore[0][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_660;WeightsStore[0][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_661;WeightsStore[0][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_662;WeightsStore[0][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_663;WeightsStore[0][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_664;WeightsStore[0][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_665;WeightsStore[0][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_666;WeightsStore[0][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_667;WeightsStore[0][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_668;WeightsStore[0][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_669;WeightsStore[0][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_670;WeightsStore[0][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_671;WeightsStore[0][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_672;WeightsStore[0][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_673;WeightsStore[0][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_674;WeightsStore[0][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_675;WeightsStore[0][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_676;WeightsStore[0][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_677;WeightsStore[0][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_678;WeightsStore[0][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_679;WeightsStore[0][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_680;WeightsStore[0][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_681;WeightsStore[0][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_682;WeightsStore[0][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_683;WeightsStore[0][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_684;WeightsStore[0][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_685;WeightsStore[0][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_686;WeightsStore[0][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_687;WeightsStore[0][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_688;WeightsStore[0][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_689;WeightsStore[0][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_690;WeightsStore[0][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_691;WeightsStore[0][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_692;WeightsStore[0][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_693;WeightsStore[0][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_694;WeightsStore[0][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_695;WeightsStore[0][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_696;WeightsStore[0][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_697;WeightsStore[0][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_698;WeightsStore[0][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_699;WeightsStore[0][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_700;WeightsStore[0][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_701;WeightsStore[0][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_702;WeightsStore[0][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_703;WeightsStore[0][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_704;WeightsStore[0][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_705;WeightsStore[0][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_706;WeightsStore[0][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_707;WeightsStore[0][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_708;WeightsStore[0][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_709;WeightsStore[0][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_710;WeightsStore[0][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_711;WeightsStore[0][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_712;WeightsStore[0][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_713;WeightsStore[0][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_714;WeightsStore[0][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_715;WeightsStore[0][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_716;WeightsStore[0][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_717;WeightsStore[0][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_718;WeightsStore[0][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_719;WeightsStore[0][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_720;WeightsStore[0][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_721;WeightsStore[0][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_722;WeightsStore[0][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_723;WeightsStore[0][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_724;WeightsStore[0][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_725;WeightsStore[0][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_726;WeightsStore[0][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_727;WeightsStore[0][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_728;WeightsStore[0][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_729;WeightsStore[0][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_730;WeightsStore[0][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_731;WeightsStore[0][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_732;WeightsStore[0][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_733;WeightsStore[0][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_734;WeightsStore[0][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_735;WeightsStore[0][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_736;WeightsStore[0][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_737;WeightsStore[0][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_738;WeightsStore[0][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_739;WeightsStore[0][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_740;WeightsStore[0][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_741;WeightsStore[0][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_742;WeightsStore[0][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_743;WeightsStore[0][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_744;WeightsStore[0][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_745;WeightsStore[0][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_746;WeightsStore[0][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_747;WeightsStore[0][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_748;WeightsStore[0][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_749;WeightsStore[0][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_750;WeightsStore[0][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_751;WeightsStore[0][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_752;WeightsStore[0][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_753;WeightsStore[0][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_754;WeightsStore[0][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_755;WeightsStore[0][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_756;WeightsStore[0][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_757;WeightsStore[0][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_758;WeightsStore[0][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_759;WeightsStore[0][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_760;WeightsStore[0][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_761;WeightsStore[0][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_762;WeightsStore[0][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_763;WeightsStore[0][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_764;WeightsStore[0][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_765;WeightsStore[0][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_766;WeightsStore[0][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_767;WeightsStore[0][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_768;WeightsStore[0][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_769;WeightsStore[0][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_770;WeightsStore[0][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_771;WeightsStore[0][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_772;WeightsStore[0][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_773;WeightsStore[0][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_774;WeightsStore[0][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_775;WeightsStore[0][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_776;WeightsStore[0][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_777;WeightsStore[0][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_778;WeightsStore[0][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_779;WeightsStore[0][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_780;WeightsStore[0][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_781;WeightsStore[0][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_782;WeightsStore[0][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_783;WeightsStore[0][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_0_784;WeightsStore[1][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_0;WeightsStore[1][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_1;WeightsStore[1][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_2;WeightsStore[1][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_3;WeightsStore[1][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_4;WeightsStore[1][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_5;WeightsStore[1][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_6;WeightsStore[1][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_7;WeightsStore[1][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_8;WeightsStore[1][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_9;WeightsStore[1][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_10;WeightsStore[1][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_11;WeightsStore[1][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_12;WeightsStore[1][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_13;WeightsStore[1][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_14;WeightsStore[1][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_15;WeightsStore[1][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_16;WeightsStore[1][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_17;WeightsStore[1][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_18;WeightsStore[1][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_19;WeightsStore[1][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_20;WeightsStore[1][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_21;WeightsStore[1][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_22;WeightsStore[1][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_23;WeightsStore[1][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_24;WeightsStore[1][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_25;WeightsStore[1][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_26;WeightsStore[1][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_27;WeightsStore[1][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_28;WeightsStore[1][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_29;WeightsStore[1][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_30;WeightsStore[1][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_31;WeightsStore[1][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_32;WeightsStore[1][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_33;WeightsStore[1][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_34;WeightsStore[1][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_35;WeightsStore[1][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_36;WeightsStore[1][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_37;WeightsStore[1][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_38;WeightsStore[1][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_39;WeightsStore[1][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_40;WeightsStore[1][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_41;WeightsStore[1][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_42;WeightsStore[1][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_43;WeightsStore[1][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_44;WeightsStore[1][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_45;WeightsStore[1][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_46;WeightsStore[1][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_47;WeightsStore[1][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_48;WeightsStore[1][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_49;WeightsStore[1][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_50;WeightsStore[1][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_51;WeightsStore[1][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_52;WeightsStore[1][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_53;WeightsStore[1][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_54;WeightsStore[1][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_55;WeightsStore[1][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_56;WeightsStore[1][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_57;WeightsStore[1][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_58;WeightsStore[1][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_59;WeightsStore[1][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_60;WeightsStore[1][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_61;WeightsStore[1][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_62;WeightsStore[1][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_63;WeightsStore[1][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_64;WeightsStore[1][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_65;WeightsStore[1][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_66;WeightsStore[1][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_67;WeightsStore[1][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_68;WeightsStore[1][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_69;WeightsStore[1][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_70;WeightsStore[1][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_71;WeightsStore[1][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_72;WeightsStore[1][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_73;WeightsStore[1][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_74;WeightsStore[1][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_75;WeightsStore[1][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_76;WeightsStore[1][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_77;WeightsStore[1][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_78;WeightsStore[1][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_79;WeightsStore[1][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_80;WeightsStore[1][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_81;WeightsStore[1][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_82;WeightsStore[1][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_83;WeightsStore[1][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_84;WeightsStore[1][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_85;WeightsStore[1][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_86;WeightsStore[1][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_87;WeightsStore[1][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_88;WeightsStore[1][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_89;WeightsStore[1][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_90;WeightsStore[1][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_91;WeightsStore[1][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_92;WeightsStore[1][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_93;WeightsStore[1][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_94;WeightsStore[1][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_95;WeightsStore[1][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_96;WeightsStore[1][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_97;WeightsStore[1][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_98;WeightsStore[1][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_99;WeightsStore[1][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_100;WeightsStore[1][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_101;WeightsStore[1][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_102;WeightsStore[1][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_103;WeightsStore[1][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_104;WeightsStore[1][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_105;WeightsStore[1][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_106;WeightsStore[1][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_107;WeightsStore[1][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_108;WeightsStore[1][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_109;WeightsStore[1][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_110;WeightsStore[1][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_111;WeightsStore[1][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_112;WeightsStore[1][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_113;WeightsStore[1][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_114;WeightsStore[1][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_115;WeightsStore[1][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_116;WeightsStore[1][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_117;WeightsStore[1][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_118;WeightsStore[1][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_119;WeightsStore[1][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_120;WeightsStore[1][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_121;WeightsStore[1][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_122;WeightsStore[1][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_123;WeightsStore[1][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_124;WeightsStore[1][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_125;WeightsStore[1][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_126;WeightsStore[1][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_127;WeightsStore[1][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_128;WeightsStore[1][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_129;WeightsStore[1][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_130;WeightsStore[1][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_131;WeightsStore[1][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_132;WeightsStore[1][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_133;WeightsStore[1][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_134;WeightsStore[1][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_135;WeightsStore[1][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_136;WeightsStore[1][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_137;WeightsStore[1][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_138;WeightsStore[1][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_139;WeightsStore[1][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_140;WeightsStore[1][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_141;WeightsStore[1][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_142;WeightsStore[1][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_143;WeightsStore[1][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_144;WeightsStore[1][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_145;WeightsStore[1][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_146;WeightsStore[1][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_147;WeightsStore[1][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_148;WeightsStore[1][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_149;WeightsStore[1][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_150;WeightsStore[1][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_151;WeightsStore[1][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_152;WeightsStore[1][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_153;WeightsStore[1][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_154;WeightsStore[1][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_155;WeightsStore[1][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_156;WeightsStore[1][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_157;WeightsStore[1][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_158;WeightsStore[1][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_159;WeightsStore[1][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_160;WeightsStore[1][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_161;WeightsStore[1][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_162;WeightsStore[1][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_163;WeightsStore[1][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_164;WeightsStore[1][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_165;WeightsStore[1][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_166;WeightsStore[1][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_167;WeightsStore[1][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_168;WeightsStore[1][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_169;WeightsStore[1][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_170;WeightsStore[1][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_171;WeightsStore[1][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_172;WeightsStore[1][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_173;WeightsStore[1][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_174;WeightsStore[1][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_175;WeightsStore[1][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_176;WeightsStore[1][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_177;WeightsStore[1][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_178;WeightsStore[1][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_179;WeightsStore[1][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_180;WeightsStore[1][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_181;WeightsStore[1][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_182;WeightsStore[1][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_183;WeightsStore[1][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_184;WeightsStore[1][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_185;WeightsStore[1][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_186;WeightsStore[1][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_187;WeightsStore[1][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_188;WeightsStore[1][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_189;WeightsStore[1][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_190;WeightsStore[1][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_191;WeightsStore[1][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_192;WeightsStore[1][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_193;WeightsStore[1][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_194;WeightsStore[1][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_195;WeightsStore[1][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_196;WeightsStore[1][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_197;WeightsStore[1][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_198;WeightsStore[1][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_199;WeightsStore[1][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_200;WeightsStore[1][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_201;WeightsStore[1][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_202;WeightsStore[1][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_203;WeightsStore[1][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_204;WeightsStore[1][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_205;WeightsStore[1][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_206;WeightsStore[1][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_207;WeightsStore[1][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_208;WeightsStore[1][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_209;WeightsStore[1][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_210;WeightsStore[1][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_211;WeightsStore[1][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_212;WeightsStore[1][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_213;WeightsStore[1][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_214;WeightsStore[1][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_215;WeightsStore[1][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_216;WeightsStore[1][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_217;WeightsStore[1][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_218;WeightsStore[1][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_219;WeightsStore[1][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_220;WeightsStore[1][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_221;WeightsStore[1][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_222;WeightsStore[1][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_223;WeightsStore[1][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_224;WeightsStore[1][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_225;WeightsStore[1][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_226;WeightsStore[1][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_227;WeightsStore[1][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_228;WeightsStore[1][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_229;WeightsStore[1][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_230;WeightsStore[1][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_231;WeightsStore[1][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_232;WeightsStore[1][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_233;WeightsStore[1][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_234;WeightsStore[1][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_235;WeightsStore[1][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_236;WeightsStore[1][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_237;WeightsStore[1][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_238;WeightsStore[1][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_239;WeightsStore[1][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_240;WeightsStore[1][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_241;WeightsStore[1][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_242;WeightsStore[1][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_243;WeightsStore[1][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_244;WeightsStore[1][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_245;WeightsStore[1][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_246;WeightsStore[1][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_247;WeightsStore[1][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_248;WeightsStore[1][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_249;WeightsStore[1][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_250;WeightsStore[1][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_251;WeightsStore[1][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_252;WeightsStore[1][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_253;WeightsStore[1][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_254;WeightsStore[1][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_255;WeightsStore[1][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_256;WeightsStore[1][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_257;WeightsStore[1][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_258;WeightsStore[1][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_259;WeightsStore[1][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_260;WeightsStore[1][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_261;WeightsStore[1][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_262;WeightsStore[1][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_263;WeightsStore[1][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_264;WeightsStore[1][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_265;WeightsStore[1][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_266;WeightsStore[1][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_267;WeightsStore[1][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_268;WeightsStore[1][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_269;WeightsStore[1][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_270;WeightsStore[1][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_271;WeightsStore[1][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_272;WeightsStore[1][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_273;WeightsStore[1][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_274;WeightsStore[1][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_275;WeightsStore[1][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_276;WeightsStore[1][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_277;WeightsStore[1][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_278;WeightsStore[1][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_279;WeightsStore[1][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_280;WeightsStore[1][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_281;WeightsStore[1][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_282;WeightsStore[1][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_283;WeightsStore[1][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_284;WeightsStore[1][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_285;WeightsStore[1][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_286;WeightsStore[1][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_287;WeightsStore[1][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_288;WeightsStore[1][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_289;WeightsStore[1][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_290;WeightsStore[1][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_291;WeightsStore[1][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_292;WeightsStore[1][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_293;WeightsStore[1][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_294;WeightsStore[1][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_295;WeightsStore[1][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_296;WeightsStore[1][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_297;WeightsStore[1][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_298;WeightsStore[1][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_299;WeightsStore[1][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_300;WeightsStore[1][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_301;WeightsStore[1][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_302;WeightsStore[1][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_303;WeightsStore[1][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_304;WeightsStore[1][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_305;WeightsStore[1][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_306;WeightsStore[1][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_307;WeightsStore[1][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_308;WeightsStore[1][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_309;WeightsStore[1][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_310;WeightsStore[1][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_311;WeightsStore[1][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_312;WeightsStore[1][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_313;WeightsStore[1][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_314;WeightsStore[1][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_315;WeightsStore[1][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_316;WeightsStore[1][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_317;WeightsStore[1][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_318;WeightsStore[1][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_319;WeightsStore[1][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_320;WeightsStore[1][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_321;WeightsStore[1][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_322;WeightsStore[1][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_323;WeightsStore[1][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_324;WeightsStore[1][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_325;WeightsStore[1][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_326;WeightsStore[1][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_327;WeightsStore[1][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_328;WeightsStore[1][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_329;WeightsStore[1][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_330;WeightsStore[1][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_331;WeightsStore[1][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_332;WeightsStore[1][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_333;WeightsStore[1][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_334;WeightsStore[1][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_335;WeightsStore[1][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_336;WeightsStore[1][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_337;WeightsStore[1][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_338;WeightsStore[1][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_339;WeightsStore[1][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_340;WeightsStore[1][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_341;WeightsStore[1][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_342;WeightsStore[1][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_343;WeightsStore[1][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_344;WeightsStore[1][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_345;WeightsStore[1][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_346;WeightsStore[1][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_347;WeightsStore[1][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_348;WeightsStore[1][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_349;WeightsStore[1][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_350;WeightsStore[1][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_351;WeightsStore[1][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_352;WeightsStore[1][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_353;WeightsStore[1][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_354;WeightsStore[1][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_355;WeightsStore[1][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_356;WeightsStore[1][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_357;WeightsStore[1][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_358;WeightsStore[1][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_359;WeightsStore[1][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_360;WeightsStore[1][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_361;WeightsStore[1][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_362;WeightsStore[1][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_363;WeightsStore[1][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_364;WeightsStore[1][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_365;WeightsStore[1][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_366;WeightsStore[1][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_367;WeightsStore[1][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_368;WeightsStore[1][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_369;WeightsStore[1][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_370;WeightsStore[1][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_371;WeightsStore[1][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_372;WeightsStore[1][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_373;WeightsStore[1][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_374;WeightsStore[1][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_375;WeightsStore[1][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_376;WeightsStore[1][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_377;WeightsStore[1][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_378;WeightsStore[1][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_379;WeightsStore[1][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_380;WeightsStore[1][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_381;WeightsStore[1][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_382;WeightsStore[1][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_383;WeightsStore[1][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_384;WeightsStore[1][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_385;WeightsStore[1][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_386;WeightsStore[1][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_387;WeightsStore[1][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_388;WeightsStore[1][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_389;WeightsStore[1][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_390;WeightsStore[1][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_391;WeightsStore[1][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_392;WeightsStore[1][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_393;WeightsStore[1][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_394;WeightsStore[1][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_395;WeightsStore[1][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_396;WeightsStore[1][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_397;WeightsStore[1][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_398;WeightsStore[1][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_399;WeightsStore[1][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_400;WeightsStore[1][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_401;WeightsStore[1][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_402;WeightsStore[1][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_403;WeightsStore[1][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_404;WeightsStore[1][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_405;WeightsStore[1][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_406;WeightsStore[1][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_407;WeightsStore[1][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_408;WeightsStore[1][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_409;WeightsStore[1][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_410;WeightsStore[1][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_411;WeightsStore[1][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_412;WeightsStore[1][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_413;WeightsStore[1][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_414;WeightsStore[1][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_415;WeightsStore[1][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_416;WeightsStore[1][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_417;WeightsStore[1][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_418;WeightsStore[1][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_419;WeightsStore[1][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_420;WeightsStore[1][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_421;WeightsStore[1][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_422;WeightsStore[1][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_423;WeightsStore[1][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_424;WeightsStore[1][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_425;WeightsStore[1][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_426;WeightsStore[1][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_427;WeightsStore[1][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_428;WeightsStore[1][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_429;WeightsStore[1][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_430;WeightsStore[1][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_431;WeightsStore[1][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_432;WeightsStore[1][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_433;WeightsStore[1][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_434;WeightsStore[1][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_435;WeightsStore[1][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_436;WeightsStore[1][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_437;WeightsStore[1][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_438;WeightsStore[1][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_439;WeightsStore[1][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_440;WeightsStore[1][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_441;WeightsStore[1][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_442;WeightsStore[1][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_443;WeightsStore[1][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_444;WeightsStore[1][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_445;WeightsStore[1][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_446;WeightsStore[1][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_447;WeightsStore[1][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_448;WeightsStore[1][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_449;WeightsStore[1][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_450;WeightsStore[1][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_451;WeightsStore[1][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_452;WeightsStore[1][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_453;WeightsStore[1][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_454;WeightsStore[1][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_455;WeightsStore[1][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_456;WeightsStore[1][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_457;WeightsStore[1][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_458;WeightsStore[1][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_459;WeightsStore[1][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_460;WeightsStore[1][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_461;WeightsStore[1][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_462;WeightsStore[1][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_463;WeightsStore[1][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_464;WeightsStore[1][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_465;WeightsStore[1][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_466;WeightsStore[1][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_467;WeightsStore[1][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_468;WeightsStore[1][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_469;WeightsStore[1][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_470;WeightsStore[1][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_471;WeightsStore[1][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_472;WeightsStore[1][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_473;WeightsStore[1][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_474;WeightsStore[1][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_475;WeightsStore[1][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_476;WeightsStore[1][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_477;WeightsStore[1][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_478;WeightsStore[1][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_479;WeightsStore[1][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_480;WeightsStore[1][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_481;WeightsStore[1][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_482;WeightsStore[1][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_483;WeightsStore[1][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_484;WeightsStore[1][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_485;WeightsStore[1][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_486;WeightsStore[1][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_487;WeightsStore[1][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_488;WeightsStore[1][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_489;WeightsStore[1][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_490;WeightsStore[1][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_491;WeightsStore[1][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_492;WeightsStore[1][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_493;WeightsStore[1][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_494;WeightsStore[1][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_495;WeightsStore[1][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_496;WeightsStore[1][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_497;WeightsStore[1][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_498;WeightsStore[1][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_499;WeightsStore[1][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_500;WeightsStore[1][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_501;WeightsStore[1][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_502;WeightsStore[1][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_503;WeightsStore[1][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_504;WeightsStore[1][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_505;WeightsStore[1][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_506;WeightsStore[1][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_507;WeightsStore[1][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_508;WeightsStore[1][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_509;WeightsStore[1][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_510;WeightsStore[1][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_511;WeightsStore[1][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_512;WeightsStore[1][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_513;WeightsStore[1][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_514;WeightsStore[1][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_515;WeightsStore[1][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_516;WeightsStore[1][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_517;WeightsStore[1][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_518;WeightsStore[1][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_519;WeightsStore[1][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_520;WeightsStore[1][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_521;WeightsStore[1][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_522;WeightsStore[1][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_523;WeightsStore[1][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_524;WeightsStore[1][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_525;WeightsStore[1][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_526;WeightsStore[1][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_527;WeightsStore[1][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_528;WeightsStore[1][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_529;WeightsStore[1][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_530;WeightsStore[1][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_531;WeightsStore[1][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_532;WeightsStore[1][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_533;WeightsStore[1][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_534;WeightsStore[1][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_535;WeightsStore[1][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_536;WeightsStore[1][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_537;WeightsStore[1][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_538;WeightsStore[1][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_539;WeightsStore[1][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_540;WeightsStore[1][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_541;WeightsStore[1][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_542;WeightsStore[1][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_543;WeightsStore[1][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_544;WeightsStore[1][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_545;WeightsStore[1][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_546;WeightsStore[1][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_547;WeightsStore[1][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_548;WeightsStore[1][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_549;WeightsStore[1][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_550;WeightsStore[1][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_551;WeightsStore[1][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_552;WeightsStore[1][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_553;WeightsStore[1][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_554;WeightsStore[1][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_555;WeightsStore[1][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_556;WeightsStore[1][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_557;WeightsStore[1][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_558;WeightsStore[1][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_559;WeightsStore[1][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_560;WeightsStore[1][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_561;WeightsStore[1][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_562;WeightsStore[1][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_563;WeightsStore[1][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_564;WeightsStore[1][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_565;WeightsStore[1][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_566;WeightsStore[1][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_567;WeightsStore[1][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_568;WeightsStore[1][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_569;WeightsStore[1][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_570;WeightsStore[1][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_571;WeightsStore[1][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_572;WeightsStore[1][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_573;WeightsStore[1][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_574;WeightsStore[1][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_575;WeightsStore[1][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_576;WeightsStore[1][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_577;WeightsStore[1][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_578;WeightsStore[1][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_579;WeightsStore[1][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_580;WeightsStore[1][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_581;WeightsStore[1][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_582;WeightsStore[1][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_583;WeightsStore[1][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_584;WeightsStore[1][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_585;WeightsStore[1][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_586;WeightsStore[1][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_587;WeightsStore[1][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_588;WeightsStore[1][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_589;WeightsStore[1][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_590;WeightsStore[1][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_591;WeightsStore[1][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_592;WeightsStore[1][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_593;WeightsStore[1][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_594;WeightsStore[1][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_595;WeightsStore[1][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_596;WeightsStore[1][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_597;WeightsStore[1][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_598;WeightsStore[1][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_599;WeightsStore[1][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_600;WeightsStore[1][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_601;WeightsStore[1][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_602;WeightsStore[1][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_603;WeightsStore[1][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_604;WeightsStore[1][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_605;WeightsStore[1][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_606;WeightsStore[1][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_607;WeightsStore[1][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_608;WeightsStore[1][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_609;WeightsStore[1][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_610;WeightsStore[1][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_611;WeightsStore[1][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_612;WeightsStore[1][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_613;WeightsStore[1][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_614;WeightsStore[1][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_615;WeightsStore[1][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_616;WeightsStore[1][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_617;WeightsStore[1][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_618;WeightsStore[1][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_619;WeightsStore[1][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_620;WeightsStore[1][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_621;WeightsStore[1][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_622;WeightsStore[1][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_623;WeightsStore[1][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_624;WeightsStore[1][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_625;WeightsStore[1][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_626;WeightsStore[1][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_627;WeightsStore[1][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_628;WeightsStore[1][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_629;WeightsStore[1][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_630;WeightsStore[1][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_631;WeightsStore[1][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_632;WeightsStore[1][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_633;WeightsStore[1][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_634;WeightsStore[1][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_635;WeightsStore[1][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_636;WeightsStore[1][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_637;WeightsStore[1][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_638;WeightsStore[1][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_639;WeightsStore[1][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_640;WeightsStore[1][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_641;WeightsStore[1][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_642;WeightsStore[1][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_643;WeightsStore[1][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_644;WeightsStore[1][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_645;WeightsStore[1][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_646;WeightsStore[1][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_647;WeightsStore[1][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_648;WeightsStore[1][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_649;WeightsStore[1][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_650;WeightsStore[1][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_651;WeightsStore[1][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_652;WeightsStore[1][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_653;WeightsStore[1][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_654;WeightsStore[1][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_655;WeightsStore[1][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_656;WeightsStore[1][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_657;WeightsStore[1][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_658;WeightsStore[1][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_659;WeightsStore[1][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_660;WeightsStore[1][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_661;WeightsStore[1][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_662;WeightsStore[1][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_663;WeightsStore[1][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_664;WeightsStore[1][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_665;WeightsStore[1][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_666;WeightsStore[1][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_667;WeightsStore[1][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_668;WeightsStore[1][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_669;WeightsStore[1][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_670;WeightsStore[1][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_671;WeightsStore[1][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_672;WeightsStore[1][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_673;WeightsStore[1][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_674;WeightsStore[1][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_675;WeightsStore[1][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_676;WeightsStore[1][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_677;WeightsStore[1][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_678;WeightsStore[1][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_679;WeightsStore[1][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_680;WeightsStore[1][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_681;WeightsStore[1][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_682;WeightsStore[1][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_683;WeightsStore[1][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_684;WeightsStore[1][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_685;WeightsStore[1][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_686;WeightsStore[1][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_687;WeightsStore[1][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_688;WeightsStore[1][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_689;WeightsStore[1][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_690;WeightsStore[1][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_691;WeightsStore[1][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_692;WeightsStore[1][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_693;WeightsStore[1][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_694;WeightsStore[1][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_695;WeightsStore[1][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_696;WeightsStore[1][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_697;WeightsStore[1][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_698;WeightsStore[1][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_699;WeightsStore[1][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_700;WeightsStore[1][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_701;WeightsStore[1][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_702;WeightsStore[1][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_703;WeightsStore[1][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_704;WeightsStore[1][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_705;WeightsStore[1][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_706;WeightsStore[1][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_707;WeightsStore[1][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_708;WeightsStore[1][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_709;WeightsStore[1][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_710;WeightsStore[1][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_711;WeightsStore[1][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_712;WeightsStore[1][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_713;WeightsStore[1][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_714;WeightsStore[1][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_715;WeightsStore[1][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_716;WeightsStore[1][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_717;WeightsStore[1][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_718;WeightsStore[1][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_719;WeightsStore[1][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_720;WeightsStore[1][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_721;WeightsStore[1][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_722;WeightsStore[1][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_723;WeightsStore[1][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_724;WeightsStore[1][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_725;WeightsStore[1][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_726;WeightsStore[1][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_727;WeightsStore[1][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_728;WeightsStore[1][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_729;WeightsStore[1][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_730;WeightsStore[1][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_731;WeightsStore[1][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_732;WeightsStore[1][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_733;WeightsStore[1][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_734;WeightsStore[1][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_735;WeightsStore[1][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_736;WeightsStore[1][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_737;WeightsStore[1][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_738;WeightsStore[1][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_739;WeightsStore[1][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_740;WeightsStore[1][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_741;WeightsStore[1][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_742;WeightsStore[1][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_743;WeightsStore[1][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_744;WeightsStore[1][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_745;WeightsStore[1][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_746;WeightsStore[1][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_747;WeightsStore[1][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_748;WeightsStore[1][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_749;WeightsStore[1][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_750;WeightsStore[1][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_751;WeightsStore[1][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_752;WeightsStore[1][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_753;WeightsStore[1][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_754;WeightsStore[1][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_755;WeightsStore[1][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_756;WeightsStore[1][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_757;WeightsStore[1][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_758;WeightsStore[1][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_759;WeightsStore[1][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_760;WeightsStore[1][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_761;WeightsStore[1][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_762;WeightsStore[1][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_763;WeightsStore[1][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_764;WeightsStore[1][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_765;WeightsStore[1][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_766;WeightsStore[1][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_767;WeightsStore[1][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_768;WeightsStore[1][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_769;WeightsStore[1][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_770;WeightsStore[1][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_771;WeightsStore[1][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_772;WeightsStore[1][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_773;WeightsStore[1][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_774;WeightsStore[1][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_775;WeightsStore[1][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_776;WeightsStore[1][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_777;WeightsStore[1][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_778;WeightsStore[1][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_779;WeightsStore[1][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_780;WeightsStore[1][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_781;WeightsStore[1][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_782;WeightsStore[1][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_783;WeightsStore[1][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_1_784;WeightsStore[2][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_0;WeightsStore[2][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_1;WeightsStore[2][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_2;WeightsStore[2][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_3;WeightsStore[2][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_4;WeightsStore[2][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_5;WeightsStore[2][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_6;WeightsStore[2][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_7;WeightsStore[2][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_8;WeightsStore[2][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_9;WeightsStore[2][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_10;WeightsStore[2][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_11;WeightsStore[2][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_12;WeightsStore[2][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_13;WeightsStore[2][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_14;WeightsStore[2][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_15;WeightsStore[2][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_16;WeightsStore[2][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_17;WeightsStore[2][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_18;WeightsStore[2][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_19;WeightsStore[2][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_20;WeightsStore[2][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_21;WeightsStore[2][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_22;WeightsStore[2][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_23;WeightsStore[2][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_24;WeightsStore[2][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_25;WeightsStore[2][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_26;WeightsStore[2][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_27;WeightsStore[2][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_28;WeightsStore[2][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_29;WeightsStore[2][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_30;WeightsStore[2][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_31;WeightsStore[2][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_32;WeightsStore[2][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_33;WeightsStore[2][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_34;WeightsStore[2][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_35;WeightsStore[2][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_36;WeightsStore[2][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_37;WeightsStore[2][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_38;WeightsStore[2][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_39;WeightsStore[2][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_40;WeightsStore[2][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_41;WeightsStore[2][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_42;WeightsStore[2][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_43;WeightsStore[2][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_44;WeightsStore[2][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_45;WeightsStore[2][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_46;WeightsStore[2][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_47;WeightsStore[2][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_48;WeightsStore[2][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_49;WeightsStore[2][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_50;WeightsStore[2][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_51;WeightsStore[2][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_52;WeightsStore[2][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_53;WeightsStore[2][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_54;WeightsStore[2][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_55;WeightsStore[2][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_56;WeightsStore[2][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_57;WeightsStore[2][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_58;WeightsStore[2][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_59;WeightsStore[2][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_60;WeightsStore[2][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_61;WeightsStore[2][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_62;WeightsStore[2][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_63;WeightsStore[2][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_64;WeightsStore[2][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_65;WeightsStore[2][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_66;WeightsStore[2][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_67;WeightsStore[2][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_68;WeightsStore[2][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_69;WeightsStore[2][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_70;WeightsStore[2][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_71;WeightsStore[2][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_72;WeightsStore[2][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_73;WeightsStore[2][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_74;WeightsStore[2][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_75;WeightsStore[2][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_76;WeightsStore[2][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_77;WeightsStore[2][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_78;WeightsStore[2][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_79;WeightsStore[2][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_80;WeightsStore[2][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_81;WeightsStore[2][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_82;WeightsStore[2][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_83;WeightsStore[2][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_84;WeightsStore[2][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_85;WeightsStore[2][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_86;WeightsStore[2][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_87;WeightsStore[2][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_88;WeightsStore[2][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_89;WeightsStore[2][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_90;WeightsStore[2][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_91;WeightsStore[2][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_92;WeightsStore[2][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_93;WeightsStore[2][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_94;WeightsStore[2][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_95;WeightsStore[2][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_96;WeightsStore[2][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_97;WeightsStore[2][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_98;WeightsStore[2][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_99;WeightsStore[2][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_100;WeightsStore[2][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_101;WeightsStore[2][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_102;WeightsStore[2][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_103;WeightsStore[2][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_104;WeightsStore[2][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_105;WeightsStore[2][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_106;WeightsStore[2][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_107;WeightsStore[2][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_108;WeightsStore[2][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_109;WeightsStore[2][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_110;WeightsStore[2][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_111;WeightsStore[2][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_112;WeightsStore[2][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_113;WeightsStore[2][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_114;WeightsStore[2][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_115;WeightsStore[2][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_116;WeightsStore[2][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_117;WeightsStore[2][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_118;WeightsStore[2][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_119;WeightsStore[2][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_120;WeightsStore[2][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_121;WeightsStore[2][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_122;WeightsStore[2][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_123;WeightsStore[2][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_124;WeightsStore[2][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_125;WeightsStore[2][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_126;WeightsStore[2][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_127;WeightsStore[2][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_128;WeightsStore[2][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_129;WeightsStore[2][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_130;WeightsStore[2][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_131;WeightsStore[2][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_132;WeightsStore[2][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_133;WeightsStore[2][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_134;WeightsStore[2][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_135;WeightsStore[2][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_136;WeightsStore[2][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_137;WeightsStore[2][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_138;WeightsStore[2][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_139;WeightsStore[2][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_140;WeightsStore[2][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_141;WeightsStore[2][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_142;WeightsStore[2][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_143;WeightsStore[2][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_144;WeightsStore[2][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_145;WeightsStore[2][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_146;WeightsStore[2][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_147;WeightsStore[2][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_148;WeightsStore[2][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_149;WeightsStore[2][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_150;WeightsStore[2][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_151;WeightsStore[2][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_152;WeightsStore[2][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_153;WeightsStore[2][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_154;WeightsStore[2][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_155;WeightsStore[2][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_156;WeightsStore[2][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_157;WeightsStore[2][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_158;WeightsStore[2][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_159;WeightsStore[2][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_160;WeightsStore[2][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_161;WeightsStore[2][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_162;WeightsStore[2][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_163;WeightsStore[2][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_164;WeightsStore[2][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_165;WeightsStore[2][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_166;WeightsStore[2][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_167;WeightsStore[2][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_168;WeightsStore[2][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_169;WeightsStore[2][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_170;WeightsStore[2][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_171;WeightsStore[2][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_172;WeightsStore[2][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_173;WeightsStore[2][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_174;WeightsStore[2][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_175;WeightsStore[2][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_176;WeightsStore[2][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_177;WeightsStore[2][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_178;WeightsStore[2][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_179;WeightsStore[2][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_180;WeightsStore[2][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_181;WeightsStore[2][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_182;WeightsStore[2][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_183;WeightsStore[2][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_184;WeightsStore[2][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_185;WeightsStore[2][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_186;WeightsStore[2][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_187;WeightsStore[2][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_188;WeightsStore[2][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_189;WeightsStore[2][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_190;WeightsStore[2][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_191;WeightsStore[2][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_192;WeightsStore[2][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_193;WeightsStore[2][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_194;WeightsStore[2][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_195;WeightsStore[2][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_196;WeightsStore[2][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_197;WeightsStore[2][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_198;WeightsStore[2][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_199;WeightsStore[2][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_200;WeightsStore[2][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_201;WeightsStore[2][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_202;WeightsStore[2][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_203;WeightsStore[2][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_204;WeightsStore[2][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_205;WeightsStore[2][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_206;WeightsStore[2][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_207;WeightsStore[2][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_208;WeightsStore[2][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_209;WeightsStore[2][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_210;WeightsStore[2][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_211;WeightsStore[2][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_212;WeightsStore[2][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_213;WeightsStore[2][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_214;WeightsStore[2][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_215;WeightsStore[2][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_216;WeightsStore[2][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_217;WeightsStore[2][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_218;WeightsStore[2][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_219;WeightsStore[2][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_220;WeightsStore[2][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_221;WeightsStore[2][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_222;WeightsStore[2][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_223;WeightsStore[2][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_224;WeightsStore[2][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_225;WeightsStore[2][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_226;WeightsStore[2][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_227;WeightsStore[2][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_228;WeightsStore[2][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_229;WeightsStore[2][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_230;WeightsStore[2][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_231;WeightsStore[2][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_232;WeightsStore[2][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_233;WeightsStore[2][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_234;WeightsStore[2][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_235;WeightsStore[2][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_236;WeightsStore[2][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_237;WeightsStore[2][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_238;WeightsStore[2][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_239;WeightsStore[2][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_240;WeightsStore[2][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_241;WeightsStore[2][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_242;WeightsStore[2][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_243;WeightsStore[2][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_244;WeightsStore[2][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_245;WeightsStore[2][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_246;WeightsStore[2][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_247;WeightsStore[2][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_248;WeightsStore[2][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_249;WeightsStore[2][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_250;WeightsStore[2][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_251;WeightsStore[2][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_252;WeightsStore[2][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_253;WeightsStore[2][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_254;WeightsStore[2][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_255;WeightsStore[2][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_256;WeightsStore[2][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_257;WeightsStore[2][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_258;WeightsStore[2][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_259;WeightsStore[2][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_260;WeightsStore[2][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_261;WeightsStore[2][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_262;WeightsStore[2][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_263;WeightsStore[2][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_264;WeightsStore[2][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_265;WeightsStore[2][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_266;WeightsStore[2][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_267;WeightsStore[2][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_268;WeightsStore[2][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_269;WeightsStore[2][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_270;WeightsStore[2][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_271;WeightsStore[2][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_272;WeightsStore[2][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_273;WeightsStore[2][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_274;WeightsStore[2][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_275;WeightsStore[2][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_276;WeightsStore[2][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_277;WeightsStore[2][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_278;WeightsStore[2][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_279;WeightsStore[2][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_280;WeightsStore[2][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_281;WeightsStore[2][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_282;WeightsStore[2][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_283;WeightsStore[2][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_284;WeightsStore[2][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_285;WeightsStore[2][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_286;WeightsStore[2][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_287;WeightsStore[2][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_288;WeightsStore[2][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_289;WeightsStore[2][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_290;WeightsStore[2][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_291;WeightsStore[2][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_292;WeightsStore[2][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_293;WeightsStore[2][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_294;WeightsStore[2][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_295;WeightsStore[2][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_296;WeightsStore[2][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_297;WeightsStore[2][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_298;WeightsStore[2][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_299;WeightsStore[2][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_300;WeightsStore[2][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_301;WeightsStore[2][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_302;WeightsStore[2][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_303;WeightsStore[2][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_304;WeightsStore[2][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_305;WeightsStore[2][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_306;WeightsStore[2][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_307;WeightsStore[2][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_308;WeightsStore[2][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_309;WeightsStore[2][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_310;WeightsStore[2][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_311;WeightsStore[2][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_312;WeightsStore[2][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_313;WeightsStore[2][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_314;WeightsStore[2][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_315;WeightsStore[2][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_316;WeightsStore[2][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_317;WeightsStore[2][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_318;WeightsStore[2][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_319;WeightsStore[2][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_320;WeightsStore[2][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_321;WeightsStore[2][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_322;WeightsStore[2][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_323;WeightsStore[2][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_324;WeightsStore[2][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_325;WeightsStore[2][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_326;WeightsStore[2][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_327;WeightsStore[2][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_328;WeightsStore[2][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_329;WeightsStore[2][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_330;WeightsStore[2][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_331;WeightsStore[2][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_332;WeightsStore[2][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_333;WeightsStore[2][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_334;WeightsStore[2][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_335;WeightsStore[2][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_336;WeightsStore[2][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_337;WeightsStore[2][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_338;WeightsStore[2][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_339;WeightsStore[2][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_340;WeightsStore[2][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_341;WeightsStore[2][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_342;WeightsStore[2][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_343;WeightsStore[2][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_344;WeightsStore[2][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_345;WeightsStore[2][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_346;WeightsStore[2][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_347;WeightsStore[2][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_348;WeightsStore[2][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_349;WeightsStore[2][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_350;WeightsStore[2][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_351;WeightsStore[2][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_352;WeightsStore[2][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_353;WeightsStore[2][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_354;WeightsStore[2][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_355;WeightsStore[2][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_356;WeightsStore[2][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_357;WeightsStore[2][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_358;WeightsStore[2][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_359;WeightsStore[2][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_360;WeightsStore[2][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_361;WeightsStore[2][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_362;WeightsStore[2][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_363;WeightsStore[2][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_364;WeightsStore[2][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_365;WeightsStore[2][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_366;WeightsStore[2][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_367;WeightsStore[2][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_368;WeightsStore[2][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_369;WeightsStore[2][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_370;WeightsStore[2][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_371;WeightsStore[2][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_372;WeightsStore[2][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_373;WeightsStore[2][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_374;WeightsStore[2][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_375;WeightsStore[2][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_376;WeightsStore[2][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_377;WeightsStore[2][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_378;WeightsStore[2][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_379;WeightsStore[2][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_380;WeightsStore[2][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_381;WeightsStore[2][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_382;WeightsStore[2][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_383;WeightsStore[2][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_384;WeightsStore[2][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_385;WeightsStore[2][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_386;WeightsStore[2][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_387;WeightsStore[2][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_388;WeightsStore[2][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_389;WeightsStore[2][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_390;WeightsStore[2][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_391;WeightsStore[2][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_392;WeightsStore[2][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_393;WeightsStore[2][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_394;WeightsStore[2][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_395;WeightsStore[2][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_396;WeightsStore[2][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_397;WeightsStore[2][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_398;WeightsStore[2][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_399;WeightsStore[2][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_400;WeightsStore[2][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_401;WeightsStore[2][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_402;WeightsStore[2][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_403;WeightsStore[2][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_404;WeightsStore[2][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_405;WeightsStore[2][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_406;WeightsStore[2][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_407;WeightsStore[2][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_408;WeightsStore[2][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_409;WeightsStore[2][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_410;WeightsStore[2][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_411;WeightsStore[2][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_412;WeightsStore[2][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_413;WeightsStore[2][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_414;WeightsStore[2][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_415;WeightsStore[2][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_416;WeightsStore[2][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_417;WeightsStore[2][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_418;WeightsStore[2][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_419;WeightsStore[2][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_420;WeightsStore[2][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_421;WeightsStore[2][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_422;WeightsStore[2][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_423;WeightsStore[2][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_424;WeightsStore[2][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_425;WeightsStore[2][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_426;WeightsStore[2][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_427;WeightsStore[2][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_428;WeightsStore[2][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_429;WeightsStore[2][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_430;WeightsStore[2][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_431;WeightsStore[2][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_432;WeightsStore[2][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_433;WeightsStore[2][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_434;WeightsStore[2][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_435;WeightsStore[2][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_436;WeightsStore[2][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_437;WeightsStore[2][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_438;WeightsStore[2][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_439;WeightsStore[2][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_440;WeightsStore[2][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_441;WeightsStore[2][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_442;WeightsStore[2][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_443;WeightsStore[2][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_444;WeightsStore[2][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_445;WeightsStore[2][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_446;WeightsStore[2][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_447;WeightsStore[2][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_448;WeightsStore[2][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_449;WeightsStore[2][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_450;WeightsStore[2][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_451;WeightsStore[2][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_452;WeightsStore[2][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_453;WeightsStore[2][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_454;WeightsStore[2][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_455;WeightsStore[2][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_456;WeightsStore[2][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_457;WeightsStore[2][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_458;WeightsStore[2][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_459;WeightsStore[2][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_460;WeightsStore[2][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_461;WeightsStore[2][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_462;WeightsStore[2][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_463;WeightsStore[2][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_464;WeightsStore[2][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_465;WeightsStore[2][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_466;WeightsStore[2][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_467;WeightsStore[2][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_468;WeightsStore[2][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_469;WeightsStore[2][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_470;WeightsStore[2][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_471;WeightsStore[2][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_472;WeightsStore[2][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_473;WeightsStore[2][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_474;WeightsStore[2][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_475;WeightsStore[2][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_476;WeightsStore[2][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_477;WeightsStore[2][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_478;WeightsStore[2][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_479;WeightsStore[2][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_480;WeightsStore[2][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_481;WeightsStore[2][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_482;WeightsStore[2][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_483;WeightsStore[2][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_484;WeightsStore[2][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_485;WeightsStore[2][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_486;WeightsStore[2][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_487;WeightsStore[2][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_488;WeightsStore[2][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_489;WeightsStore[2][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_490;WeightsStore[2][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_491;WeightsStore[2][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_492;WeightsStore[2][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_493;WeightsStore[2][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_494;WeightsStore[2][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_495;WeightsStore[2][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_496;WeightsStore[2][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_497;WeightsStore[2][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_498;WeightsStore[2][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_499;WeightsStore[2][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_500;WeightsStore[2][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_501;WeightsStore[2][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_502;WeightsStore[2][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_503;WeightsStore[2][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_504;WeightsStore[2][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_505;WeightsStore[2][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_506;WeightsStore[2][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_507;WeightsStore[2][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_508;WeightsStore[2][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_509;WeightsStore[2][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_510;WeightsStore[2][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_511;WeightsStore[2][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_512;WeightsStore[2][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_513;WeightsStore[2][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_514;WeightsStore[2][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_515;WeightsStore[2][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_516;WeightsStore[2][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_517;WeightsStore[2][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_518;WeightsStore[2][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_519;WeightsStore[2][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_520;WeightsStore[2][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_521;WeightsStore[2][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_522;WeightsStore[2][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_523;WeightsStore[2][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_524;WeightsStore[2][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_525;WeightsStore[2][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_526;WeightsStore[2][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_527;WeightsStore[2][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_528;WeightsStore[2][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_529;WeightsStore[2][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_530;WeightsStore[2][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_531;WeightsStore[2][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_532;WeightsStore[2][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_533;WeightsStore[2][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_534;WeightsStore[2][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_535;WeightsStore[2][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_536;WeightsStore[2][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_537;WeightsStore[2][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_538;WeightsStore[2][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_539;WeightsStore[2][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_540;WeightsStore[2][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_541;WeightsStore[2][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_542;WeightsStore[2][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_543;WeightsStore[2][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_544;WeightsStore[2][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_545;WeightsStore[2][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_546;WeightsStore[2][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_547;WeightsStore[2][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_548;WeightsStore[2][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_549;WeightsStore[2][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_550;WeightsStore[2][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_551;WeightsStore[2][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_552;WeightsStore[2][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_553;WeightsStore[2][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_554;WeightsStore[2][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_555;WeightsStore[2][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_556;WeightsStore[2][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_557;WeightsStore[2][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_558;WeightsStore[2][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_559;WeightsStore[2][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_560;WeightsStore[2][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_561;WeightsStore[2][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_562;WeightsStore[2][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_563;WeightsStore[2][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_564;WeightsStore[2][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_565;WeightsStore[2][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_566;WeightsStore[2][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_567;WeightsStore[2][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_568;WeightsStore[2][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_569;WeightsStore[2][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_570;WeightsStore[2][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_571;WeightsStore[2][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_572;WeightsStore[2][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_573;WeightsStore[2][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_574;WeightsStore[2][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_575;WeightsStore[2][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_576;WeightsStore[2][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_577;WeightsStore[2][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_578;WeightsStore[2][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_579;WeightsStore[2][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_580;WeightsStore[2][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_581;WeightsStore[2][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_582;WeightsStore[2][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_583;WeightsStore[2][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_584;WeightsStore[2][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_585;WeightsStore[2][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_586;WeightsStore[2][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_587;WeightsStore[2][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_588;WeightsStore[2][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_589;WeightsStore[2][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_590;WeightsStore[2][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_591;WeightsStore[2][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_592;WeightsStore[2][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_593;WeightsStore[2][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_594;WeightsStore[2][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_595;WeightsStore[2][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_596;WeightsStore[2][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_597;WeightsStore[2][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_598;WeightsStore[2][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_599;WeightsStore[2][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_600;WeightsStore[2][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_601;WeightsStore[2][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_602;WeightsStore[2][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_603;WeightsStore[2][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_604;WeightsStore[2][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_605;WeightsStore[2][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_606;WeightsStore[2][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_607;WeightsStore[2][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_608;WeightsStore[2][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_609;WeightsStore[2][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_610;WeightsStore[2][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_611;WeightsStore[2][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_612;WeightsStore[2][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_613;WeightsStore[2][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_614;WeightsStore[2][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_615;WeightsStore[2][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_616;WeightsStore[2][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_617;WeightsStore[2][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_618;WeightsStore[2][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_619;WeightsStore[2][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_620;WeightsStore[2][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_621;WeightsStore[2][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_622;WeightsStore[2][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_623;WeightsStore[2][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_624;WeightsStore[2][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_625;WeightsStore[2][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_626;WeightsStore[2][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_627;WeightsStore[2][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_628;WeightsStore[2][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_629;WeightsStore[2][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_630;WeightsStore[2][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_631;WeightsStore[2][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_632;WeightsStore[2][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_633;WeightsStore[2][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_634;WeightsStore[2][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_635;WeightsStore[2][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_636;WeightsStore[2][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_637;WeightsStore[2][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_638;WeightsStore[2][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_639;WeightsStore[2][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_640;WeightsStore[2][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_641;WeightsStore[2][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_642;WeightsStore[2][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_643;WeightsStore[2][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_644;WeightsStore[2][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_645;WeightsStore[2][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_646;WeightsStore[2][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_647;WeightsStore[2][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_648;WeightsStore[2][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_649;WeightsStore[2][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_650;WeightsStore[2][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_651;WeightsStore[2][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_652;WeightsStore[2][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_653;WeightsStore[2][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_654;WeightsStore[2][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_655;WeightsStore[2][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_656;WeightsStore[2][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_657;WeightsStore[2][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_658;WeightsStore[2][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_659;WeightsStore[2][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_660;WeightsStore[2][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_661;WeightsStore[2][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_662;WeightsStore[2][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_663;WeightsStore[2][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_664;WeightsStore[2][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_665;WeightsStore[2][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_666;WeightsStore[2][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_667;WeightsStore[2][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_668;WeightsStore[2][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_669;WeightsStore[2][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_670;WeightsStore[2][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_671;WeightsStore[2][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_672;WeightsStore[2][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_673;WeightsStore[2][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_674;WeightsStore[2][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_675;WeightsStore[2][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_676;WeightsStore[2][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_677;WeightsStore[2][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_678;WeightsStore[2][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_679;WeightsStore[2][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_680;WeightsStore[2][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_681;WeightsStore[2][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_682;WeightsStore[2][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_683;WeightsStore[2][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_684;WeightsStore[2][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_685;WeightsStore[2][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_686;WeightsStore[2][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_687;WeightsStore[2][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_688;WeightsStore[2][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_689;WeightsStore[2][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_690;WeightsStore[2][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_691;WeightsStore[2][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_692;WeightsStore[2][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_693;WeightsStore[2][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_694;WeightsStore[2][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_695;WeightsStore[2][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_696;WeightsStore[2][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_697;WeightsStore[2][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_698;WeightsStore[2][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_699;WeightsStore[2][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_700;WeightsStore[2][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_701;WeightsStore[2][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_702;WeightsStore[2][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_703;WeightsStore[2][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_704;WeightsStore[2][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_705;WeightsStore[2][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_706;WeightsStore[2][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_707;WeightsStore[2][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_708;WeightsStore[2][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_709;WeightsStore[2][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_710;WeightsStore[2][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_711;WeightsStore[2][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_712;WeightsStore[2][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_713;WeightsStore[2][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_714;WeightsStore[2][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_715;WeightsStore[2][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_716;WeightsStore[2][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_717;WeightsStore[2][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_718;WeightsStore[2][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_719;WeightsStore[2][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_720;WeightsStore[2][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_721;WeightsStore[2][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_722;WeightsStore[2][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_723;WeightsStore[2][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_724;WeightsStore[2][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_725;WeightsStore[2][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_726;WeightsStore[2][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_727;WeightsStore[2][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_728;WeightsStore[2][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_729;WeightsStore[2][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_730;WeightsStore[2][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_731;WeightsStore[2][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_732;WeightsStore[2][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_733;WeightsStore[2][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_734;WeightsStore[2][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_735;WeightsStore[2][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_736;WeightsStore[2][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_737;WeightsStore[2][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_738;WeightsStore[2][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_739;WeightsStore[2][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_740;WeightsStore[2][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_741;WeightsStore[2][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_742;WeightsStore[2][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_743;WeightsStore[2][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_744;WeightsStore[2][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_745;WeightsStore[2][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_746;WeightsStore[2][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_747;WeightsStore[2][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_748;WeightsStore[2][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_749;WeightsStore[2][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_750;WeightsStore[2][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_751;WeightsStore[2][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_752;WeightsStore[2][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_753;WeightsStore[2][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_754;WeightsStore[2][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_755;WeightsStore[2][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_756;WeightsStore[2][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_757;WeightsStore[2][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_758;WeightsStore[2][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_759;WeightsStore[2][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_760;WeightsStore[2][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_761;WeightsStore[2][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_762;WeightsStore[2][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_763;WeightsStore[2][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_764;WeightsStore[2][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_765;WeightsStore[2][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_766;WeightsStore[2][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_767;WeightsStore[2][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_768;WeightsStore[2][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_769;WeightsStore[2][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_770;WeightsStore[2][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_771;WeightsStore[2][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_772;WeightsStore[2][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_773;WeightsStore[2][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_774;WeightsStore[2][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_775;WeightsStore[2][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_776;WeightsStore[2][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_777;WeightsStore[2][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_778;WeightsStore[2][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_779;WeightsStore[2][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_780;WeightsStore[2][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_781;WeightsStore[2][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_782;WeightsStore[2][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_783;WeightsStore[2][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_2_784;WeightsStore[3][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_0;WeightsStore[3][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_1;WeightsStore[3][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_2;WeightsStore[3][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_3;WeightsStore[3][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_4;WeightsStore[3][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_5;WeightsStore[3][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_6;WeightsStore[3][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_7;WeightsStore[3][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_8;WeightsStore[3][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_9;WeightsStore[3][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_10;WeightsStore[3][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_11;WeightsStore[3][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_12;WeightsStore[3][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_13;WeightsStore[3][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_14;WeightsStore[3][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_15;WeightsStore[3][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_16;WeightsStore[3][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_17;WeightsStore[3][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_18;WeightsStore[3][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_19;WeightsStore[3][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_20;WeightsStore[3][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_21;WeightsStore[3][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_22;WeightsStore[3][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_23;WeightsStore[3][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_24;WeightsStore[3][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_25;WeightsStore[3][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_26;WeightsStore[3][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_27;WeightsStore[3][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_28;WeightsStore[3][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_29;WeightsStore[3][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_30;WeightsStore[3][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_31;WeightsStore[3][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_32;WeightsStore[3][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_33;WeightsStore[3][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_34;WeightsStore[3][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_35;WeightsStore[3][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_36;WeightsStore[3][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_37;WeightsStore[3][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_38;WeightsStore[3][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_39;WeightsStore[3][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_40;WeightsStore[3][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_41;WeightsStore[3][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_42;WeightsStore[3][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_43;WeightsStore[3][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_44;WeightsStore[3][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_45;WeightsStore[3][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_46;WeightsStore[3][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_47;WeightsStore[3][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_48;WeightsStore[3][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_49;WeightsStore[3][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_50;WeightsStore[3][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_51;WeightsStore[3][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_52;WeightsStore[3][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_53;WeightsStore[3][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_54;WeightsStore[3][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_55;WeightsStore[3][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_56;WeightsStore[3][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_57;WeightsStore[3][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_58;WeightsStore[3][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_59;WeightsStore[3][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_60;WeightsStore[3][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_61;WeightsStore[3][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_62;WeightsStore[3][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_63;WeightsStore[3][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_64;WeightsStore[3][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_65;WeightsStore[3][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_66;WeightsStore[3][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_67;WeightsStore[3][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_68;WeightsStore[3][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_69;WeightsStore[3][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_70;WeightsStore[3][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_71;WeightsStore[3][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_72;WeightsStore[3][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_73;WeightsStore[3][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_74;WeightsStore[3][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_75;WeightsStore[3][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_76;WeightsStore[3][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_77;WeightsStore[3][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_78;WeightsStore[3][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_79;WeightsStore[3][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_80;WeightsStore[3][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_81;WeightsStore[3][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_82;WeightsStore[3][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_83;WeightsStore[3][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_84;WeightsStore[3][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_85;WeightsStore[3][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_86;WeightsStore[3][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_87;WeightsStore[3][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_88;WeightsStore[3][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_89;WeightsStore[3][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_90;WeightsStore[3][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_91;WeightsStore[3][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_92;WeightsStore[3][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_93;WeightsStore[3][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_94;WeightsStore[3][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_95;WeightsStore[3][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_96;WeightsStore[3][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_97;WeightsStore[3][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_98;WeightsStore[3][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_99;WeightsStore[3][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_100;WeightsStore[3][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_101;WeightsStore[3][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_102;WeightsStore[3][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_103;WeightsStore[3][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_104;WeightsStore[3][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_105;WeightsStore[3][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_106;WeightsStore[3][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_107;WeightsStore[3][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_108;WeightsStore[3][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_109;WeightsStore[3][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_110;WeightsStore[3][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_111;WeightsStore[3][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_112;WeightsStore[3][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_113;WeightsStore[3][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_114;WeightsStore[3][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_115;WeightsStore[3][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_116;WeightsStore[3][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_117;WeightsStore[3][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_118;WeightsStore[3][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_119;WeightsStore[3][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_120;WeightsStore[3][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_121;WeightsStore[3][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_122;WeightsStore[3][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_123;WeightsStore[3][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_124;WeightsStore[3][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_125;WeightsStore[3][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_126;WeightsStore[3][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_127;WeightsStore[3][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_128;WeightsStore[3][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_129;WeightsStore[3][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_130;WeightsStore[3][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_131;WeightsStore[3][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_132;WeightsStore[3][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_133;WeightsStore[3][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_134;WeightsStore[3][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_135;WeightsStore[3][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_136;WeightsStore[3][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_137;WeightsStore[3][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_138;WeightsStore[3][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_139;WeightsStore[3][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_140;WeightsStore[3][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_141;WeightsStore[3][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_142;WeightsStore[3][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_143;WeightsStore[3][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_144;WeightsStore[3][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_145;WeightsStore[3][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_146;WeightsStore[3][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_147;WeightsStore[3][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_148;WeightsStore[3][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_149;WeightsStore[3][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_150;WeightsStore[3][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_151;WeightsStore[3][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_152;WeightsStore[3][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_153;WeightsStore[3][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_154;WeightsStore[3][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_155;WeightsStore[3][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_156;WeightsStore[3][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_157;WeightsStore[3][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_158;WeightsStore[3][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_159;WeightsStore[3][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_160;WeightsStore[3][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_161;WeightsStore[3][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_162;WeightsStore[3][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_163;WeightsStore[3][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_164;WeightsStore[3][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_165;WeightsStore[3][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_166;WeightsStore[3][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_167;WeightsStore[3][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_168;WeightsStore[3][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_169;WeightsStore[3][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_170;WeightsStore[3][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_171;WeightsStore[3][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_172;WeightsStore[3][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_173;WeightsStore[3][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_174;WeightsStore[3][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_175;WeightsStore[3][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_176;WeightsStore[3][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_177;WeightsStore[3][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_178;WeightsStore[3][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_179;WeightsStore[3][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_180;WeightsStore[3][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_181;WeightsStore[3][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_182;WeightsStore[3][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_183;WeightsStore[3][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_184;WeightsStore[3][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_185;WeightsStore[3][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_186;WeightsStore[3][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_187;WeightsStore[3][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_188;WeightsStore[3][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_189;WeightsStore[3][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_190;WeightsStore[3][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_191;WeightsStore[3][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_192;WeightsStore[3][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_193;WeightsStore[3][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_194;WeightsStore[3][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_195;WeightsStore[3][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_196;WeightsStore[3][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_197;WeightsStore[3][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_198;WeightsStore[3][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_199;WeightsStore[3][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_200;WeightsStore[3][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_201;WeightsStore[3][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_202;WeightsStore[3][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_203;WeightsStore[3][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_204;WeightsStore[3][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_205;WeightsStore[3][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_206;WeightsStore[3][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_207;WeightsStore[3][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_208;WeightsStore[3][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_209;WeightsStore[3][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_210;WeightsStore[3][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_211;WeightsStore[3][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_212;WeightsStore[3][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_213;WeightsStore[3][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_214;WeightsStore[3][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_215;WeightsStore[3][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_216;WeightsStore[3][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_217;WeightsStore[3][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_218;WeightsStore[3][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_219;WeightsStore[3][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_220;WeightsStore[3][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_221;WeightsStore[3][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_222;WeightsStore[3][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_223;WeightsStore[3][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_224;WeightsStore[3][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_225;WeightsStore[3][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_226;WeightsStore[3][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_227;WeightsStore[3][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_228;WeightsStore[3][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_229;WeightsStore[3][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_230;WeightsStore[3][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_231;WeightsStore[3][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_232;WeightsStore[3][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_233;WeightsStore[3][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_234;WeightsStore[3][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_235;WeightsStore[3][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_236;WeightsStore[3][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_237;WeightsStore[3][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_238;WeightsStore[3][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_239;WeightsStore[3][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_240;WeightsStore[3][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_241;WeightsStore[3][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_242;WeightsStore[3][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_243;WeightsStore[3][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_244;WeightsStore[3][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_245;WeightsStore[3][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_246;WeightsStore[3][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_247;WeightsStore[3][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_248;WeightsStore[3][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_249;WeightsStore[3][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_250;WeightsStore[3][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_251;WeightsStore[3][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_252;WeightsStore[3][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_253;WeightsStore[3][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_254;WeightsStore[3][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_255;WeightsStore[3][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_256;WeightsStore[3][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_257;WeightsStore[3][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_258;WeightsStore[3][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_259;WeightsStore[3][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_260;WeightsStore[3][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_261;WeightsStore[3][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_262;WeightsStore[3][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_263;WeightsStore[3][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_264;WeightsStore[3][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_265;WeightsStore[3][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_266;WeightsStore[3][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_267;WeightsStore[3][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_268;WeightsStore[3][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_269;WeightsStore[3][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_270;WeightsStore[3][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_271;WeightsStore[3][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_272;WeightsStore[3][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_273;WeightsStore[3][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_274;WeightsStore[3][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_275;WeightsStore[3][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_276;WeightsStore[3][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_277;WeightsStore[3][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_278;WeightsStore[3][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_279;WeightsStore[3][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_280;WeightsStore[3][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_281;WeightsStore[3][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_282;WeightsStore[3][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_283;WeightsStore[3][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_284;WeightsStore[3][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_285;WeightsStore[3][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_286;WeightsStore[3][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_287;WeightsStore[3][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_288;WeightsStore[3][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_289;WeightsStore[3][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_290;WeightsStore[3][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_291;WeightsStore[3][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_292;WeightsStore[3][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_293;WeightsStore[3][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_294;WeightsStore[3][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_295;WeightsStore[3][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_296;WeightsStore[3][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_297;WeightsStore[3][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_298;WeightsStore[3][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_299;WeightsStore[3][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_300;WeightsStore[3][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_301;WeightsStore[3][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_302;WeightsStore[3][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_303;WeightsStore[3][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_304;WeightsStore[3][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_305;WeightsStore[3][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_306;WeightsStore[3][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_307;WeightsStore[3][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_308;WeightsStore[3][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_309;WeightsStore[3][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_310;WeightsStore[3][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_311;WeightsStore[3][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_312;WeightsStore[3][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_313;WeightsStore[3][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_314;WeightsStore[3][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_315;WeightsStore[3][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_316;WeightsStore[3][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_317;WeightsStore[3][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_318;WeightsStore[3][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_319;WeightsStore[3][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_320;WeightsStore[3][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_321;WeightsStore[3][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_322;WeightsStore[3][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_323;WeightsStore[3][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_324;WeightsStore[3][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_325;WeightsStore[3][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_326;WeightsStore[3][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_327;WeightsStore[3][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_328;WeightsStore[3][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_329;WeightsStore[3][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_330;WeightsStore[3][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_331;WeightsStore[3][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_332;WeightsStore[3][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_333;WeightsStore[3][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_334;WeightsStore[3][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_335;WeightsStore[3][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_336;WeightsStore[3][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_337;WeightsStore[3][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_338;WeightsStore[3][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_339;WeightsStore[3][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_340;WeightsStore[3][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_341;WeightsStore[3][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_342;WeightsStore[3][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_343;WeightsStore[3][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_344;WeightsStore[3][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_345;WeightsStore[3][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_346;WeightsStore[3][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_347;WeightsStore[3][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_348;WeightsStore[3][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_349;WeightsStore[3][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_350;WeightsStore[3][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_351;WeightsStore[3][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_352;WeightsStore[3][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_353;WeightsStore[3][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_354;WeightsStore[3][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_355;WeightsStore[3][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_356;WeightsStore[3][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_357;WeightsStore[3][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_358;WeightsStore[3][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_359;WeightsStore[3][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_360;WeightsStore[3][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_361;WeightsStore[3][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_362;WeightsStore[3][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_363;WeightsStore[3][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_364;WeightsStore[3][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_365;WeightsStore[3][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_366;WeightsStore[3][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_367;WeightsStore[3][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_368;WeightsStore[3][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_369;WeightsStore[3][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_370;WeightsStore[3][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_371;WeightsStore[3][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_372;WeightsStore[3][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_373;WeightsStore[3][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_374;WeightsStore[3][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_375;WeightsStore[3][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_376;WeightsStore[3][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_377;WeightsStore[3][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_378;WeightsStore[3][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_379;WeightsStore[3][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_380;WeightsStore[3][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_381;WeightsStore[3][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_382;WeightsStore[3][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_383;WeightsStore[3][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_384;WeightsStore[3][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_385;WeightsStore[3][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_386;WeightsStore[3][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_387;WeightsStore[3][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_388;WeightsStore[3][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_389;WeightsStore[3][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_390;WeightsStore[3][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_391;WeightsStore[3][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_392;WeightsStore[3][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_393;WeightsStore[3][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_394;WeightsStore[3][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_395;WeightsStore[3][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_396;WeightsStore[3][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_397;WeightsStore[3][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_398;WeightsStore[3][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_399;WeightsStore[3][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_400;WeightsStore[3][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_401;WeightsStore[3][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_402;WeightsStore[3][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_403;WeightsStore[3][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_404;WeightsStore[3][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_405;WeightsStore[3][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_406;WeightsStore[3][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_407;WeightsStore[3][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_408;WeightsStore[3][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_409;WeightsStore[3][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_410;WeightsStore[3][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_411;WeightsStore[3][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_412;WeightsStore[3][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_413;WeightsStore[3][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_414;WeightsStore[3][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_415;WeightsStore[3][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_416;WeightsStore[3][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_417;WeightsStore[3][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_418;WeightsStore[3][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_419;WeightsStore[3][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_420;WeightsStore[3][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_421;WeightsStore[3][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_422;WeightsStore[3][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_423;WeightsStore[3][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_424;WeightsStore[3][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_425;WeightsStore[3][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_426;WeightsStore[3][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_427;WeightsStore[3][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_428;WeightsStore[3][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_429;WeightsStore[3][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_430;WeightsStore[3][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_431;WeightsStore[3][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_432;WeightsStore[3][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_433;WeightsStore[3][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_434;WeightsStore[3][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_435;WeightsStore[3][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_436;WeightsStore[3][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_437;WeightsStore[3][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_438;WeightsStore[3][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_439;WeightsStore[3][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_440;WeightsStore[3][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_441;WeightsStore[3][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_442;WeightsStore[3][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_443;WeightsStore[3][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_444;WeightsStore[3][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_445;WeightsStore[3][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_446;WeightsStore[3][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_447;WeightsStore[3][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_448;WeightsStore[3][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_449;WeightsStore[3][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_450;WeightsStore[3][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_451;WeightsStore[3][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_452;WeightsStore[3][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_453;WeightsStore[3][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_454;WeightsStore[3][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_455;WeightsStore[3][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_456;WeightsStore[3][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_457;WeightsStore[3][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_458;WeightsStore[3][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_459;WeightsStore[3][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_460;WeightsStore[3][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_461;WeightsStore[3][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_462;WeightsStore[3][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_463;WeightsStore[3][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_464;WeightsStore[3][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_465;WeightsStore[3][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_466;WeightsStore[3][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_467;WeightsStore[3][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_468;WeightsStore[3][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_469;WeightsStore[3][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_470;WeightsStore[3][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_471;WeightsStore[3][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_472;WeightsStore[3][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_473;WeightsStore[3][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_474;WeightsStore[3][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_475;WeightsStore[3][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_476;WeightsStore[3][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_477;WeightsStore[3][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_478;WeightsStore[3][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_479;WeightsStore[3][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_480;WeightsStore[3][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_481;WeightsStore[3][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_482;WeightsStore[3][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_483;WeightsStore[3][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_484;WeightsStore[3][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_485;WeightsStore[3][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_486;WeightsStore[3][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_487;WeightsStore[3][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_488;WeightsStore[3][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_489;WeightsStore[3][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_490;WeightsStore[3][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_491;WeightsStore[3][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_492;WeightsStore[3][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_493;WeightsStore[3][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_494;WeightsStore[3][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_495;WeightsStore[3][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_496;WeightsStore[3][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_497;WeightsStore[3][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_498;WeightsStore[3][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_499;WeightsStore[3][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_500;WeightsStore[3][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_501;WeightsStore[3][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_502;WeightsStore[3][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_503;WeightsStore[3][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_504;WeightsStore[3][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_505;WeightsStore[3][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_506;WeightsStore[3][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_507;WeightsStore[3][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_508;WeightsStore[3][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_509;WeightsStore[3][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_510;WeightsStore[3][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_511;WeightsStore[3][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_512;WeightsStore[3][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_513;WeightsStore[3][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_514;WeightsStore[3][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_515;WeightsStore[3][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_516;WeightsStore[3][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_517;WeightsStore[3][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_518;WeightsStore[3][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_519;WeightsStore[3][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_520;WeightsStore[3][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_521;WeightsStore[3][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_522;WeightsStore[3][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_523;WeightsStore[3][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_524;WeightsStore[3][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_525;WeightsStore[3][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_526;WeightsStore[3][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_527;WeightsStore[3][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_528;WeightsStore[3][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_529;WeightsStore[3][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_530;WeightsStore[3][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_531;WeightsStore[3][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_532;WeightsStore[3][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_533;WeightsStore[3][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_534;WeightsStore[3][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_535;WeightsStore[3][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_536;WeightsStore[3][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_537;WeightsStore[3][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_538;WeightsStore[3][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_539;WeightsStore[3][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_540;WeightsStore[3][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_541;WeightsStore[3][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_542;WeightsStore[3][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_543;WeightsStore[3][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_544;WeightsStore[3][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_545;WeightsStore[3][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_546;WeightsStore[3][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_547;WeightsStore[3][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_548;WeightsStore[3][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_549;WeightsStore[3][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_550;WeightsStore[3][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_551;WeightsStore[3][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_552;WeightsStore[3][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_553;WeightsStore[3][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_554;WeightsStore[3][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_555;WeightsStore[3][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_556;WeightsStore[3][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_557;WeightsStore[3][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_558;WeightsStore[3][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_559;WeightsStore[3][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_560;WeightsStore[3][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_561;WeightsStore[3][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_562;WeightsStore[3][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_563;WeightsStore[3][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_564;WeightsStore[3][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_565;WeightsStore[3][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_566;WeightsStore[3][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_567;WeightsStore[3][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_568;WeightsStore[3][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_569;WeightsStore[3][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_570;WeightsStore[3][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_571;WeightsStore[3][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_572;WeightsStore[3][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_573;WeightsStore[3][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_574;WeightsStore[3][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_575;WeightsStore[3][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_576;WeightsStore[3][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_577;WeightsStore[3][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_578;WeightsStore[3][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_579;WeightsStore[3][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_580;WeightsStore[3][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_581;WeightsStore[3][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_582;WeightsStore[3][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_583;WeightsStore[3][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_584;WeightsStore[3][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_585;WeightsStore[3][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_586;WeightsStore[3][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_587;WeightsStore[3][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_588;WeightsStore[3][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_589;WeightsStore[3][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_590;WeightsStore[3][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_591;WeightsStore[3][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_592;WeightsStore[3][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_593;WeightsStore[3][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_594;WeightsStore[3][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_595;WeightsStore[3][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_596;WeightsStore[3][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_597;WeightsStore[3][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_598;WeightsStore[3][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_599;WeightsStore[3][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_600;WeightsStore[3][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_601;WeightsStore[3][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_602;WeightsStore[3][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_603;WeightsStore[3][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_604;WeightsStore[3][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_605;WeightsStore[3][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_606;WeightsStore[3][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_607;WeightsStore[3][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_608;WeightsStore[3][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_609;WeightsStore[3][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_610;WeightsStore[3][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_611;WeightsStore[3][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_612;WeightsStore[3][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_613;WeightsStore[3][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_614;WeightsStore[3][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_615;WeightsStore[3][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_616;WeightsStore[3][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_617;WeightsStore[3][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_618;WeightsStore[3][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_619;WeightsStore[3][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_620;WeightsStore[3][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_621;WeightsStore[3][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_622;WeightsStore[3][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_623;WeightsStore[3][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_624;WeightsStore[3][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_625;WeightsStore[3][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_626;WeightsStore[3][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_627;WeightsStore[3][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_628;WeightsStore[3][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_629;WeightsStore[3][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_630;WeightsStore[3][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_631;WeightsStore[3][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_632;WeightsStore[3][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_633;WeightsStore[3][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_634;WeightsStore[3][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_635;WeightsStore[3][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_636;WeightsStore[3][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_637;WeightsStore[3][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_638;WeightsStore[3][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_639;WeightsStore[3][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_640;WeightsStore[3][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_641;WeightsStore[3][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_642;WeightsStore[3][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_643;WeightsStore[3][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_644;WeightsStore[3][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_645;WeightsStore[3][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_646;WeightsStore[3][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_647;WeightsStore[3][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_648;WeightsStore[3][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_649;WeightsStore[3][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_650;WeightsStore[3][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_651;WeightsStore[3][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_652;WeightsStore[3][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_653;WeightsStore[3][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_654;WeightsStore[3][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_655;WeightsStore[3][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_656;WeightsStore[3][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_657;WeightsStore[3][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_658;WeightsStore[3][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_659;WeightsStore[3][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_660;WeightsStore[3][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_661;WeightsStore[3][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_662;WeightsStore[3][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_663;WeightsStore[3][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_664;WeightsStore[3][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_665;WeightsStore[3][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_666;WeightsStore[3][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_667;WeightsStore[3][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_668;WeightsStore[3][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_669;WeightsStore[3][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_670;WeightsStore[3][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_671;WeightsStore[3][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_672;WeightsStore[3][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_673;WeightsStore[3][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_674;WeightsStore[3][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_675;WeightsStore[3][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_676;WeightsStore[3][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_677;WeightsStore[3][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_678;WeightsStore[3][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_679;WeightsStore[3][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_680;WeightsStore[3][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_681;WeightsStore[3][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_682;WeightsStore[3][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_683;WeightsStore[3][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_684;WeightsStore[3][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_685;WeightsStore[3][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_686;WeightsStore[3][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_687;WeightsStore[3][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_688;WeightsStore[3][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_689;WeightsStore[3][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_690;WeightsStore[3][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_691;WeightsStore[3][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_692;WeightsStore[3][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_693;WeightsStore[3][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_694;WeightsStore[3][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_695;WeightsStore[3][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_696;WeightsStore[3][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_697;WeightsStore[3][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_698;WeightsStore[3][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_699;WeightsStore[3][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_700;WeightsStore[3][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_701;WeightsStore[3][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_702;WeightsStore[3][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_703;WeightsStore[3][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_704;WeightsStore[3][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_705;WeightsStore[3][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_706;WeightsStore[3][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_707;WeightsStore[3][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_708;WeightsStore[3][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_709;WeightsStore[3][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_710;WeightsStore[3][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_711;WeightsStore[3][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_712;WeightsStore[3][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_713;WeightsStore[3][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_714;WeightsStore[3][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_715;WeightsStore[3][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_716;WeightsStore[3][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_717;WeightsStore[3][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_718;WeightsStore[3][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_719;WeightsStore[3][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_720;WeightsStore[3][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_721;WeightsStore[3][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_722;WeightsStore[3][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_723;WeightsStore[3][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_724;WeightsStore[3][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_725;WeightsStore[3][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_726;WeightsStore[3][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_727;WeightsStore[3][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_728;WeightsStore[3][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_729;WeightsStore[3][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_730;WeightsStore[3][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_731;WeightsStore[3][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_732;WeightsStore[3][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_733;WeightsStore[3][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_734;WeightsStore[3][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_735;WeightsStore[3][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_736;WeightsStore[3][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_737;WeightsStore[3][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_738;WeightsStore[3][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_739;WeightsStore[3][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_740;WeightsStore[3][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_741;WeightsStore[3][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_742;WeightsStore[3][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_743;WeightsStore[3][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_744;WeightsStore[3][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_745;WeightsStore[3][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_746;WeightsStore[3][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_747;WeightsStore[3][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_748;WeightsStore[3][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_749;WeightsStore[3][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_750;WeightsStore[3][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_751;WeightsStore[3][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_752;WeightsStore[3][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_753;WeightsStore[3][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_754;WeightsStore[3][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_755;WeightsStore[3][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_756;WeightsStore[3][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_757;WeightsStore[3][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_758;WeightsStore[3][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_759;WeightsStore[3][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_760;WeightsStore[3][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_761;WeightsStore[3][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_762;WeightsStore[3][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_763;WeightsStore[3][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_764;WeightsStore[3][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_765;WeightsStore[3][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_766;WeightsStore[3][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_767;WeightsStore[3][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_768;WeightsStore[3][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_769;WeightsStore[3][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_770;WeightsStore[3][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_771;WeightsStore[3][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_772;WeightsStore[3][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_773;WeightsStore[3][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_774;WeightsStore[3][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_775;WeightsStore[3][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_776;WeightsStore[3][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_777;WeightsStore[3][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_778;WeightsStore[3][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_779;WeightsStore[3][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_780;WeightsStore[3][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_781;WeightsStore[3][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_782;WeightsStore[3][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_783;WeightsStore[3][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_3_784;WeightsStore[4][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_0;WeightsStore[4][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_1;WeightsStore[4][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_2;WeightsStore[4][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_3;WeightsStore[4][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_4;WeightsStore[4][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_5;WeightsStore[4][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_6;WeightsStore[4][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_7;WeightsStore[4][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_8;WeightsStore[4][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_9;WeightsStore[4][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_10;WeightsStore[4][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_11;WeightsStore[4][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_12;WeightsStore[4][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_13;WeightsStore[4][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_14;WeightsStore[4][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_15;WeightsStore[4][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_16;WeightsStore[4][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_17;WeightsStore[4][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_18;WeightsStore[4][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_19;WeightsStore[4][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_20;WeightsStore[4][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_21;WeightsStore[4][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_22;WeightsStore[4][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_23;WeightsStore[4][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_24;WeightsStore[4][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_25;WeightsStore[4][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_26;WeightsStore[4][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_27;WeightsStore[4][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_28;WeightsStore[4][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_29;WeightsStore[4][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_30;WeightsStore[4][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_31;WeightsStore[4][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_32;WeightsStore[4][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_33;WeightsStore[4][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_34;WeightsStore[4][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_35;WeightsStore[4][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_36;WeightsStore[4][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_37;WeightsStore[4][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_38;WeightsStore[4][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_39;WeightsStore[4][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_40;WeightsStore[4][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_41;WeightsStore[4][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_42;WeightsStore[4][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_43;WeightsStore[4][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_44;WeightsStore[4][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_45;WeightsStore[4][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_46;WeightsStore[4][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_47;WeightsStore[4][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_48;WeightsStore[4][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_49;WeightsStore[4][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_50;WeightsStore[4][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_51;WeightsStore[4][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_52;WeightsStore[4][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_53;WeightsStore[4][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_54;WeightsStore[4][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_55;WeightsStore[4][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_56;WeightsStore[4][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_57;WeightsStore[4][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_58;WeightsStore[4][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_59;WeightsStore[4][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_60;WeightsStore[4][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_61;WeightsStore[4][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_62;WeightsStore[4][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_63;WeightsStore[4][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_64;WeightsStore[4][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_65;WeightsStore[4][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_66;WeightsStore[4][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_67;WeightsStore[4][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_68;WeightsStore[4][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_69;WeightsStore[4][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_70;WeightsStore[4][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_71;WeightsStore[4][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_72;WeightsStore[4][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_73;WeightsStore[4][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_74;WeightsStore[4][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_75;WeightsStore[4][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_76;WeightsStore[4][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_77;WeightsStore[4][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_78;WeightsStore[4][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_79;WeightsStore[4][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_80;WeightsStore[4][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_81;WeightsStore[4][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_82;WeightsStore[4][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_83;WeightsStore[4][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_84;WeightsStore[4][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_85;WeightsStore[4][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_86;WeightsStore[4][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_87;WeightsStore[4][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_88;WeightsStore[4][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_89;WeightsStore[4][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_90;WeightsStore[4][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_91;WeightsStore[4][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_92;WeightsStore[4][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_93;WeightsStore[4][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_94;WeightsStore[4][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_95;WeightsStore[4][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_96;WeightsStore[4][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_97;WeightsStore[4][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_98;WeightsStore[4][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_99;WeightsStore[4][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_100;WeightsStore[4][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_101;WeightsStore[4][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_102;WeightsStore[4][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_103;WeightsStore[4][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_104;WeightsStore[4][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_105;WeightsStore[4][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_106;WeightsStore[4][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_107;WeightsStore[4][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_108;WeightsStore[4][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_109;WeightsStore[4][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_110;WeightsStore[4][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_111;WeightsStore[4][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_112;WeightsStore[4][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_113;WeightsStore[4][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_114;WeightsStore[4][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_115;WeightsStore[4][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_116;WeightsStore[4][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_117;WeightsStore[4][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_118;WeightsStore[4][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_119;WeightsStore[4][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_120;WeightsStore[4][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_121;WeightsStore[4][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_122;WeightsStore[4][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_123;WeightsStore[4][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_124;WeightsStore[4][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_125;WeightsStore[4][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_126;WeightsStore[4][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_127;WeightsStore[4][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_128;WeightsStore[4][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_129;WeightsStore[4][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_130;WeightsStore[4][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_131;WeightsStore[4][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_132;WeightsStore[4][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_133;WeightsStore[4][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_134;WeightsStore[4][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_135;WeightsStore[4][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_136;WeightsStore[4][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_137;WeightsStore[4][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_138;WeightsStore[4][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_139;WeightsStore[4][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_140;WeightsStore[4][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_141;WeightsStore[4][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_142;WeightsStore[4][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_143;WeightsStore[4][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_144;WeightsStore[4][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_145;WeightsStore[4][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_146;WeightsStore[4][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_147;WeightsStore[4][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_148;WeightsStore[4][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_149;WeightsStore[4][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_150;WeightsStore[4][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_151;WeightsStore[4][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_152;WeightsStore[4][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_153;WeightsStore[4][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_154;WeightsStore[4][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_155;WeightsStore[4][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_156;WeightsStore[4][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_157;WeightsStore[4][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_158;WeightsStore[4][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_159;WeightsStore[4][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_160;WeightsStore[4][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_161;WeightsStore[4][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_162;WeightsStore[4][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_163;WeightsStore[4][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_164;WeightsStore[4][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_165;WeightsStore[4][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_166;WeightsStore[4][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_167;WeightsStore[4][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_168;WeightsStore[4][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_169;WeightsStore[4][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_170;WeightsStore[4][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_171;WeightsStore[4][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_172;WeightsStore[4][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_173;WeightsStore[4][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_174;WeightsStore[4][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_175;WeightsStore[4][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_176;WeightsStore[4][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_177;WeightsStore[4][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_178;WeightsStore[4][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_179;WeightsStore[4][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_180;WeightsStore[4][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_181;WeightsStore[4][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_182;WeightsStore[4][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_183;WeightsStore[4][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_184;WeightsStore[4][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_185;WeightsStore[4][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_186;WeightsStore[4][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_187;WeightsStore[4][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_188;WeightsStore[4][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_189;WeightsStore[4][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_190;WeightsStore[4][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_191;WeightsStore[4][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_192;WeightsStore[4][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_193;WeightsStore[4][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_194;WeightsStore[4][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_195;WeightsStore[4][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_196;WeightsStore[4][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_197;WeightsStore[4][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_198;WeightsStore[4][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_199;WeightsStore[4][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_200;WeightsStore[4][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_201;WeightsStore[4][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_202;WeightsStore[4][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_203;WeightsStore[4][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_204;WeightsStore[4][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_205;WeightsStore[4][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_206;WeightsStore[4][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_207;WeightsStore[4][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_208;WeightsStore[4][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_209;WeightsStore[4][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_210;WeightsStore[4][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_211;WeightsStore[4][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_212;WeightsStore[4][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_213;WeightsStore[4][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_214;WeightsStore[4][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_215;WeightsStore[4][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_216;WeightsStore[4][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_217;WeightsStore[4][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_218;WeightsStore[4][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_219;WeightsStore[4][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_220;WeightsStore[4][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_221;WeightsStore[4][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_222;WeightsStore[4][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_223;WeightsStore[4][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_224;WeightsStore[4][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_225;WeightsStore[4][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_226;WeightsStore[4][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_227;WeightsStore[4][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_228;WeightsStore[4][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_229;WeightsStore[4][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_230;WeightsStore[4][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_231;WeightsStore[4][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_232;WeightsStore[4][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_233;WeightsStore[4][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_234;WeightsStore[4][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_235;WeightsStore[4][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_236;WeightsStore[4][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_237;WeightsStore[4][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_238;WeightsStore[4][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_239;WeightsStore[4][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_240;WeightsStore[4][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_241;WeightsStore[4][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_242;WeightsStore[4][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_243;WeightsStore[4][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_244;WeightsStore[4][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_245;WeightsStore[4][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_246;WeightsStore[4][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_247;WeightsStore[4][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_248;WeightsStore[4][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_249;WeightsStore[4][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_250;WeightsStore[4][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_251;WeightsStore[4][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_252;WeightsStore[4][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_253;WeightsStore[4][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_254;WeightsStore[4][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_255;WeightsStore[4][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_256;WeightsStore[4][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_257;WeightsStore[4][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_258;WeightsStore[4][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_259;WeightsStore[4][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_260;WeightsStore[4][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_261;WeightsStore[4][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_262;WeightsStore[4][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_263;WeightsStore[4][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_264;WeightsStore[4][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_265;WeightsStore[4][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_266;WeightsStore[4][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_267;WeightsStore[4][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_268;WeightsStore[4][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_269;WeightsStore[4][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_270;WeightsStore[4][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_271;WeightsStore[4][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_272;WeightsStore[4][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_273;WeightsStore[4][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_274;WeightsStore[4][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_275;WeightsStore[4][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_276;WeightsStore[4][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_277;WeightsStore[4][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_278;WeightsStore[4][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_279;WeightsStore[4][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_280;WeightsStore[4][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_281;WeightsStore[4][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_282;WeightsStore[4][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_283;WeightsStore[4][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_284;WeightsStore[4][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_285;WeightsStore[4][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_286;WeightsStore[4][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_287;WeightsStore[4][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_288;WeightsStore[4][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_289;WeightsStore[4][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_290;WeightsStore[4][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_291;WeightsStore[4][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_292;WeightsStore[4][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_293;WeightsStore[4][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_294;WeightsStore[4][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_295;WeightsStore[4][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_296;WeightsStore[4][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_297;WeightsStore[4][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_298;WeightsStore[4][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_299;WeightsStore[4][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_300;WeightsStore[4][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_301;WeightsStore[4][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_302;WeightsStore[4][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_303;WeightsStore[4][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_304;WeightsStore[4][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_305;WeightsStore[4][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_306;WeightsStore[4][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_307;WeightsStore[4][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_308;WeightsStore[4][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_309;WeightsStore[4][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_310;WeightsStore[4][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_311;WeightsStore[4][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_312;WeightsStore[4][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_313;WeightsStore[4][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_314;WeightsStore[4][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_315;WeightsStore[4][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_316;WeightsStore[4][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_317;WeightsStore[4][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_318;WeightsStore[4][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_319;WeightsStore[4][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_320;WeightsStore[4][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_321;WeightsStore[4][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_322;WeightsStore[4][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_323;WeightsStore[4][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_324;WeightsStore[4][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_325;WeightsStore[4][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_326;WeightsStore[4][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_327;WeightsStore[4][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_328;WeightsStore[4][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_329;WeightsStore[4][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_330;WeightsStore[4][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_331;WeightsStore[4][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_332;WeightsStore[4][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_333;WeightsStore[4][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_334;WeightsStore[4][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_335;WeightsStore[4][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_336;WeightsStore[4][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_337;WeightsStore[4][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_338;WeightsStore[4][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_339;WeightsStore[4][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_340;WeightsStore[4][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_341;WeightsStore[4][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_342;WeightsStore[4][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_343;WeightsStore[4][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_344;WeightsStore[4][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_345;WeightsStore[4][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_346;WeightsStore[4][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_347;WeightsStore[4][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_348;WeightsStore[4][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_349;WeightsStore[4][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_350;WeightsStore[4][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_351;WeightsStore[4][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_352;WeightsStore[4][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_353;WeightsStore[4][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_354;WeightsStore[4][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_355;WeightsStore[4][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_356;WeightsStore[4][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_357;WeightsStore[4][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_358;WeightsStore[4][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_359;WeightsStore[4][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_360;WeightsStore[4][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_361;WeightsStore[4][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_362;WeightsStore[4][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_363;WeightsStore[4][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_364;WeightsStore[4][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_365;WeightsStore[4][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_366;WeightsStore[4][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_367;WeightsStore[4][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_368;WeightsStore[4][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_369;WeightsStore[4][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_370;WeightsStore[4][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_371;WeightsStore[4][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_372;WeightsStore[4][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_373;WeightsStore[4][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_374;WeightsStore[4][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_375;WeightsStore[4][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_376;WeightsStore[4][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_377;WeightsStore[4][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_378;WeightsStore[4][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_379;WeightsStore[4][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_380;WeightsStore[4][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_381;WeightsStore[4][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_382;WeightsStore[4][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_383;WeightsStore[4][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_384;WeightsStore[4][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_385;WeightsStore[4][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_386;WeightsStore[4][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_387;WeightsStore[4][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_388;WeightsStore[4][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_389;WeightsStore[4][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_390;WeightsStore[4][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_391;WeightsStore[4][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_392;WeightsStore[4][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_393;WeightsStore[4][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_394;WeightsStore[4][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_395;WeightsStore[4][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_396;WeightsStore[4][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_397;WeightsStore[4][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_398;WeightsStore[4][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_399;WeightsStore[4][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_400;WeightsStore[4][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_401;WeightsStore[4][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_402;WeightsStore[4][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_403;WeightsStore[4][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_404;WeightsStore[4][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_405;WeightsStore[4][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_406;WeightsStore[4][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_407;WeightsStore[4][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_408;WeightsStore[4][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_409;WeightsStore[4][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_410;WeightsStore[4][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_411;WeightsStore[4][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_412;WeightsStore[4][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_413;WeightsStore[4][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_414;WeightsStore[4][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_415;WeightsStore[4][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_416;WeightsStore[4][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_417;WeightsStore[4][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_418;WeightsStore[4][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_419;WeightsStore[4][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_420;WeightsStore[4][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_421;WeightsStore[4][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_422;WeightsStore[4][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_423;WeightsStore[4][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_424;WeightsStore[4][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_425;WeightsStore[4][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_426;WeightsStore[4][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_427;WeightsStore[4][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_428;WeightsStore[4][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_429;WeightsStore[4][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_430;WeightsStore[4][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_431;WeightsStore[4][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_432;WeightsStore[4][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_433;WeightsStore[4][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_434;WeightsStore[4][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_435;WeightsStore[4][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_436;WeightsStore[4][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_437;WeightsStore[4][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_438;WeightsStore[4][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_439;WeightsStore[4][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_440;WeightsStore[4][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_441;WeightsStore[4][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_442;WeightsStore[4][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_443;WeightsStore[4][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_444;WeightsStore[4][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_445;WeightsStore[4][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_446;WeightsStore[4][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_447;WeightsStore[4][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_448;WeightsStore[4][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_449;WeightsStore[4][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_450;WeightsStore[4][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_451;WeightsStore[4][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_452;WeightsStore[4][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_453;WeightsStore[4][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_454;WeightsStore[4][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_455;WeightsStore[4][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_456;WeightsStore[4][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_457;WeightsStore[4][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_458;WeightsStore[4][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_459;WeightsStore[4][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_460;WeightsStore[4][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_461;WeightsStore[4][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_462;WeightsStore[4][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_463;WeightsStore[4][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_464;WeightsStore[4][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_465;WeightsStore[4][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_466;WeightsStore[4][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_467;WeightsStore[4][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_468;WeightsStore[4][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_469;WeightsStore[4][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_470;WeightsStore[4][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_471;WeightsStore[4][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_472;WeightsStore[4][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_473;WeightsStore[4][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_474;WeightsStore[4][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_475;WeightsStore[4][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_476;WeightsStore[4][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_477;WeightsStore[4][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_478;WeightsStore[4][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_479;WeightsStore[4][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_480;WeightsStore[4][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_481;WeightsStore[4][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_482;WeightsStore[4][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_483;WeightsStore[4][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_484;WeightsStore[4][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_485;WeightsStore[4][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_486;WeightsStore[4][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_487;WeightsStore[4][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_488;WeightsStore[4][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_489;WeightsStore[4][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_490;WeightsStore[4][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_491;WeightsStore[4][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_492;WeightsStore[4][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_493;WeightsStore[4][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_494;WeightsStore[4][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_495;WeightsStore[4][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_496;WeightsStore[4][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_497;WeightsStore[4][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_498;WeightsStore[4][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_499;WeightsStore[4][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_500;WeightsStore[4][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_501;WeightsStore[4][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_502;WeightsStore[4][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_503;WeightsStore[4][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_504;WeightsStore[4][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_505;WeightsStore[4][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_506;WeightsStore[4][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_507;WeightsStore[4][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_508;WeightsStore[4][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_509;WeightsStore[4][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_510;WeightsStore[4][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_511;WeightsStore[4][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_512;WeightsStore[4][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_513;WeightsStore[4][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_514;WeightsStore[4][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_515;WeightsStore[4][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_516;WeightsStore[4][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_517;WeightsStore[4][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_518;WeightsStore[4][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_519;WeightsStore[4][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_520;WeightsStore[4][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_521;WeightsStore[4][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_522;WeightsStore[4][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_523;WeightsStore[4][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_524;WeightsStore[4][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_525;WeightsStore[4][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_526;WeightsStore[4][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_527;WeightsStore[4][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_528;WeightsStore[4][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_529;WeightsStore[4][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_530;WeightsStore[4][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_531;WeightsStore[4][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_532;WeightsStore[4][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_533;WeightsStore[4][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_534;WeightsStore[4][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_535;WeightsStore[4][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_536;WeightsStore[4][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_537;WeightsStore[4][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_538;WeightsStore[4][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_539;WeightsStore[4][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_540;WeightsStore[4][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_541;WeightsStore[4][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_542;WeightsStore[4][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_543;WeightsStore[4][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_544;WeightsStore[4][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_545;WeightsStore[4][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_546;WeightsStore[4][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_547;WeightsStore[4][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_548;WeightsStore[4][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_549;WeightsStore[4][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_550;WeightsStore[4][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_551;WeightsStore[4][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_552;WeightsStore[4][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_553;WeightsStore[4][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_554;WeightsStore[4][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_555;WeightsStore[4][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_556;WeightsStore[4][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_557;WeightsStore[4][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_558;WeightsStore[4][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_559;WeightsStore[4][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_560;WeightsStore[4][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_561;WeightsStore[4][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_562;WeightsStore[4][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_563;WeightsStore[4][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_564;WeightsStore[4][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_565;WeightsStore[4][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_566;WeightsStore[4][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_567;WeightsStore[4][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_568;WeightsStore[4][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_569;WeightsStore[4][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_570;WeightsStore[4][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_571;WeightsStore[4][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_572;WeightsStore[4][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_573;WeightsStore[4][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_574;WeightsStore[4][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_575;WeightsStore[4][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_576;WeightsStore[4][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_577;WeightsStore[4][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_578;WeightsStore[4][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_579;WeightsStore[4][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_580;WeightsStore[4][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_581;WeightsStore[4][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_582;WeightsStore[4][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_583;WeightsStore[4][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_584;WeightsStore[4][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_585;WeightsStore[4][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_586;WeightsStore[4][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_587;WeightsStore[4][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_588;WeightsStore[4][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_589;WeightsStore[4][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_590;WeightsStore[4][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_591;WeightsStore[4][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_592;WeightsStore[4][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_593;WeightsStore[4][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_594;WeightsStore[4][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_595;WeightsStore[4][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_596;WeightsStore[4][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_597;WeightsStore[4][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_598;WeightsStore[4][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_599;WeightsStore[4][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_600;WeightsStore[4][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_601;WeightsStore[4][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_602;WeightsStore[4][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_603;WeightsStore[4][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_604;WeightsStore[4][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_605;WeightsStore[4][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_606;WeightsStore[4][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_607;WeightsStore[4][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_608;WeightsStore[4][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_609;WeightsStore[4][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_610;WeightsStore[4][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_611;WeightsStore[4][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_612;WeightsStore[4][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_613;WeightsStore[4][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_614;WeightsStore[4][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_615;WeightsStore[4][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_616;WeightsStore[4][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_617;WeightsStore[4][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_618;WeightsStore[4][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_619;WeightsStore[4][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_620;WeightsStore[4][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_621;WeightsStore[4][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_622;WeightsStore[4][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_623;WeightsStore[4][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_624;WeightsStore[4][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_625;WeightsStore[4][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_626;WeightsStore[4][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_627;WeightsStore[4][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_628;WeightsStore[4][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_629;WeightsStore[4][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_630;WeightsStore[4][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_631;WeightsStore[4][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_632;WeightsStore[4][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_633;WeightsStore[4][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_634;WeightsStore[4][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_635;WeightsStore[4][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_636;WeightsStore[4][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_637;WeightsStore[4][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_638;WeightsStore[4][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_639;WeightsStore[4][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_640;WeightsStore[4][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_641;WeightsStore[4][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_642;WeightsStore[4][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_643;WeightsStore[4][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_644;WeightsStore[4][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_645;WeightsStore[4][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_646;WeightsStore[4][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_647;WeightsStore[4][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_648;WeightsStore[4][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_649;WeightsStore[4][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_650;WeightsStore[4][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_651;WeightsStore[4][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_652;WeightsStore[4][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_653;WeightsStore[4][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_654;WeightsStore[4][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_655;WeightsStore[4][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_656;WeightsStore[4][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_657;WeightsStore[4][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_658;WeightsStore[4][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_659;WeightsStore[4][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_660;WeightsStore[4][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_661;WeightsStore[4][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_662;WeightsStore[4][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_663;WeightsStore[4][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_664;WeightsStore[4][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_665;WeightsStore[4][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_666;WeightsStore[4][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_667;WeightsStore[4][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_668;WeightsStore[4][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_669;WeightsStore[4][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_670;WeightsStore[4][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_671;WeightsStore[4][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_672;WeightsStore[4][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_673;WeightsStore[4][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_674;WeightsStore[4][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_675;WeightsStore[4][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_676;WeightsStore[4][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_677;WeightsStore[4][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_678;WeightsStore[4][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_679;WeightsStore[4][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_680;WeightsStore[4][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_681;WeightsStore[4][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_682;WeightsStore[4][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_683;WeightsStore[4][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_684;WeightsStore[4][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_685;WeightsStore[4][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_686;WeightsStore[4][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_687;WeightsStore[4][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_688;WeightsStore[4][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_689;WeightsStore[4][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_690;WeightsStore[4][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_691;WeightsStore[4][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_692;WeightsStore[4][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_693;WeightsStore[4][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_694;WeightsStore[4][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_695;WeightsStore[4][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_696;WeightsStore[4][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_697;WeightsStore[4][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_698;WeightsStore[4][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_699;WeightsStore[4][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_700;WeightsStore[4][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_701;WeightsStore[4][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_702;WeightsStore[4][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_703;WeightsStore[4][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_704;WeightsStore[4][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_705;WeightsStore[4][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_706;WeightsStore[4][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_707;WeightsStore[4][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_708;WeightsStore[4][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_709;WeightsStore[4][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_710;WeightsStore[4][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_711;WeightsStore[4][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_712;WeightsStore[4][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_713;WeightsStore[4][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_714;WeightsStore[4][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_715;WeightsStore[4][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_716;WeightsStore[4][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_717;WeightsStore[4][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_718;WeightsStore[4][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_719;WeightsStore[4][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_720;WeightsStore[4][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_721;WeightsStore[4][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_722;WeightsStore[4][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_723;WeightsStore[4][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_724;WeightsStore[4][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_725;WeightsStore[4][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_726;WeightsStore[4][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_727;WeightsStore[4][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_728;WeightsStore[4][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_729;WeightsStore[4][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_730;WeightsStore[4][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_731;WeightsStore[4][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_732;WeightsStore[4][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_733;WeightsStore[4][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_734;WeightsStore[4][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_735;WeightsStore[4][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_736;WeightsStore[4][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_737;WeightsStore[4][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_738;WeightsStore[4][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_739;WeightsStore[4][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_740;WeightsStore[4][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_741;WeightsStore[4][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_742;WeightsStore[4][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_743;WeightsStore[4][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_744;WeightsStore[4][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_745;WeightsStore[4][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_746;WeightsStore[4][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_747;WeightsStore[4][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_748;WeightsStore[4][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_749;WeightsStore[4][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_750;WeightsStore[4][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_751;WeightsStore[4][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_752;WeightsStore[4][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_753;WeightsStore[4][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_754;WeightsStore[4][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_755;WeightsStore[4][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_756;WeightsStore[4][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_757;WeightsStore[4][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_758;WeightsStore[4][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_759;WeightsStore[4][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_760;WeightsStore[4][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_761;WeightsStore[4][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_762;WeightsStore[4][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_763;WeightsStore[4][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_764;WeightsStore[4][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_765;WeightsStore[4][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_766;WeightsStore[4][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_767;WeightsStore[4][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_768;WeightsStore[4][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_769;WeightsStore[4][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_770;WeightsStore[4][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_771;WeightsStore[4][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_772;WeightsStore[4][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_773;WeightsStore[4][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_774;WeightsStore[4][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_775;WeightsStore[4][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_776;WeightsStore[4][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_777;WeightsStore[4][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_778;WeightsStore[4][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_779;WeightsStore[4][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_780;WeightsStore[4][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_781;WeightsStore[4][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_782;WeightsStore[4][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_783;WeightsStore[4][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_4_784;WeightsStore[5][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_0;WeightsStore[5][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_1;WeightsStore[5][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_2;WeightsStore[5][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_3;WeightsStore[5][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_4;WeightsStore[5][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_5;WeightsStore[5][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_6;WeightsStore[5][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_7;WeightsStore[5][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_8;WeightsStore[5][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_9;WeightsStore[5][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_10;WeightsStore[5][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_11;WeightsStore[5][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_12;WeightsStore[5][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_13;WeightsStore[5][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_14;WeightsStore[5][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_15;WeightsStore[5][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_16;WeightsStore[5][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_17;WeightsStore[5][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_18;WeightsStore[5][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_19;WeightsStore[5][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_20;WeightsStore[5][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_21;WeightsStore[5][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_22;WeightsStore[5][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_23;WeightsStore[5][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_24;WeightsStore[5][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_25;WeightsStore[5][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_26;WeightsStore[5][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_27;WeightsStore[5][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_28;WeightsStore[5][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_29;WeightsStore[5][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_30;WeightsStore[5][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_31;WeightsStore[5][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_32;WeightsStore[5][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_33;WeightsStore[5][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_34;WeightsStore[5][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_35;WeightsStore[5][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_36;WeightsStore[5][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_37;WeightsStore[5][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_38;WeightsStore[5][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_39;WeightsStore[5][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_40;WeightsStore[5][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_41;WeightsStore[5][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_42;WeightsStore[5][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_43;WeightsStore[5][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_44;WeightsStore[5][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_45;WeightsStore[5][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_46;WeightsStore[5][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_47;WeightsStore[5][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_48;WeightsStore[5][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_49;WeightsStore[5][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_50;WeightsStore[5][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_51;WeightsStore[5][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_52;WeightsStore[5][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_53;WeightsStore[5][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_54;WeightsStore[5][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_55;WeightsStore[5][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_56;WeightsStore[5][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_57;WeightsStore[5][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_58;WeightsStore[5][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_59;WeightsStore[5][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_60;WeightsStore[5][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_61;WeightsStore[5][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_62;WeightsStore[5][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_63;WeightsStore[5][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_64;WeightsStore[5][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_65;WeightsStore[5][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_66;WeightsStore[5][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_67;WeightsStore[5][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_68;WeightsStore[5][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_69;WeightsStore[5][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_70;WeightsStore[5][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_71;WeightsStore[5][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_72;WeightsStore[5][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_73;WeightsStore[5][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_74;WeightsStore[5][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_75;WeightsStore[5][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_76;WeightsStore[5][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_77;WeightsStore[5][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_78;WeightsStore[5][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_79;WeightsStore[5][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_80;WeightsStore[5][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_81;WeightsStore[5][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_82;WeightsStore[5][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_83;WeightsStore[5][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_84;WeightsStore[5][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_85;WeightsStore[5][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_86;WeightsStore[5][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_87;WeightsStore[5][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_88;WeightsStore[5][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_89;WeightsStore[5][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_90;WeightsStore[5][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_91;WeightsStore[5][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_92;WeightsStore[5][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_93;WeightsStore[5][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_94;WeightsStore[5][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_95;WeightsStore[5][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_96;WeightsStore[5][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_97;WeightsStore[5][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_98;WeightsStore[5][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_99;WeightsStore[5][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_100;WeightsStore[5][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_101;WeightsStore[5][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_102;WeightsStore[5][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_103;WeightsStore[5][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_104;WeightsStore[5][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_105;WeightsStore[5][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_106;WeightsStore[5][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_107;WeightsStore[5][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_108;WeightsStore[5][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_109;WeightsStore[5][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_110;WeightsStore[5][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_111;WeightsStore[5][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_112;WeightsStore[5][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_113;WeightsStore[5][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_114;WeightsStore[5][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_115;WeightsStore[5][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_116;WeightsStore[5][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_117;WeightsStore[5][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_118;WeightsStore[5][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_119;WeightsStore[5][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_120;WeightsStore[5][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_121;WeightsStore[5][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_122;WeightsStore[5][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_123;WeightsStore[5][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_124;WeightsStore[5][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_125;WeightsStore[5][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_126;WeightsStore[5][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_127;WeightsStore[5][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_128;WeightsStore[5][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_129;WeightsStore[5][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_130;WeightsStore[5][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_131;WeightsStore[5][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_132;WeightsStore[5][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_133;WeightsStore[5][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_134;WeightsStore[5][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_135;WeightsStore[5][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_136;WeightsStore[5][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_137;WeightsStore[5][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_138;WeightsStore[5][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_139;WeightsStore[5][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_140;WeightsStore[5][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_141;WeightsStore[5][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_142;WeightsStore[5][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_143;WeightsStore[5][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_144;WeightsStore[5][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_145;WeightsStore[5][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_146;WeightsStore[5][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_147;WeightsStore[5][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_148;WeightsStore[5][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_149;WeightsStore[5][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_150;WeightsStore[5][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_151;WeightsStore[5][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_152;WeightsStore[5][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_153;WeightsStore[5][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_154;WeightsStore[5][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_155;WeightsStore[5][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_156;WeightsStore[5][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_157;WeightsStore[5][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_158;WeightsStore[5][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_159;WeightsStore[5][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_160;WeightsStore[5][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_161;WeightsStore[5][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_162;WeightsStore[5][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_163;WeightsStore[5][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_164;WeightsStore[5][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_165;WeightsStore[5][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_166;WeightsStore[5][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_167;WeightsStore[5][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_168;WeightsStore[5][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_169;WeightsStore[5][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_170;WeightsStore[5][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_171;WeightsStore[5][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_172;WeightsStore[5][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_173;WeightsStore[5][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_174;WeightsStore[5][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_175;WeightsStore[5][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_176;WeightsStore[5][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_177;WeightsStore[5][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_178;WeightsStore[5][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_179;WeightsStore[5][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_180;WeightsStore[5][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_181;WeightsStore[5][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_182;WeightsStore[5][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_183;WeightsStore[5][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_184;WeightsStore[5][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_185;WeightsStore[5][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_186;WeightsStore[5][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_187;WeightsStore[5][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_188;WeightsStore[5][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_189;WeightsStore[5][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_190;WeightsStore[5][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_191;WeightsStore[5][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_192;WeightsStore[5][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_193;WeightsStore[5][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_194;WeightsStore[5][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_195;WeightsStore[5][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_196;WeightsStore[5][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_197;WeightsStore[5][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_198;WeightsStore[5][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_199;WeightsStore[5][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_200;WeightsStore[5][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_201;WeightsStore[5][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_202;WeightsStore[5][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_203;WeightsStore[5][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_204;WeightsStore[5][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_205;WeightsStore[5][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_206;WeightsStore[5][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_207;WeightsStore[5][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_208;WeightsStore[5][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_209;WeightsStore[5][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_210;WeightsStore[5][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_211;WeightsStore[5][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_212;WeightsStore[5][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_213;WeightsStore[5][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_214;WeightsStore[5][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_215;WeightsStore[5][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_216;WeightsStore[5][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_217;WeightsStore[5][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_218;WeightsStore[5][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_219;WeightsStore[5][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_220;WeightsStore[5][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_221;WeightsStore[5][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_222;WeightsStore[5][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_223;WeightsStore[5][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_224;WeightsStore[5][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_225;WeightsStore[5][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_226;WeightsStore[5][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_227;WeightsStore[5][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_228;WeightsStore[5][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_229;WeightsStore[5][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_230;WeightsStore[5][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_231;WeightsStore[5][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_232;WeightsStore[5][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_233;WeightsStore[5][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_234;WeightsStore[5][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_235;WeightsStore[5][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_236;WeightsStore[5][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_237;WeightsStore[5][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_238;WeightsStore[5][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_239;WeightsStore[5][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_240;WeightsStore[5][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_241;WeightsStore[5][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_242;WeightsStore[5][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_243;WeightsStore[5][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_244;WeightsStore[5][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_245;WeightsStore[5][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_246;WeightsStore[5][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_247;WeightsStore[5][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_248;WeightsStore[5][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_249;WeightsStore[5][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_250;WeightsStore[5][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_251;WeightsStore[5][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_252;WeightsStore[5][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_253;WeightsStore[5][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_254;WeightsStore[5][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_255;WeightsStore[5][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_256;WeightsStore[5][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_257;WeightsStore[5][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_258;WeightsStore[5][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_259;WeightsStore[5][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_260;WeightsStore[5][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_261;WeightsStore[5][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_262;WeightsStore[5][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_263;WeightsStore[5][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_264;WeightsStore[5][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_265;WeightsStore[5][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_266;WeightsStore[5][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_267;WeightsStore[5][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_268;WeightsStore[5][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_269;WeightsStore[5][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_270;WeightsStore[5][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_271;WeightsStore[5][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_272;WeightsStore[5][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_273;WeightsStore[5][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_274;WeightsStore[5][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_275;WeightsStore[5][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_276;WeightsStore[5][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_277;WeightsStore[5][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_278;WeightsStore[5][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_279;WeightsStore[5][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_280;WeightsStore[5][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_281;WeightsStore[5][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_282;WeightsStore[5][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_283;WeightsStore[5][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_284;WeightsStore[5][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_285;WeightsStore[5][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_286;WeightsStore[5][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_287;WeightsStore[5][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_288;WeightsStore[5][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_289;WeightsStore[5][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_290;WeightsStore[5][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_291;WeightsStore[5][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_292;WeightsStore[5][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_293;WeightsStore[5][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_294;WeightsStore[5][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_295;WeightsStore[5][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_296;WeightsStore[5][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_297;WeightsStore[5][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_298;WeightsStore[5][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_299;WeightsStore[5][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_300;WeightsStore[5][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_301;WeightsStore[5][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_302;WeightsStore[5][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_303;WeightsStore[5][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_304;WeightsStore[5][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_305;WeightsStore[5][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_306;WeightsStore[5][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_307;WeightsStore[5][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_308;WeightsStore[5][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_309;WeightsStore[5][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_310;WeightsStore[5][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_311;WeightsStore[5][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_312;WeightsStore[5][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_313;WeightsStore[5][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_314;WeightsStore[5][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_315;WeightsStore[5][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_316;WeightsStore[5][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_317;WeightsStore[5][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_318;WeightsStore[5][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_319;WeightsStore[5][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_320;WeightsStore[5][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_321;WeightsStore[5][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_322;WeightsStore[5][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_323;WeightsStore[5][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_324;WeightsStore[5][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_325;WeightsStore[5][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_326;WeightsStore[5][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_327;WeightsStore[5][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_328;WeightsStore[5][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_329;WeightsStore[5][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_330;WeightsStore[5][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_331;WeightsStore[5][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_332;WeightsStore[5][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_333;WeightsStore[5][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_334;WeightsStore[5][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_335;WeightsStore[5][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_336;WeightsStore[5][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_337;WeightsStore[5][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_338;WeightsStore[5][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_339;WeightsStore[5][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_340;WeightsStore[5][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_341;WeightsStore[5][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_342;WeightsStore[5][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_343;WeightsStore[5][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_344;WeightsStore[5][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_345;WeightsStore[5][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_346;WeightsStore[5][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_347;WeightsStore[5][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_348;WeightsStore[5][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_349;WeightsStore[5][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_350;WeightsStore[5][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_351;WeightsStore[5][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_352;WeightsStore[5][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_353;WeightsStore[5][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_354;WeightsStore[5][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_355;WeightsStore[5][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_356;WeightsStore[5][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_357;WeightsStore[5][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_358;WeightsStore[5][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_359;WeightsStore[5][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_360;WeightsStore[5][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_361;WeightsStore[5][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_362;WeightsStore[5][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_363;WeightsStore[5][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_364;WeightsStore[5][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_365;WeightsStore[5][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_366;WeightsStore[5][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_367;WeightsStore[5][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_368;WeightsStore[5][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_369;WeightsStore[5][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_370;WeightsStore[5][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_371;WeightsStore[5][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_372;WeightsStore[5][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_373;WeightsStore[5][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_374;WeightsStore[5][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_375;WeightsStore[5][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_376;WeightsStore[5][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_377;WeightsStore[5][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_378;WeightsStore[5][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_379;WeightsStore[5][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_380;WeightsStore[5][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_381;WeightsStore[5][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_382;WeightsStore[5][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_383;WeightsStore[5][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_384;WeightsStore[5][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_385;WeightsStore[5][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_386;WeightsStore[5][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_387;WeightsStore[5][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_388;WeightsStore[5][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_389;WeightsStore[5][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_390;WeightsStore[5][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_391;WeightsStore[5][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_392;WeightsStore[5][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_393;WeightsStore[5][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_394;WeightsStore[5][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_395;WeightsStore[5][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_396;WeightsStore[5][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_397;WeightsStore[5][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_398;WeightsStore[5][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_399;WeightsStore[5][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_400;WeightsStore[5][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_401;WeightsStore[5][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_402;WeightsStore[5][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_403;WeightsStore[5][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_404;WeightsStore[5][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_405;WeightsStore[5][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_406;WeightsStore[5][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_407;WeightsStore[5][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_408;WeightsStore[5][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_409;WeightsStore[5][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_410;WeightsStore[5][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_411;WeightsStore[5][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_412;WeightsStore[5][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_413;WeightsStore[5][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_414;WeightsStore[5][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_415;WeightsStore[5][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_416;WeightsStore[5][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_417;WeightsStore[5][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_418;WeightsStore[5][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_419;WeightsStore[5][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_420;WeightsStore[5][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_421;WeightsStore[5][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_422;WeightsStore[5][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_423;WeightsStore[5][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_424;WeightsStore[5][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_425;WeightsStore[5][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_426;WeightsStore[5][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_427;WeightsStore[5][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_428;WeightsStore[5][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_429;WeightsStore[5][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_430;WeightsStore[5][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_431;WeightsStore[5][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_432;WeightsStore[5][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_433;WeightsStore[5][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_434;WeightsStore[5][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_435;WeightsStore[5][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_436;WeightsStore[5][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_437;WeightsStore[5][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_438;WeightsStore[5][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_439;WeightsStore[5][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_440;WeightsStore[5][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_441;WeightsStore[5][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_442;WeightsStore[5][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_443;WeightsStore[5][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_444;WeightsStore[5][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_445;WeightsStore[5][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_446;WeightsStore[5][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_447;WeightsStore[5][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_448;WeightsStore[5][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_449;WeightsStore[5][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_450;WeightsStore[5][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_451;WeightsStore[5][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_452;WeightsStore[5][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_453;WeightsStore[5][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_454;WeightsStore[5][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_455;WeightsStore[5][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_456;WeightsStore[5][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_457;WeightsStore[5][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_458;WeightsStore[5][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_459;WeightsStore[5][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_460;WeightsStore[5][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_461;WeightsStore[5][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_462;WeightsStore[5][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_463;WeightsStore[5][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_464;WeightsStore[5][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_465;WeightsStore[5][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_466;WeightsStore[5][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_467;WeightsStore[5][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_468;WeightsStore[5][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_469;WeightsStore[5][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_470;WeightsStore[5][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_471;WeightsStore[5][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_472;WeightsStore[5][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_473;WeightsStore[5][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_474;WeightsStore[5][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_475;WeightsStore[5][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_476;WeightsStore[5][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_477;WeightsStore[5][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_478;WeightsStore[5][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_479;WeightsStore[5][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_480;WeightsStore[5][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_481;WeightsStore[5][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_482;WeightsStore[5][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_483;WeightsStore[5][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_484;WeightsStore[5][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_485;WeightsStore[5][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_486;WeightsStore[5][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_487;WeightsStore[5][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_488;WeightsStore[5][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_489;WeightsStore[5][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_490;WeightsStore[5][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_491;WeightsStore[5][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_492;WeightsStore[5][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_493;WeightsStore[5][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_494;WeightsStore[5][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_495;WeightsStore[5][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_496;WeightsStore[5][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_497;WeightsStore[5][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_498;WeightsStore[5][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_499;WeightsStore[5][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_500;WeightsStore[5][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_501;WeightsStore[5][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_502;WeightsStore[5][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_503;WeightsStore[5][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_504;WeightsStore[5][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_505;WeightsStore[5][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_506;WeightsStore[5][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_507;WeightsStore[5][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_508;WeightsStore[5][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_509;WeightsStore[5][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_510;WeightsStore[5][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_511;WeightsStore[5][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_512;WeightsStore[5][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_513;WeightsStore[5][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_514;WeightsStore[5][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_515;WeightsStore[5][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_516;WeightsStore[5][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_517;WeightsStore[5][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_518;WeightsStore[5][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_519;WeightsStore[5][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_520;WeightsStore[5][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_521;WeightsStore[5][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_522;WeightsStore[5][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_523;WeightsStore[5][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_524;WeightsStore[5][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_525;WeightsStore[5][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_526;WeightsStore[5][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_527;WeightsStore[5][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_528;WeightsStore[5][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_529;WeightsStore[5][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_530;WeightsStore[5][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_531;WeightsStore[5][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_532;WeightsStore[5][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_533;WeightsStore[5][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_534;WeightsStore[5][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_535;WeightsStore[5][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_536;WeightsStore[5][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_537;WeightsStore[5][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_538;WeightsStore[5][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_539;WeightsStore[5][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_540;WeightsStore[5][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_541;WeightsStore[5][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_542;WeightsStore[5][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_543;WeightsStore[5][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_544;WeightsStore[5][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_545;WeightsStore[5][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_546;WeightsStore[5][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_547;WeightsStore[5][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_548;WeightsStore[5][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_549;WeightsStore[5][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_550;WeightsStore[5][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_551;WeightsStore[5][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_552;WeightsStore[5][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_553;WeightsStore[5][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_554;WeightsStore[5][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_555;WeightsStore[5][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_556;WeightsStore[5][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_557;WeightsStore[5][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_558;WeightsStore[5][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_559;WeightsStore[5][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_560;WeightsStore[5][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_561;WeightsStore[5][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_562;WeightsStore[5][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_563;WeightsStore[5][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_564;WeightsStore[5][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_565;WeightsStore[5][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_566;WeightsStore[5][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_567;WeightsStore[5][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_568;WeightsStore[5][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_569;WeightsStore[5][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_570;WeightsStore[5][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_571;WeightsStore[5][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_572;WeightsStore[5][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_573;WeightsStore[5][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_574;WeightsStore[5][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_575;WeightsStore[5][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_576;WeightsStore[5][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_577;WeightsStore[5][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_578;WeightsStore[5][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_579;WeightsStore[5][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_580;WeightsStore[5][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_581;WeightsStore[5][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_582;WeightsStore[5][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_583;WeightsStore[5][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_584;WeightsStore[5][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_585;WeightsStore[5][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_586;WeightsStore[5][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_587;WeightsStore[5][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_588;WeightsStore[5][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_589;WeightsStore[5][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_590;WeightsStore[5][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_591;WeightsStore[5][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_592;WeightsStore[5][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_593;WeightsStore[5][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_594;WeightsStore[5][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_595;WeightsStore[5][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_596;WeightsStore[5][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_597;WeightsStore[5][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_598;WeightsStore[5][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_599;WeightsStore[5][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_600;WeightsStore[5][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_601;WeightsStore[5][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_602;WeightsStore[5][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_603;WeightsStore[5][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_604;WeightsStore[5][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_605;WeightsStore[5][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_606;WeightsStore[5][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_607;WeightsStore[5][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_608;WeightsStore[5][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_609;WeightsStore[5][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_610;WeightsStore[5][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_611;WeightsStore[5][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_612;WeightsStore[5][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_613;WeightsStore[5][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_614;WeightsStore[5][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_615;WeightsStore[5][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_616;WeightsStore[5][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_617;WeightsStore[5][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_618;WeightsStore[5][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_619;WeightsStore[5][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_620;WeightsStore[5][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_621;WeightsStore[5][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_622;WeightsStore[5][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_623;WeightsStore[5][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_624;WeightsStore[5][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_625;WeightsStore[5][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_626;WeightsStore[5][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_627;WeightsStore[5][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_628;WeightsStore[5][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_629;WeightsStore[5][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_630;WeightsStore[5][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_631;WeightsStore[5][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_632;WeightsStore[5][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_633;WeightsStore[5][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_634;WeightsStore[5][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_635;WeightsStore[5][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_636;WeightsStore[5][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_637;WeightsStore[5][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_638;WeightsStore[5][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_639;WeightsStore[5][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_640;WeightsStore[5][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_641;WeightsStore[5][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_642;WeightsStore[5][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_643;WeightsStore[5][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_644;WeightsStore[5][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_645;WeightsStore[5][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_646;WeightsStore[5][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_647;WeightsStore[5][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_648;WeightsStore[5][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_649;WeightsStore[5][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_650;WeightsStore[5][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_651;WeightsStore[5][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_652;WeightsStore[5][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_653;WeightsStore[5][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_654;WeightsStore[5][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_655;WeightsStore[5][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_656;WeightsStore[5][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_657;WeightsStore[5][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_658;WeightsStore[5][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_659;WeightsStore[5][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_660;WeightsStore[5][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_661;WeightsStore[5][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_662;WeightsStore[5][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_663;WeightsStore[5][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_664;WeightsStore[5][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_665;WeightsStore[5][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_666;WeightsStore[5][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_667;WeightsStore[5][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_668;WeightsStore[5][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_669;WeightsStore[5][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_670;WeightsStore[5][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_671;WeightsStore[5][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_672;WeightsStore[5][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_673;WeightsStore[5][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_674;WeightsStore[5][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_675;WeightsStore[5][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_676;WeightsStore[5][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_677;WeightsStore[5][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_678;WeightsStore[5][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_679;WeightsStore[5][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_680;WeightsStore[5][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_681;WeightsStore[5][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_682;WeightsStore[5][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_683;WeightsStore[5][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_684;WeightsStore[5][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_685;WeightsStore[5][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_686;WeightsStore[5][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_687;WeightsStore[5][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_688;WeightsStore[5][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_689;WeightsStore[5][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_690;WeightsStore[5][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_691;WeightsStore[5][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_692;WeightsStore[5][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_693;WeightsStore[5][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_694;WeightsStore[5][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_695;WeightsStore[5][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_696;WeightsStore[5][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_697;WeightsStore[5][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_698;WeightsStore[5][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_699;WeightsStore[5][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_700;WeightsStore[5][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_701;WeightsStore[5][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_702;WeightsStore[5][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_703;WeightsStore[5][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_704;WeightsStore[5][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_705;WeightsStore[5][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_706;WeightsStore[5][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_707;WeightsStore[5][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_708;WeightsStore[5][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_709;WeightsStore[5][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_710;WeightsStore[5][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_711;WeightsStore[5][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_712;WeightsStore[5][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_713;WeightsStore[5][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_714;WeightsStore[5][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_715;WeightsStore[5][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_716;WeightsStore[5][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_717;WeightsStore[5][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_718;WeightsStore[5][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_719;WeightsStore[5][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_720;WeightsStore[5][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_721;WeightsStore[5][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_722;WeightsStore[5][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_723;WeightsStore[5][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_724;WeightsStore[5][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_725;WeightsStore[5][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_726;WeightsStore[5][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_727;WeightsStore[5][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_728;WeightsStore[5][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_729;WeightsStore[5][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_730;WeightsStore[5][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_731;WeightsStore[5][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_732;WeightsStore[5][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_733;WeightsStore[5][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_734;WeightsStore[5][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_735;WeightsStore[5][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_736;WeightsStore[5][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_737;WeightsStore[5][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_738;WeightsStore[5][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_739;WeightsStore[5][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_740;WeightsStore[5][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_741;WeightsStore[5][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_742;WeightsStore[5][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_743;WeightsStore[5][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_744;WeightsStore[5][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_745;WeightsStore[5][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_746;WeightsStore[5][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_747;WeightsStore[5][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_748;WeightsStore[5][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_749;WeightsStore[5][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_750;WeightsStore[5][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_751;WeightsStore[5][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_752;WeightsStore[5][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_753;WeightsStore[5][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_754;WeightsStore[5][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_755;WeightsStore[5][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_756;WeightsStore[5][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_757;WeightsStore[5][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_758;WeightsStore[5][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_759;WeightsStore[5][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_760;WeightsStore[5][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_761;WeightsStore[5][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_762;WeightsStore[5][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_763;WeightsStore[5][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_764;WeightsStore[5][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_765;WeightsStore[5][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_766;WeightsStore[5][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_767;WeightsStore[5][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_768;WeightsStore[5][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_769;WeightsStore[5][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_770;WeightsStore[5][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_771;WeightsStore[5][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_772;WeightsStore[5][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_773;WeightsStore[5][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_774;WeightsStore[5][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_775;WeightsStore[5][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_776;WeightsStore[5][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_777;WeightsStore[5][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_778;WeightsStore[5][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_779;WeightsStore[5][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_780;WeightsStore[5][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_781;WeightsStore[5][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_782;WeightsStore[5][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_783;WeightsStore[5][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_5_784;WeightsStore[6][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_0;WeightsStore[6][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_1;WeightsStore[6][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_2;WeightsStore[6][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_3;WeightsStore[6][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_4;WeightsStore[6][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_5;WeightsStore[6][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_6;WeightsStore[6][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_7;WeightsStore[6][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_8;WeightsStore[6][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_9;WeightsStore[6][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_10;WeightsStore[6][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_11;WeightsStore[6][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_12;WeightsStore[6][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_13;WeightsStore[6][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_14;WeightsStore[6][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_15;WeightsStore[6][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_16;WeightsStore[6][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_17;WeightsStore[6][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_18;WeightsStore[6][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_19;WeightsStore[6][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_20;WeightsStore[6][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_21;WeightsStore[6][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_22;WeightsStore[6][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_23;WeightsStore[6][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_24;WeightsStore[6][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_25;WeightsStore[6][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_26;WeightsStore[6][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_27;WeightsStore[6][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_28;WeightsStore[6][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_29;WeightsStore[6][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_30;WeightsStore[6][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_31;WeightsStore[6][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_32;WeightsStore[6][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_33;WeightsStore[6][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_34;WeightsStore[6][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_35;WeightsStore[6][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_36;WeightsStore[6][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_37;WeightsStore[6][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_38;WeightsStore[6][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_39;WeightsStore[6][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_40;WeightsStore[6][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_41;WeightsStore[6][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_42;WeightsStore[6][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_43;WeightsStore[6][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_44;WeightsStore[6][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_45;WeightsStore[6][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_46;WeightsStore[6][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_47;WeightsStore[6][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_48;WeightsStore[6][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_49;WeightsStore[6][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_50;WeightsStore[6][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_51;WeightsStore[6][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_52;WeightsStore[6][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_53;WeightsStore[6][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_54;WeightsStore[6][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_55;WeightsStore[6][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_56;WeightsStore[6][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_57;WeightsStore[6][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_58;WeightsStore[6][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_59;WeightsStore[6][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_60;WeightsStore[6][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_61;WeightsStore[6][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_62;WeightsStore[6][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_63;WeightsStore[6][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_64;WeightsStore[6][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_65;WeightsStore[6][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_66;WeightsStore[6][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_67;WeightsStore[6][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_68;WeightsStore[6][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_69;WeightsStore[6][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_70;WeightsStore[6][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_71;WeightsStore[6][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_72;WeightsStore[6][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_73;WeightsStore[6][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_74;WeightsStore[6][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_75;WeightsStore[6][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_76;WeightsStore[6][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_77;WeightsStore[6][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_78;WeightsStore[6][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_79;WeightsStore[6][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_80;WeightsStore[6][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_81;WeightsStore[6][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_82;WeightsStore[6][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_83;WeightsStore[6][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_84;WeightsStore[6][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_85;WeightsStore[6][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_86;WeightsStore[6][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_87;WeightsStore[6][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_88;WeightsStore[6][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_89;WeightsStore[6][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_90;WeightsStore[6][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_91;WeightsStore[6][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_92;WeightsStore[6][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_93;WeightsStore[6][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_94;WeightsStore[6][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_95;WeightsStore[6][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_96;WeightsStore[6][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_97;WeightsStore[6][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_98;WeightsStore[6][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_99;WeightsStore[6][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_100;WeightsStore[6][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_101;WeightsStore[6][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_102;WeightsStore[6][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_103;WeightsStore[6][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_104;WeightsStore[6][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_105;WeightsStore[6][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_106;WeightsStore[6][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_107;WeightsStore[6][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_108;WeightsStore[6][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_109;WeightsStore[6][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_110;WeightsStore[6][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_111;WeightsStore[6][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_112;WeightsStore[6][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_113;WeightsStore[6][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_114;WeightsStore[6][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_115;WeightsStore[6][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_116;WeightsStore[6][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_117;WeightsStore[6][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_118;WeightsStore[6][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_119;WeightsStore[6][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_120;WeightsStore[6][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_121;WeightsStore[6][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_122;WeightsStore[6][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_123;WeightsStore[6][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_124;WeightsStore[6][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_125;WeightsStore[6][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_126;WeightsStore[6][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_127;WeightsStore[6][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_128;WeightsStore[6][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_129;WeightsStore[6][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_130;WeightsStore[6][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_131;WeightsStore[6][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_132;WeightsStore[6][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_133;WeightsStore[6][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_134;WeightsStore[6][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_135;WeightsStore[6][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_136;WeightsStore[6][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_137;WeightsStore[6][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_138;WeightsStore[6][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_139;WeightsStore[6][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_140;WeightsStore[6][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_141;WeightsStore[6][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_142;WeightsStore[6][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_143;WeightsStore[6][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_144;WeightsStore[6][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_145;WeightsStore[6][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_146;WeightsStore[6][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_147;WeightsStore[6][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_148;WeightsStore[6][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_149;WeightsStore[6][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_150;WeightsStore[6][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_151;WeightsStore[6][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_152;WeightsStore[6][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_153;WeightsStore[6][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_154;WeightsStore[6][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_155;WeightsStore[6][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_156;WeightsStore[6][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_157;WeightsStore[6][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_158;WeightsStore[6][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_159;WeightsStore[6][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_160;WeightsStore[6][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_161;WeightsStore[6][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_162;WeightsStore[6][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_163;WeightsStore[6][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_164;WeightsStore[6][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_165;WeightsStore[6][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_166;WeightsStore[6][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_167;WeightsStore[6][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_168;WeightsStore[6][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_169;WeightsStore[6][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_170;WeightsStore[6][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_171;WeightsStore[6][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_172;WeightsStore[6][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_173;WeightsStore[6][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_174;WeightsStore[6][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_175;WeightsStore[6][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_176;WeightsStore[6][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_177;WeightsStore[6][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_178;WeightsStore[6][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_179;WeightsStore[6][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_180;WeightsStore[6][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_181;WeightsStore[6][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_182;WeightsStore[6][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_183;WeightsStore[6][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_184;WeightsStore[6][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_185;WeightsStore[6][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_186;WeightsStore[6][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_187;WeightsStore[6][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_188;WeightsStore[6][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_189;WeightsStore[6][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_190;WeightsStore[6][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_191;WeightsStore[6][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_192;WeightsStore[6][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_193;WeightsStore[6][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_194;WeightsStore[6][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_195;WeightsStore[6][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_196;WeightsStore[6][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_197;WeightsStore[6][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_198;WeightsStore[6][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_199;WeightsStore[6][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_200;WeightsStore[6][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_201;WeightsStore[6][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_202;WeightsStore[6][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_203;WeightsStore[6][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_204;WeightsStore[6][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_205;WeightsStore[6][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_206;WeightsStore[6][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_207;WeightsStore[6][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_208;WeightsStore[6][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_209;WeightsStore[6][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_210;WeightsStore[6][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_211;WeightsStore[6][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_212;WeightsStore[6][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_213;WeightsStore[6][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_214;WeightsStore[6][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_215;WeightsStore[6][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_216;WeightsStore[6][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_217;WeightsStore[6][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_218;WeightsStore[6][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_219;WeightsStore[6][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_220;WeightsStore[6][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_221;WeightsStore[6][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_222;WeightsStore[6][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_223;WeightsStore[6][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_224;WeightsStore[6][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_225;WeightsStore[6][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_226;WeightsStore[6][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_227;WeightsStore[6][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_228;WeightsStore[6][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_229;WeightsStore[6][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_230;WeightsStore[6][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_231;WeightsStore[6][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_232;WeightsStore[6][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_233;WeightsStore[6][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_234;WeightsStore[6][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_235;WeightsStore[6][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_236;WeightsStore[6][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_237;WeightsStore[6][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_238;WeightsStore[6][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_239;WeightsStore[6][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_240;WeightsStore[6][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_241;WeightsStore[6][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_242;WeightsStore[6][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_243;WeightsStore[6][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_244;WeightsStore[6][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_245;WeightsStore[6][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_246;WeightsStore[6][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_247;WeightsStore[6][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_248;WeightsStore[6][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_249;WeightsStore[6][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_250;WeightsStore[6][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_251;WeightsStore[6][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_252;WeightsStore[6][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_253;WeightsStore[6][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_254;WeightsStore[6][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_255;WeightsStore[6][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_256;WeightsStore[6][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_257;WeightsStore[6][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_258;WeightsStore[6][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_259;WeightsStore[6][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_260;WeightsStore[6][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_261;WeightsStore[6][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_262;WeightsStore[6][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_263;WeightsStore[6][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_264;WeightsStore[6][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_265;WeightsStore[6][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_266;WeightsStore[6][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_267;WeightsStore[6][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_268;WeightsStore[6][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_269;WeightsStore[6][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_270;WeightsStore[6][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_271;WeightsStore[6][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_272;WeightsStore[6][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_273;WeightsStore[6][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_274;WeightsStore[6][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_275;WeightsStore[6][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_276;WeightsStore[6][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_277;WeightsStore[6][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_278;WeightsStore[6][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_279;WeightsStore[6][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_280;WeightsStore[6][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_281;WeightsStore[6][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_282;WeightsStore[6][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_283;WeightsStore[6][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_284;WeightsStore[6][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_285;WeightsStore[6][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_286;WeightsStore[6][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_287;WeightsStore[6][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_288;WeightsStore[6][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_289;WeightsStore[6][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_290;WeightsStore[6][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_291;WeightsStore[6][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_292;WeightsStore[6][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_293;WeightsStore[6][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_294;WeightsStore[6][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_295;WeightsStore[6][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_296;WeightsStore[6][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_297;WeightsStore[6][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_298;WeightsStore[6][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_299;WeightsStore[6][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_300;WeightsStore[6][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_301;WeightsStore[6][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_302;WeightsStore[6][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_303;WeightsStore[6][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_304;WeightsStore[6][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_305;WeightsStore[6][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_306;WeightsStore[6][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_307;WeightsStore[6][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_308;WeightsStore[6][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_309;WeightsStore[6][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_310;WeightsStore[6][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_311;WeightsStore[6][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_312;WeightsStore[6][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_313;WeightsStore[6][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_314;WeightsStore[6][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_315;WeightsStore[6][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_316;WeightsStore[6][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_317;WeightsStore[6][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_318;WeightsStore[6][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_319;WeightsStore[6][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_320;WeightsStore[6][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_321;WeightsStore[6][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_322;WeightsStore[6][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_323;WeightsStore[6][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_324;WeightsStore[6][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_325;WeightsStore[6][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_326;WeightsStore[6][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_327;WeightsStore[6][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_328;WeightsStore[6][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_329;WeightsStore[6][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_330;WeightsStore[6][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_331;WeightsStore[6][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_332;WeightsStore[6][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_333;WeightsStore[6][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_334;WeightsStore[6][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_335;WeightsStore[6][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_336;WeightsStore[6][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_337;WeightsStore[6][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_338;WeightsStore[6][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_339;WeightsStore[6][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_340;WeightsStore[6][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_341;WeightsStore[6][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_342;WeightsStore[6][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_343;WeightsStore[6][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_344;WeightsStore[6][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_345;WeightsStore[6][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_346;WeightsStore[6][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_347;WeightsStore[6][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_348;WeightsStore[6][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_349;WeightsStore[6][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_350;WeightsStore[6][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_351;WeightsStore[6][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_352;WeightsStore[6][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_353;WeightsStore[6][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_354;WeightsStore[6][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_355;WeightsStore[6][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_356;WeightsStore[6][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_357;WeightsStore[6][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_358;WeightsStore[6][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_359;WeightsStore[6][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_360;WeightsStore[6][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_361;WeightsStore[6][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_362;WeightsStore[6][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_363;WeightsStore[6][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_364;WeightsStore[6][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_365;WeightsStore[6][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_366;WeightsStore[6][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_367;WeightsStore[6][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_368;WeightsStore[6][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_369;WeightsStore[6][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_370;WeightsStore[6][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_371;WeightsStore[6][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_372;WeightsStore[6][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_373;WeightsStore[6][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_374;WeightsStore[6][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_375;WeightsStore[6][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_376;WeightsStore[6][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_377;WeightsStore[6][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_378;WeightsStore[6][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_379;WeightsStore[6][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_380;WeightsStore[6][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_381;WeightsStore[6][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_382;WeightsStore[6][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_383;WeightsStore[6][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_384;WeightsStore[6][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_385;WeightsStore[6][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_386;WeightsStore[6][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_387;WeightsStore[6][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_388;WeightsStore[6][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_389;WeightsStore[6][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_390;WeightsStore[6][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_391;WeightsStore[6][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_392;WeightsStore[6][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_393;WeightsStore[6][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_394;WeightsStore[6][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_395;WeightsStore[6][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_396;WeightsStore[6][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_397;WeightsStore[6][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_398;WeightsStore[6][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_399;WeightsStore[6][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_400;WeightsStore[6][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_401;WeightsStore[6][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_402;WeightsStore[6][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_403;WeightsStore[6][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_404;WeightsStore[6][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_405;WeightsStore[6][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_406;WeightsStore[6][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_407;WeightsStore[6][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_408;WeightsStore[6][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_409;WeightsStore[6][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_410;WeightsStore[6][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_411;WeightsStore[6][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_412;WeightsStore[6][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_413;WeightsStore[6][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_414;WeightsStore[6][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_415;WeightsStore[6][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_416;WeightsStore[6][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_417;WeightsStore[6][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_418;WeightsStore[6][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_419;WeightsStore[6][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_420;WeightsStore[6][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_421;WeightsStore[6][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_422;WeightsStore[6][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_423;WeightsStore[6][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_424;WeightsStore[6][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_425;WeightsStore[6][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_426;WeightsStore[6][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_427;WeightsStore[6][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_428;WeightsStore[6][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_429;WeightsStore[6][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_430;WeightsStore[6][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_431;WeightsStore[6][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_432;WeightsStore[6][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_433;WeightsStore[6][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_434;WeightsStore[6][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_435;WeightsStore[6][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_436;WeightsStore[6][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_437;WeightsStore[6][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_438;WeightsStore[6][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_439;WeightsStore[6][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_440;WeightsStore[6][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_441;WeightsStore[6][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_442;WeightsStore[6][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_443;WeightsStore[6][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_444;WeightsStore[6][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_445;WeightsStore[6][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_446;WeightsStore[6][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_447;WeightsStore[6][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_448;WeightsStore[6][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_449;WeightsStore[6][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_450;WeightsStore[6][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_451;WeightsStore[6][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_452;WeightsStore[6][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_453;WeightsStore[6][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_454;WeightsStore[6][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_455;WeightsStore[6][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_456;WeightsStore[6][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_457;WeightsStore[6][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_458;WeightsStore[6][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_459;WeightsStore[6][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_460;WeightsStore[6][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_461;WeightsStore[6][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_462;WeightsStore[6][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_463;WeightsStore[6][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_464;WeightsStore[6][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_465;WeightsStore[6][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_466;WeightsStore[6][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_467;WeightsStore[6][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_468;WeightsStore[6][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_469;WeightsStore[6][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_470;WeightsStore[6][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_471;WeightsStore[6][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_472;WeightsStore[6][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_473;WeightsStore[6][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_474;WeightsStore[6][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_475;WeightsStore[6][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_476;WeightsStore[6][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_477;WeightsStore[6][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_478;WeightsStore[6][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_479;WeightsStore[6][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_480;WeightsStore[6][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_481;WeightsStore[6][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_482;WeightsStore[6][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_483;WeightsStore[6][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_484;WeightsStore[6][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_485;WeightsStore[6][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_486;WeightsStore[6][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_487;WeightsStore[6][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_488;WeightsStore[6][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_489;WeightsStore[6][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_490;WeightsStore[6][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_491;WeightsStore[6][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_492;WeightsStore[6][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_493;WeightsStore[6][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_494;WeightsStore[6][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_495;WeightsStore[6][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_496;WeightsStore[6][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_497;WeightsStore[6][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_498;WeightsStore[6][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_499;WeightsStore[6][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_500;WeightsStore[6][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_501;WeightsStore[6][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_502;WeightsStore[6][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_503;WeightsStore[6][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_504;WeightsStore[6][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_505;WeightsStore[6][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_506;WeightsStore[6][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_507;WeightsStore[6][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_508;WeightsStore[6][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_509;WeightsStore[6][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_510;WeightsStore[6][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_511;WeightsStore[6][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_512;WeightsStore[6][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_513;WeightsStore[6][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_514;WeightsStore[6][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_515;WeightsStore[6][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_516;WeightsStore[6][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_517;WeightsStore[6][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_518;WeightsStore[6][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_519;WeightsStore[6][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_520;WeightsStore[6][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_521;WeightsStore[6][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_522;WeightsStore[6][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_523;WeightsStore[6][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_524;WeightsStore[6][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_525;WeightsStore[6][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_526;WeightsStore[6][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_527;WeightsStore[6][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_528;WeightsStore[6][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_529;WeightsStore[6][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_530;WeightsStore[6][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_531;WeightsStore[6][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_532;WeightsStore[6][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_533;WeightsStore[6][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_534;WeightsStore[6][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_535;WeightsStore[6][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_536;WeightsStore[6][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_537;WeightsStore[6][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_538;WeightsStore[6][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_539;WeightsStore[6][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_540;WeightsStore[6][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_541;WeightsStore[6][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_542;WeightsStore[6][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_543;WeightsStore[6][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_544;WeightsStore[6][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_545;WeightsStore[6][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_546;WeightsStore[6][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_547;WeightsStore[6][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_548;WeightsStore[6][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_549;WeightsStore[6][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_550;WeightsStore[6][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_551;WeightsStore[6][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_552;WeightsStore[6][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_553;WeightsStore[6][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_554;WeightsStore[6][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_555;WeightsStore[6][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_556;WeightsStore[6][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_557;WeightsStore[6][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_558;WeightsStore[6][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_559;WeightsStore[6][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_560;WeightsStore[6][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_561;WeightsStore[6][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_562;WeightsStore[6][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_563;WeightsStore[6][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_564;WeightsStore[6][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_565;WeightsStore[6][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_566;WeightsStore[6][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_567;WeightsStore[6][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_568;WeightsStore[6][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_569;WeightsStore[6][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_570;WeightsStore[6][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_571;WeightsStore[6][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_572;WeightsStore[6][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_573;WeightsStore[6][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_574;WeightsStore[6][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_575;WeightsStore[6][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_576;WeightsStore[6][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_577;WeightsStore[6][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_578;WeightsStore[6][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_579;WeightsStore[6][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_580;WeightsStore[6][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_581;WeightsStore[6][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_582;WeightsStore[6][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_583;WeightsStore[6][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_584;WeightsStore[6][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_585;WeightsStore[6][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_586;WeightsStore[6][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_587;WeightsStore[6][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_588;WeightsStore[6][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_589;WeightsStore[6][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_590;WeightsStore[6][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_591;WeightsStore[6][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_592;WeightsStore[6][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_593;WeightsStore[6][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_594;WeightsStore[6][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_595;WeightsStore[6][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_596;WeightsStore[6][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_597;WeightsStore[6][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_598;WeightsStore[6][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_599;WeightsStore[6][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_600;WeightsStore[6][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_601;WeightsStore[6][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_602;WeightsStore[6][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_603;WeightsStore[6][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_604;WeightsStore[6][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_605;WeightsStore[6][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_606;WeightsStore[6][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_607;WeightsStore[6][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_608;WeightsStore[6][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_609;WeightsStore[6][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_610;WeightsStore[6][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_611;WeightsStore[6][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_612;WeightsStore[6][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_613;WeightsStore[6][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_614;WeightsStore[6][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_615;WeightsStore[6][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_616;WeightsStore[6][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_617;WeightsStore[6][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_618;WeightsStore[6][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_619;WeightsStore[6][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_620;WeightsStore[6][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_621;WeightsStore[6][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_622;WeightsStore[6][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_623;WeightsStore[6][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_624;WeightsStore[6][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_625;WeightsStore[6][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_626;WeightsStore[6][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_627;WeightsStore[6][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_628;WeightsStore[6][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_629;WeightsStore[6][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_630;WeightsStore[6][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_631;WeightsStore[6][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_632;WeightsStore[6][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_633;WeightsStore[6][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_634;WeightsStore[6][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_635;WeightsStore[6][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_636;WeightsStore[6][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_637;WeightsStore[6][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_638;WeightsStore[6][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_639;WeightsStore[6][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_640;WeightsStore[6][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_641;WeightsStore[6][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_642;WeightsStore[6][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_643;WeightsStore[6][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_644;WeightsStore[6][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_645;WeightsStore[6][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_646;WeightsStore[6][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_647;WeightsStore[6][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_648;WeightsStore[6][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_649;WeightsStore[6][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_650;WeightsStore[6][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_651;WeightsStore[6][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_652;WeightsStore[6][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_653;WeightsStore[6][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_654;WeightsStore[6][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_655;WeightsStore[6][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_656;WeightsStore[6][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_657;WeightsStore[6][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_658;WeightsStore[6][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_659;WeightsStore[6][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_660;WeightsStore[6][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_661;WeightsStore[6][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_662;WeightsStore[6][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_663;WeightsStore[6][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_664;WeightsStore[6][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_665;WeightsStore[6][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_666;WeightsStore[6][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_667;WeightsStore[6][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_668;WeightsStore[6][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_669;WeightsStore[6][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_670;WeightsStore[6][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_671;WeightsStore[6][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_672;WeightsStore[6][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_673;WeightsStore[6][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_674;WeightsStore[6][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_675;WeightsStore[6][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_676;WeightsStore[6][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_677;WeightsStore[6][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_678;WeightsStore[6][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_679;WeightsStore[6][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_680;WeightsStore[6][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_681;WeightsStore[6][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_682;WeightsStore[6][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_683;WeightsStore[6][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_684;WeightsStore[6][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_685;WeightsStore[6][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_686;WeightsStore[6][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_687;WeightsStore[6][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_688;WeightsStore[6][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_689;WeightsStore[6][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_690;WeightsStore[6][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_691;WeightsStore[6][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_692;WeightsStore[6][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_693;WeightsStore[6][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_694;WeightsStore[6][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_695;WeightsStore[6][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_696;WeightsStore[6][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_697;WeightsStore[6][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_698;WeightsStore[6][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_699;WeightsStore[6][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_700;WeightsStore[6][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_701;WeightsStore[6][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_702;WeightsStore[6][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_703;WeightsStore[6][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_704;WeightsStore[6][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_705;WeightsStore[6][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_706;WeightsStore[6][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_707;WeightsStore[6][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_708;WeightsStore[6][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_709;WeightsStore[6][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_710;WeightsStore[6][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_711;WeightsStore[6][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_712;WeightsStore[6][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_713;WeightsStore[6][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_714;WeightsStore[6][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_715;WeightsStore[6][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_716;WeightsStore[6][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_717;WeightsStore[6][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_718;WeightsStore[6][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_719;WeightsStore[6][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_720;WeightsStore[6][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_721;WeightsStore[6][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_722;WeightsStore[6][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_723;WeightsStore[6][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_724;WeightsStore[6][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_725;WeightsStore[6][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_726;WeightsStore[6][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_727;WeightsStore[6][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_728;WeightsStore[6][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_729;WeightsStore[6][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_730;WeightsStore[6][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_731;WeightsStore[6][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_732;WeightsStore[6][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_733;WeightsStore[6][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_734;WeightsStore[6][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_735;WeightsStore[6][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_736;WeightsStore[6][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_737;WeightsStore[6][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_738;WeightsStore[6][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_739;WeightsStore[6][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_740;WeightsStore[6][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_741;WeightsStore[6][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_742;WeightsStore[6][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_743;WeightsStore[6][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_744;WeightsStore[6][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_745;WeightsStore[6][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_746;WeightsStore[6][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_747;WeightsStore[6][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_748;WeightsStore[6][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_749;WeightsStore[6][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_750;WeightsStore[6][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_751;WeightsStore[6][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_752;WeightsStore[6][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_753;WeightsStore[6][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_754;WeightsStore[6][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_755;WeightsStore[6][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_756;WeightsStore[6][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_757;WeightsStore[6][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_758;WeightsStore[6][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_759;WeightsStore[6][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_760;WeightsStore[6][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_761;WeightsStore[6][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_762;WeightsStore[6][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_763;WeightsStore[6][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_764;WeightsStore[6][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_765;WeightsStore[6][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_766;WeightsStore[6][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_767;WeightsStore[6][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_768;WeightsStore[6][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_769;WeightsStore[6][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_770;WeightsStore[6][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_771;WeightsStore[6][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_772;WeightsStore[6][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_773;WeightsStore[6][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_774;WeightsStore[6][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_775;WeightsStore[6][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_776;WeightsStore[6][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_777;WeightsStore[6][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_778;WeightsStore[6][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_779;WeightsStore[6][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_780;WeightsStore[6][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_781;WeightsStore[6][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_782;WeightsStore[6][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_783;WeightsStore[6][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_6_784;WeightsStore[7][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_0;WeightsStore[7][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_1;WeightsStore[7][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_2;WeightsStore[7][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_3;WeightsStore[7][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_4;WeightsStore[7][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_5;WeightsStore[7][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_6;WeightsStore[7][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_7;WeightsStore[7][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_8;WeightsStore[7][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_9;WeightsStore[7][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_10;WeightsStore[7][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_11;WeightsStore[7][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_12;WeightsStore[7][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_13;WeightsStore[7][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_14;WeightsStore[7][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_15;WeightsStore[7][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_16;WeightsStore[7][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_17;WeightsStore[7][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_18;WeightsStore[7][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_19;WeightsStore[7][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_20;WeightsStore[7][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_21;WeightsStore[7][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_22;WeightsStore[7][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_23;WeightsStore[7][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_24;WeightsStore[7][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_25;WeightsStore[7][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_26;WeightsStore[7][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_27;WeightsStore[7][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_28;WeightsStore[7][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_29;WeightsStore[7][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_30;WeightsStore[7][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_31;WeightsStore[7][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_32;WeightsStore[7][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_33;WeightsStore[7][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_34;WeightsStore[7][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_35;WeightsStore[7][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_36;WeightsStore[7][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_37;WeightsStore[7][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_38;WeightsStore[7][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_39;WeightsStore[7][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_40;WeightsStore[7][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_41;WeightsStore[7][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_42;WeightsStore[7][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_43;WeightsStore[7][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_44;WeightsStore[7][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_45;WeightsStore[7][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_46;WeightsStore[7][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_47;WeightsStore[7][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_48;WeightsStore[7][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_49;WeightsStore[7][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_50;WeightsStore[7][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_51;WeightsStore[7][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_52;WeightsStore[7][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_53;WeightsStore[7][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_54;WeightsStore[7][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_55;WeightsStore[7][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_56;WeightsStore[7][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_57;WeightsStore[7][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_58;WeightsStore[7][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_59;WeightsStore[7][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_60;WeightsStore[7][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_61;WeightsStore[7][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_62;WeightsStore[7][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_63;WeightsStore[7][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_64;WeightsStore[7][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_65;WeightsStore[7][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_66;WeightsStore[7][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_67;WeightsStore[7][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_68;WeightsStore[7][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_69;WeightsStore[7][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_70;WeightsStore[7][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_71;WeightsStore[7][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_72;WeightsStore[7][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_73;WeightsStore[7][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_74;WeightsStore[7][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_75;WeightsStore[7][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_76;WeightsStore[7][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_77;WeightsStore[7][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_78;WeightsStore[7][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_79;WeightsStore[7][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_80;WeightsStore[7][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_81;WeightsStore[7][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_82;WeightsStore[7][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_83;WeightsStore[7][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_84;WeightsStore[7][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_85;WeightsStore[7][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_86;WeightsStore[7][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_87;WeightsStore[7][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_88;WeightsStore[7][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_89;WeightsStore[7][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_90;WeightsStore[7][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_91;WeightsStore[7][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_92;WeightsStore[7][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_93;WeightsStore[7][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_94;WeightsStore[7][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_95;WeightsStore[7][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_96;WeightsStore[7][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_97;WeightsStore[7][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_98;WeightsStore[7][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_99;WeightsStore[7][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_100;WeightsStore[7][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_101;WeightsStore[7][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_102;WeightsStore[7][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_103;WeightsStore[7][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_104;WeightsStore[7][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_105;WeightsStore[7][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_106;WeightsStore[7][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_107;WeightsStore[7][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_108;WeightsStore[7][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_109;WeightsStore[7][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_110;WeightsStore[7][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_111;WeightsStore[7][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_112;WeightsStore[7][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_113;WeightsStore[7][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_114;WeightsStore[7][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_115;WeightsStore[7][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_116;WeightsStore[7][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_117;WeightsStore[7][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_118;WeightsStore[7][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_119;WeightsStore[7][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_120;WeightsStore[7][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_121;WeightsStore[7][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_122;WeightsStore[7][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_123;WeightsStore[7][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_124;WeightsStore[7][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_125;WeightsStore[7][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_126;WeightsStore[7][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_127;WeightsStore[7][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_128;WeightsStore[7][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_129;WeightsStore[7][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_130;WeightsStore[7][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_131;WeightsStore[7][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_132;WeightsStore[7][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_133;WeightsStore[7][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_134;WeightsStore[7][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_135;WeightsStore[7][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_136;WeightsStore[7][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_137;WeightsStore[7][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_138;WeightsStore[7][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_139;WeightsStore[7][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_140;WeightsStore[7][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_141;WeightsStore[7][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_142;WeightsStore[7][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_143;WeightsStore[7][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_144;WeightsStore[7][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_145;WeightsStore[7][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_146;WeightsStore[7][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_147;WeightsStore[7][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_148;WeightsStore[7][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_149;WeightsStore[7][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_150;WeightsStore[7][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_151;WeightsStore[7][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_152;WeightsStore[7][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_153;WeightsStore[7][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_154;WeightsStore[7][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_155;WeightsStore[7][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_156;WeightsStore[7][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_157;WeightsStore[7][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_158;WeightsStore[7][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_159;WeightsStore[7][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_160;WeightsStore[7][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_161;WeightsStore[7][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_162;WeightsStore[7][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_163;WeightsStore[7][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_164;WeightsStore[7][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_165;WeightsStore[7][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_166;WeightsStore[7][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_167;WeightsStore[7][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_168;WeightsStore[7][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_169;WeightsStore[7][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_170;WeightsStore[7][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_171;WeightsStore[7][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_172;WeightsStore[7][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_173;WeightsStore[7][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_174;WeightsStore[7][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_175;WeightsStore[7][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_176;WeightsStore[7][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_177;WeightsStore[7][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_178;WeightsStore[7][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_179;WeightsStore[7][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_180;WeightsStore[7][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_181;WeightsStore[7][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_182;WeightsStore[7][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_183;WeightsStore[7][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_184;WeightsStore[7][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_185;WeightsStore[7][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_186;WeightsStore[7][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_187;WeightsStore[7][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_188;WeightsStore[7][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_189;WeightsStore[7][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_190;WeightsStore[7][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_191;WeightsStore[7][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_192;WeightsStore[7][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_193;WeightsStore[7][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_194;WeightsStore[7][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_195;WeightsStore[7][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_196;WeightsStore[7][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_197;WeightsStore[7][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_198;WeightsStore[7][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_199;WeightsStore[7][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_200;WeightsStore[7][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_201;WeightsStore[7][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_202;WeightsStore[7][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_203;WeightsStore[7][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_204;WeightsStore[7][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_205;WeightsStore[7][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_206;WeightsStore[7][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_207;WeightsStore[7][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_208;WeightsStore[7][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_209;WeightsStore[7][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_210;WeightsStore[7][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_211;WeightsStore[7][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_212;WeightsStore[7][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_213;WeightsStore[7][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_214;WeightsStore[7][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_215;WeightsStore[7][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_216;WeightsStore[7][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_217;WeightsStore[7][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_218;WeightsStore[7][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_219;WeightsStore[7][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_220;WeightsStore[7][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_221;WeightsStore[7][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_222;WeightsStore[7][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_223;WeightsStore[7][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_224;WeightsStore[7][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_225;WeightsStore[7][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_226;WeightsStore[7][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_227;WeightsStore[7][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_228;WeightsStore[7][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_229;WeightsStore[7][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_230;WeightsStore[7][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_231;WeightsStore[7][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_232;WeightsStore[7][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_233;WeightsStore[7][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_234;WeightsStore[7][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_235;WeightsStore[7][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_236;WeightsStore[7][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_237;WeightsStore[7][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_238;WeightsStore[7][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_239;WeightsStore[7][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_240;WeightsStore[7][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_241;WeightsStore[7][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_242;WeightsStore[7][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_243;WeightsStore[7][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_244;WeightsStore[7][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_245;WeightsStore[7][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_246;WeightsStore[7][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_247;WeightsStore[7][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_248;WeightsStore[7][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_249;WeightsStore[7][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_250;WeightsStore[7][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_251;WeightsStore[7][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_252;WeightsStore[7][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_253;WeightsStore[7][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_254;WeightsStore[7][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_255;WeightsStore[7][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_256;WeightsStore[7][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_257;WeightsStore[7][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_258;WeightsStore[7][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_259;WeightsStore[7][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_260;WeightsStore[7][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_261;WeightsStore[7][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_262;WeightsStore[7][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_263;WeightsStore[7][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_264;WeightsStore[7][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_265;WeightsStore[7][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_266;WeightsStore[7][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_267;WeightsStore[7][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_268;WeightsStore[7][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_269;WeightsStore[7][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_270;WeightsStore[7][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_271;WeightsStore[7][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_272;WeightsStore[7][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_273;WeightsStore[7][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_274;WeightsStore[7][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_275;WeightsStore[7][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_276;WeightsStore[7][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_277;WeightsStore[7][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_278;WeightsStore[7][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_279;WeightsStore[7][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_280;WeightsStore[7][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_281;WeightsStore[7][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_282;WeightsStore[7][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_283;WeightsStore[7][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_284;WeightsStore[7][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_285;WeightsStore[7][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_286;WeightsStore[7][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_287;WeightsStore[7][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_288;WeightsStore[7][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_289;WeightsStore[7][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_290;WeightsStore[7][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_291;WeightsStore[7][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_292;WeightsStore[7][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_293;WeightsStore[7][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_294;WeightsStore[7][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_295;WeightsStore[7][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_296;WeightsStore[7][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_297;WeightsStore[7][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_298;WeightsStore[7][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_299;WeightsStore[7][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_300;WeightsStore[7][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_301;WeightsStore[7][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_302;WeightsStore[7][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_303;WeightsStore[7][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_304;WeightsStore[7][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_305;WeightsStore[7][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_306;WeightsStore[7][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_307;WeightsStore[7][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_308;WeightsStore[7][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_309;WeightsStore[7][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_310;WeightsStore[7][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_311;WeightsStore[7][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_312;WeightsStore[7][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_313;WeightsStore[7][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_314;WeightsStore[7][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_315;WeightsStore[7][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_316;WeightsStore[7][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_317;WeightsStore[7][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_318;WeightsStore[7][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_319;WeightsStore[7][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_320;WeightsStore[7][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_321;WeightsStore[7][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_322;WeightsStore[7][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_323;WeightsStore[7][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_324;WeightsStore[7][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_325;WeightsStore[7][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_326;WeightsStore[7][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_327;WeightsStore[7][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_328;WeightsStore[7][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_329;WeightsStore[7][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_330;WeightsStore[7][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_331;WeightsStore[7][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_332;WeightsStore[7][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_333;WeightsStore[7][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_334;WeightsStore[7][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_335;WeightsStore[7][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_336;WeightsStore[7][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_337;WeightsStore[7][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_338;WeightsStore[7][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_339;WeightsStore[7][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_340;WeightsStore[7][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_341;WeightsStore[7][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_342;WeightsStore[7][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_343;WeightsStore[7][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_344;WeightsStore[7][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_345;WeightsStore[7][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_346;WeightsStore[7][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_347;WeightsStore[7][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_348;WeightsStore[7][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_349;WeightsStore[7][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_350;WeightsStore[7][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_351;WeightsStore[7][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_352;WeightsStore[7][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_353;WeightsStore[7][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_354;WeightsStore[7][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_355;WeightsStore[7][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_356;WeightsStore[7][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_357;WeightsStore[7][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_358;WeightsStore[7][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_359;WeightsStore[7][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_360;WeightsStore[7][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_361;WeightsStore[7][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_362;WeightsStore[7][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_363;WeightsStore[7][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_364;WeightsStore[7][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_365;WeightsStore[7][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_366;WeightsStore[7][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_367;WeightsStore[7][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_368;WeightsStore[7][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_369;WeightsStore[7][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_370;WeightsStore[7][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_371;WeightsStore[7][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_372;WeightsStore[7][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_373;WeightsStore[7][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_374;WeightsStore[7][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_375;WeightsStore[7][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_376;WeightsStore[7][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_377;WeightsStore[7][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_378;WeightsStore[7][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_379;WeightsStore[7][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_380;WeightsStore[7][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_381;WeightsStore[7][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_382;WeightsStore[7][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_383;WeightsStore[7][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_384;WeightsStore[7][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_385;WeightsStore[7][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_386;WeightsStore[7][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_387;WeightsStore[7][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_388;WeightsStore[7][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_389;WeightsStore[7][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_390;WeightsStore[7][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_391;WeightsStore[7][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_392;WeightsStore[7][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_393;WeightsStore[7][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_394;WeightsStore[7][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_395;WeightsStore[7][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_396;WeightsStore[7][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_397;WeightsStore[7][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_398;WeightsStore[7][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_399;WeightsStore[7][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_400;WeightsStore[7][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_401;WeightsStore[7][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_402;WeightsStore[7][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_403;WeightsStore[7][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_404;WeightsStore[7][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_405;WeightsStore[7][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_406;WeightsStore[7][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_407;WeightsStore[7][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_408;WeightsStore[7][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_409;WeightsStore[7][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_410;WeightsStore[7][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_411;WeightsStore[7][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_412;WeightsStore[7][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_413;WeightsStore[7][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_414;WeightsStore[7][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_415;WeightsStore[7][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_416;WeightsStore[7][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_417;WeightsStore[7][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_418;WeightsStore[7][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_419;WeightsStore[7][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_420;WeightsStore[7][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_421;WeightsStore[7][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_422;WeightsStore[7][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_423;WeightsStore[7][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_424;WeightsStore[7][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_425;WeightsStore[7][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_426;WeightsStore[7][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_427;WeightsStore[7][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_428;WeightsStore[7][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_429;WeightsStore[7][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_430;WeightsStore[7][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_431;WeightsStore[7][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_432;WeightsStore[7][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_433;WeightsStore[7][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_434;WeightsStore[7][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_435;WeightsStore[7][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_436;WeightsStore[7][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_437;WeightsStore[7][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_438;WeightsStore[7][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_439;WeightsStore[7][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_440;WeightsStore[7][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_441;WeightsStore[7][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_442;WeightsStore[7][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_443;WeightsStore[7][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_444;WeightsStore[7][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_445;WeightsStore[7][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_446;WeightsStore[7][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_447;WeightsStore[7][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_448;WeightsStore[7][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_449;WeightsStore[7][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_450;WeightsStore[7][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_451;WeightsStore[7][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_452;WeightsStore[7][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_453;WeightsStore[7][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_454;WeightsStore[7][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_455;WeightsStore[7][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_456;WeightsStore[7][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_457;WeightsStore[7][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_458;WeightsStore[7][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_459;WeightsStore[7][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_460;WeightsStore[7][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_461;WeightsStore[7][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_462;WeightsStore[7][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_463;WeightsStore[7][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_464;WeightsStore[7][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_465;WeightsStore[7][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_466;WeightsStore[7][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_467;WeightsStore[7][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_468;WeightsStore[7][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_469;WeightsStore[7][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_470;WeightsStore[7][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_471;WeightsStore[7][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_472;WeightsStore[7][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_473;WeightsStore[7][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_474;WeightsStore[7][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_475;WeightsStore[7][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_476;WeightsStore[7][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_477;WeightsStore[7][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_478;WeightsStore[7][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_479;WeightsStore[7][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_480;WeightsStore[7][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_481;WeightsStore[7][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_482;WeightsStore[7][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_483;WeightsStore[7][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_484;WeightsStore[7][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_485;WeightsStore[7][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_486;WeightsStore[7][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_487;WeightsStore[7][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_488;WeightsStore[7][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_489;WeightsStore[7][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_490;WeightsStore[7][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_491;WeightsStore[7][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_492;WeightsStore[7][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_493;WeightsStore[7][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_494;WeightsStore[7][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_495;WeightsStore[7][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_496;WeightsStore[7][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_497;WeightsStore[7][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_498;WeightsStore[7][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_499;WeightsStore[7][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_500;WeightsStore[7][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_501;WeightsStore[7][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_502;WeightsStore[7][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_503;WeightsStore[7][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_504;WeightsStore[7][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_505;WeightsStore[7][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_506;WeightsStore[7][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_507;WeightsStore[7][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_508;WeightsStore[7][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_509;WeightsStore[7][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_510;WeightsStore[7][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_511;WeightsStore[7][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_512;WeightsStore[7][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_513;WeightsStore[7][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_514;WeightsStore[7][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_515;WeightsStore[7][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_516;WeightsStore[7][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_517;WeightsStore[7][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_518;WeightsStore[7][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_519;WeightsStore[7][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_520;WeightsStore[7][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_521;WeightsStore[7][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_522;WeightsStore[7][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_523;WeightsStore[7][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_524;WeightsStore[7][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_525;WeightsStore[7][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_526;WeightsStore[7][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_527;WeightsStore[7][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_528;WeightsStore[7][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_529;WeightsStore[7][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_530;WeightsStore[7][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_531;WeightsStore[7][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_532;WeightsStore[7][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_533;WeightsStore[7][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_534;WeightsStore[7][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_535;WeightsStore[7][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_536;WeightsStore[7][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_537;WeightsStore[7][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_538;WeightsStore[7][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_539;WeightsStore[7][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_540;WeightsStore[7][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_541;WeightsStore[7][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_542;WeightsStore[7][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_543;WeightsStore[7][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_544;WeightsStore[7][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_545;WeightsStore[7][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_546;WeightsStore[7][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_547;WeightsStore[7][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_548;WeightsStore[7][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_549;WeightsStore[7][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_550;WeightsStore[7][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_551;WeightsStore[7][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_552;WeightsStore[7][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_553;WeightsStore[7][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_554;WeightsStore[7][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_555;WeightsStore[7][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_556;WeightsStore[7][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_557;WeightsStore[7][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_558;WeightsStore[7][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_559;WeightsStore[7][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_560;WeightsStore[7][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_561;WeightsStore[7][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_562;WeightsStore[7][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_563;WeightsStore[7][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_564;WeightsStore[7][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_565;WeightsStore[7][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_566;WeightsStore[7][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_567;WeightsStore[7][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_568;WeightsStore[7][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_569;WeightsStore[7][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_570;WeightsStore[7][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_571;WeightsStore[7][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_572;WeightsStore[7][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_573;WeightsStore[7][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_574;WeightsStore[7][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_575;WeightsStore[7][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_576;WeightsStore[7][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_577;WeightsStore[7][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_578;WeightsStore[7][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_579;WeightsStore[7][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_580;WeightsStore[7][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_581;WeightsStore[7][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_582;WeightsStore[7][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_583;WeightsStore[7][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_584;WeightsStore[7][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_585;WeightsStore[7][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_586;WeightsStore[7][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_587;WeightsStore[7][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_588;WeightsStore[7][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_589;WeightsStore[7][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_590;WeightsStore[7][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_591;WeightsStore[7][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_592;WeightsStore[7][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_593;WeightsStore[7][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_594;WeightsStore[7][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_595;WeightsStore[7][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_596;WeightsStore[7][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_597;WeightsStore[7][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_598;WeightsStore[7][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_599;WeightsStore[7][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_600;WeightsStore[7][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_601;WeightsStore[7][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_602;WeightsStore[7][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_603;WeightsStore[7][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_604;WeightsStore[7][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_605;WeightsStore[7][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_606;WeightsStore[7][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_607;WeightsStore[7][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_608;WeightsStore[7][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_609;WeightsStore[7][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_610;WeightsStore[7][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_611;WeightsStore[7][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_612;WeightsStore[7][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_613;WeightsStore[7][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_614;WeightsStore[7][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_615;WeightsStore[7][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_616;WeightsStore[7][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_617;WeightsStore[7][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_618;WeightsStore[7][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_619;WeightsStore[7][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_620;WeightsStore[7][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_621;WeightsStore[7][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_622;WeightsStore[7][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_623;WeightsStore[7][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_624;WeightsStore[7][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_625;WeightsStore[7][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_626;WeightsStore[7][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_627;WeightsStore[7][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_628;WeightsStore[7][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_629;WeightsStore[7][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_630;WeightsStore[7][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_631;WeightsStore[7][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_632;WeightsStore[7][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_633;WeightsStore[7][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_634;WeightsStore[7][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_635;WeightsStore[7][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_636;WeightsStore[7][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_637;WeightsStore[7][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_638;WeightsStore[7][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_639;WeightsStore[7][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_640;WeightsStore[7][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_641;WeightsStore[7][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_642;WeightsStore[7][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_643;WeightsStore[7][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_644;WeightsStore[7][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_645;WeightsStore[7][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_646;WeightsStore[7][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_647;WeightsStore[7][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_648;WeightsStore[7][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_649;WeightsStore[7][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_650;WeightsStore[7][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_651;WeightsStore[7][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_652;WeightsStore[7][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_653;WeightsStore[7][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_654;WeightsStore[7][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_655;WeightsStore[7][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_656;WeightsStore[7][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_657;WeightsStore[7][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_658;WeightsStore[7][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_659;WeightsStore[7][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_660;WeightsStore[7][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_661;WeightsStore[7][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_662;WeightsStore[7][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_663;WeightsStore[7][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_664;WeightsStore[7][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_665;WeightsStore[7][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_666;WeightsStore[7][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_667;WeightsStore[7][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_668;WeightsStore[7][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_669;WeightsStore[7][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_670;WeightsStore[7][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_671;WeightsStore[7][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_672;WeightsStore[7][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_673;WeightsStore[7][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_674;WeightsStore[7][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_675;WeightsStore[7][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_676;WeightsStore[7][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_677;WeightsStore[7][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_678;WeightsStore[7][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_679;WeightsStore[7][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_680;WeightsStore[7][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_681;WeightsStore[7][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_682;WeightsStore[7][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_683;WeightsStore[7][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_684;WeightsStore[7][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_685;WeightsStore[7][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_686;WeightsStore[7][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_687;WeightsStore[7][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_688;WeightsStore[7][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_689;WeightsStore[7][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_690;WeightsStore[7][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_691;WeightsStore[7][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_692;WeightsStore[7][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_693;WeightsStore[7][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_694;WeightsStore[7][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_695;WeightsStore[7][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_696;WeightsStore[7][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_697;WeightsStore[7][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_698;WeightsStore[7][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_699;WeightsStore[7][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_700;WeightsStore[7][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_701;WeightsStore[7][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_702;WeightsStore[7][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_703;WeightsStore[7][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_704;WeightsStore[7][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_705;WeightsStore[7][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_706;WeightsStore[7][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_707;WeightsStore[7][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_708;WeightsStore[7][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_709;WeightsStore[7][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_710;WeightsStore[7][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_711;WeightsStore[7][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_712;WeightsStore[7][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_713;WeightsStore[7][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_714;WeightsStore[7][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_715;WeightsStore[7][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_716;WeightsStore[7][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_717;WeightsStore[7][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_718;WeightsStore[7][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_719;WeightsStore[7][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_720;WeightsStore[7][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_721;WeightsStore[7][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_722;WeightsStore[7][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_723;WeightsStore[7][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_724;WeightsStore[7][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_725;WeightsStore[7][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_726;WeightsStore[7][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_727;WeightsStore[7][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_728;WeightsStore[7][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_729;WeightsStore[7][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_730;WeightsStore[7][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_731;WeightsStore[7][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_732;WeightsStore[7][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_733;WeightsStore[7][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_734;WeightsStore[7][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_735;WeightsStore[7][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_736;WeightsStore[7][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_737;WeightsStore[7][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_738;WeightsStore[7][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_739;WeightsStore[7][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_740;WeightsStore[7][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_741;WeightsStore[7][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_742;WeightsStore[7][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_743;WeightsStore[7][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_744;WeightsStore[7][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_745;WeightsStore[7][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_746;WeightsStore[7][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_747;WeightsStore[7][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_748;WeightsStore[7][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_749;WeightsStore[7][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_750;WeightsStore[7][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_751;WeightsStore[7][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_752;WeightsStore[7][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_753;WeightsStore[7][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_754;WeightsStore[7][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_755;WeightsStore[7][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_756;WeightsStore[7][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_757;WeightsStore[7][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_758;WeightsStore[7][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_759;WeightsStore[7][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_760;WeightsStore[7][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_761;WeightsStore[7][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_762;WeightsStore[7][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_763;WeightsStore[7][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_764;WeightsStore[7][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_765;WeightsStore[7][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_766;WeightsStore[7][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_767;WeightsStore[7][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_768;WeightsStore[7][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_769;WeightsStore[7][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_770;WeightsStore[7][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_771;WeightsStore[7][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_772;WeightsStore[7][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_773;WeightsStore[7][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_774;WeightsStore[7][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_775;WeightsStore[7][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_776;WeightsStore[7][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_777;WeightsStore[7][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_778;WeightsStore[7][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_779;WeightsStore[7][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_780;WeightsStore[7][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_781;WeightsStore[7][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_782;WeightsStore[7][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_783;WeightsStore[7][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_7_784;WeightsStore[8][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_0;WeightsStore[8][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_1;WeightsStore[8][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_2;WeightsStore[8][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_3;WeightsStore[8][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_4;WeightsStore[8][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_5;WeightsStore[8][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_6;WeightsStore[8][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_7;WeightsStore[8][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_8;WeightsStore[8][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_9;WeightsStore[8][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_10;WeightsStore[8][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_11;WeightsStore[8][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_12;WeightsStore[8][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_13;WeightsStore[8][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_14;WeightsStore[8][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_15;WeightsStore[8][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_16;WeightsStore[8][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_17;WeightsStore[8][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_18;WeightsStore[8][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_19;WeightsStore[8][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_20;WeightsStore[8][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_21;WeightsStore[8][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_22;WeightsStore[8][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_23;WeightsStore[8][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_24;WeightsStore[8][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_25;WeightsStore[8][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_26;WeightsStore[8][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_27;WeightsStore[8][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_28;WeightsStore[8][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_29;WeightsStore[8][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_30;WeightsStore[8][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_31;WeightsStore[8][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_32;WeightsStore[8][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_33;WeightsStore[8][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_34;WeightsStore[8][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_35;WeightsStore[8][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_36;WeightsStore[8][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_37;WeightsStore[8][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_38;WeightsStore[8][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_39;WeightsStore[8][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_40;WeightsStore[8][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_41;WeightsStore[8][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_42;WeightsStore[8][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_43;WeightsStore[8][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_44;WeightsStore[8][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_45;WeightsStore[8][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_46;WeightsStore[8][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_47;WeightsStore[8][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_48;WeightsStore[8][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_49;WeightsStore[8][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_50;WeightsStore[8][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_51;WeightsStore[8][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_52;WeightsStore[8][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_53;WeightsStore[8][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_54;WeightsStore[8][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_55;WeightsStore[8][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_56;WeightsStore[8][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_57;WeightsStore[8][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_58;WeightsStore[8][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_59;WeightsStore[8][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_60;WeightsStore[8][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_61;WeightsStore[8][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_62;WeightsStore[8][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_63;WeightsStore[8][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_64;WeightsStore[8][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_65;WeightsStore[8][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_66;WeightsStore[8][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_67;WeightsStore[8][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_68;WeightsStore[8][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_69;WeightsStore[8][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_70;WeightsStore[8][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_71;WeightsStore[8][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_72;WeightsStore[8][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_73;WeightsStore[8][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_74;WeightsStore[8][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_75;WeightsStore[8][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_76;WeightsStore[8][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_77;WeightsStore[8][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_78;WeightsStore[8][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_79;WeightsStore[8][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_80;WeightsStore[8][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_81;WeightsStore[8][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_82;WeightsStore[8][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_83;WeightsStore[8][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_84;WeightsStore[8][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_85;WeightsStore[8][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_86;WeightsStore[8][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_87;WeightsStore[8][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_88;WeightsStore[8][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_89;WeightsStore[8][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_90;WeightsStore[8][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_91;WeightsStore[8][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_92;WeightsStore[8][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_93;WeightsStore[8][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_94;WeightsStore[8][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_95;WeightsStore[8][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_96;WeightsStore[8][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_97;WeightsStore[8][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_98;WeightsStore[8][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_99;WeightsStore[8][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_100;WeightsStore[8][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_101;WeightsStore[8][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_102;WeightsStore[8][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_103;WeightsStore[8][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_104;WeightsStore[8][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_105;WeightsStore[8][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_106;WeightsStore[8][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_107;WeightsStore[8][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_108;WeightsStore[8][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_109;WeightsStore[8][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_110;WeightsStore[8][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_111;WeightsStore[8][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_112;WeightsStore[8][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_113;WeightsStore[8][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_114;WeightsStore[8][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_115;WeightsStore[8][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_116;WeightsStore[8][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_117;WeightsStore[8][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_118;WeightsStore[8][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_119;WeightsStore[8][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_120;WeightsStore[8][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_121;WeightsStore[8][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_122;WeightsStore[8][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_123;WeightsStore[8][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_124;WeightsStore[8][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_125;WeightsStore[8][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_126;WeightsStore[8][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_127;WeightsStore[8][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_128;WeightsStore[8][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_129;WeightsStore[8][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_130;WeightsStore[8][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_131;WeightsStore[8][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_132;WeightsStore[8][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_133;WeightsStore[8][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_134;WeightsStore[8][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_135;WeightsStore[8][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_136;WeightsStore[8][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_137;WeightsStore[8][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_138;WeightsStore[8][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_139;WeightsStore[8][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_140;WeightsStore[8][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_141;WeightsStore[8][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_142;WeightsStore[8][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_143;WeightsStore[8][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_144;WeightsStore[8][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_145;WeightsStore[8][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_146;WeightsStore[8][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_147;WeightsStore[8][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_148;WeightsStore[8][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_149;WeightsStore[8][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_150;WeightsStore[8][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_151;WeightsStore[8][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_152;WeightsStore[8][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_153;WeightsStore[8][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_154;WeightsStore[8][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_155;WeightsStore[8][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_156;WeightsStore[8][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_157;WeightsStore[8][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_158;WeightsStore[8][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_159;WeightsStore[8][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_160;WeightsStore[8][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_161;WeightsStore[8][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_162;WeightsStore[8][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_163;WeightsStore[8][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_164;WeightsStore[8][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_165;WeightsStore[8][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_166;WeightsStore[8][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_167;WeightsStore[8][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_168;WeightsStore[8][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_169;WeightsStore[8][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_170;WeightsStore[8][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_171;WeightsStore[8][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_172;WeightsStore[8][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_173;WeightsStore[8][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_174;WeightsStore[8][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_175;WeightsStore[8][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_176;WeightsStore[8][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_177;WeightsStore[8][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_178;WeightsStore[8][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_179;WeightsStore[8][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_180;WeightsStore[8][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_181;WeightsStore[8][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_182;WeightsStore[8][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_183;WeightsStore[8][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_184;WeightsStore[8][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_185;WeightsStore[8][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_186;WeightsStore[8][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_187;WeightsStore[8][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_188;WeightsStore[8][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_189;WeightsStore[8][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_190;WeightsStore[8][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_191;WeightsStore[8][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_192;WeightsStore[8][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_193;WeightsStore[8][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_194;WeightsStore[8][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_195;WeightsStore[8][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_196;WeightsStore[8][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_197;WeightsStore[8][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_198;WeightsStore[8][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_199;WeightsStore[8][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_200;WeightsStore[8][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_201;WeightsStore[8][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_202;WeightsStore[8][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_203;WeightsStore[8][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_204;WeightsStore[8][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_205;WeightsStore[8][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_206;WeightsStore[8][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_207;WeightsStore[8][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_208;WeightsStore[8][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_209;WeightsStore[8][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_210;WeightsStore[8][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_211;WeightsStore[8][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_212;WeightsStore[8][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_213;WeightsStore[8][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_214;WeightsStore[8][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_215;WeightsStore[8][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_216;WeightsStore[8][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_217;WeightsStore[8][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_218;WeightsStore[8][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_219;WeightsStore[8][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_220;WeightsStore[8][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_221;WeightsStore[8][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_222;WeightsStore[8][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_223;WeightsStore[8][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_224;WeightsStore[8][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_225;WeightsStore[8][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_226;WeightsStore[8][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_227;WeightsStore[8][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_228;WeightsStore[8][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_229;WeightsStore[8][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_230;WeightsStore[8][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_231;WeightsStore[8][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_232;WeightsStore[8][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_233;WeightsStore[8][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_234;WeightsStore[8][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_235;WeightsStore[8][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_236;WeightsStore[8][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_237;WeightsStore[8][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_238;WeightsStore[8][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_239;WeightsStore[8][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_240;WeightsStore[8][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_241;WeightsStore[8][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_242;WeightsStore[8][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_243;WeightsStore[8][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_244;WeightsStore[8][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_245;WeightsStore[8][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_246;WeightsStore[8][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_247;WeightsStore[8][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_248;WeightsStore[8][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_249;WeightsStore[8][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_250;WeightsStore[8][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_251;WeightsStore[8][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_252;WeightsStore[8][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_253;WeightsStore[8][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_254;WeightsStore[8][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_255;WeightsStore[8][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_256;WeightsStore[8][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_257;WeightsStore[8][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_258;WeightsStore[8][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_259;WeightsStore[8][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_260;WeightsStore[8][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_261;WeightsStore[8][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_262;WeightsStore[8][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_263;WeightsStore[8][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_264;WeightsStore[8][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_265;WeightsStore[8][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_266;WeightsStore[8][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_267;WeightsStore[8][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_268;WeightsStore[8][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_269;WeightsStore[8][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_270;WeightsStore[8][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_271;WeightsStore[8][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_272;WeightsStore[8][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_273;WeightsStore[8][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_274;WeightsStore[8][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_275;WeightsStore[8][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_276;WeightsStore[8][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_277;WeightsStore[8][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_278;WeightsStore[8][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_279;WeightsStore[8][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_280;WeightsStore[8][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_281;WeightsStore[8][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_282;WeightsStore[8][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_283;WeightsStore[8][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_284;WeightsStore[8][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_285;WeightsStore[8][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_286;WeightsStore[8][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_287;WeightsStore[8][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_288;WeightsStore[8][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_289;WeightsStore[8][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_290;WeightsStore[8][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_291;WeightsStore[8][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_292;WeightsStore[8][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_293;WeightsStore[8][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_294;WeightsStore[8][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_295;WeightsStore[8][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_296;WeightsStore[8][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_297;WeightsStore[8][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_298;WeightsStore[8][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_299;WeightsStore[8][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_300;WeightsStore[8][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_301;WeightsStore[8][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_302;WeightsStore[8][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_303;WeightsStore[8][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_304;WeightsStore[8][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_305;WeightsStore[8][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_306;WeightsStore[8][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_307;WeightsStore[8][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_308;WeightsStore[8][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_309;WeightsStore[8][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_310;WeightsStore[8][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_311;WeightsStore[8][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_312;WeightsStore[8][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_313;WeightsStore[8][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_314;WeightsStore[8][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_315;WeightsStore[8][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_316;WeightsStore[8][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_317;WeightsStore[8][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_318;WeightsStore[8][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_319;WeightsStore[8][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_320;WeightsStore[8][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_321;WeightsStore[8][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_322;WeightsStore[8][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_323;WeightsStore[8][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_324;WeightsStore[8][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_325;WeightsStore[8][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_326;WeightsStore[8][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_327;WeightsStore[8][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_328;WeightsStore[8][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_329;WeightsStore[8][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_330;WeightsStore[8][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_331;WeightsStore[8][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_332;WeightsStore[8][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_333;WeightsStore[8][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_334;WeightsStore[8][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_335;WeightsStore[8][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_336;WeightsStore[8][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_337;WeightsStore[8][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_338;WeightsStore[8][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_339;WeightsStore[8][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_340;WeightsStore[8][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_341;WeightsStore[8][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_342;WeightsStore[8][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_343;WeightsStore[8][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_344;WeightsStore[8][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_345;WeightsStore[8][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_346;WeightsStore[8][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_347;WeightsStore[8][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_348;WeightsStore[8][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_349;WeightsStore[8][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_350;WeightsStore[8][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_351;WeightsStore[8][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_352;WeightsStore[8][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_353;WeightsStore[8][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_354;WeightsStore[8][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_355;WeightsStore[8][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_356;WeightsStore[8][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_357;WeightsStore[8][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_358;WeightsStore[8][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_359;WeightsStore[8][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_360;WeightsStore[8][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_361;WeightsStore[8][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_362;WeightsStore[8][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_363;WeightsStore[8][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_364;WeightsStore[8][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_365;WeightsStore[8][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_366;WeightsStore[8][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_367;WeightsStore[8][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_368;WeightsStore[8][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_369;WeightsStore[8][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_370;WeightsStore[8][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_371;WeightsStore[8][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_372;WeightsStore[8][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_373;WeightsStore[8][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_374;WeightsStore[8][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_375;WeightsStore[8][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_376;WeightsStore[8][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_377;WeightsStore[8][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_378;WeightsStore[8][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_379;WeightsStore[8][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_380;WeightsStore[8][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_381;WeightsStore[8][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_382;WeightsStore[8][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_383;WeightsStore[8][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_384;WeightsStore[8][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_385;WeightsStore[8][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_386;WeightsStore[8][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_387;WeightsStore[8][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_388;WeightsStore[8][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_389;WeightsStore[8][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_390;WeightsStore[8][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_391;WeightsStore[8][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_392;WeightsStore[8][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_393;WeightsStore[8][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_394;WeightsStore[8][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_395;WeightsStore[8][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_396;WeightsStore[8][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_397;WeightsStore[8][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_398;WeightsStore[8][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_399;WeightsStore[8][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_400;WeightsStore[8][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_401;WeightsStore[8][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_402;WeightsStore[8][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_403;WeightsStore[8][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_404;WeightsStore[8][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_405;WeightsStore[8][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_406;WeightsStore[8][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_407;WeightsStore[8][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_408;WeightsStore[8][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_409;WeightsStore[8][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_410;WeightsStore[8][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_411;WeightsStore[8][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_412;WeightsStore[8][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_413;WeightsStore[8][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_414;WeightsStore[8][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_415;WeightsStore[8][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_416;WeightsStore[8][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_417;WeightsStore[8][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_418;WeightsStore[8][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_419;WeightsStore[8][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_420;WeightsStore[8][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_421;WeightsStore[8][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_422;WeightsStore[8][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_423;WeightsStore[8][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_424;WeightsStore[8][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_425;WeightsStore[8][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_426;WeightsStore[8][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_427;WeightsStore[8][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_428;WeightsStore[8][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_429;WeightsStore[8][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_430;WeightsStore[8][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_431;WeightsStore[8][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_432;WeightsStore[8][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_433;WeightsStore[8][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_434;WeightsStore[8][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_435;WeightsStore[8][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_436;WeightsStore[8][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_437;WeightsStore[8][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_438;WeightsStore[8][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_439;WeightsStore[8][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_440;WeightsStore[8][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_441;WeightsStore[8][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_442;WeightsStore[8][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_443;WeightsStore[8][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_444;WeightsStore[8][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_445;WeightsStore[8][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_446;WeightsStore[8][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_447;WeightsStore[8][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_448;WeightsStore[8][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_449;WeightsStore[8][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_450;WeightsStore[8][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_451;WeightsStore[8][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_452;WeightsStore[8][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_453;WeightsStore[8][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_454;WeightsStore[8][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_455;WeightsStore[8][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_456;WeightsStore[8][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_457;WeightsStore[8][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_458;WeightsStore[8][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_459;WeightsStore[8][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_460;WeightsStore[8][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_461;WeightsStore[8][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_462;WeightsStore[8][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_463;WeightsStore[8][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_464;WeightsStore[8][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_465;WeightsStore[8][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_466;WeightsStore[8][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_467;WeightsStore[8][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_468;WeightsStore[8][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_469;WeightsStore[8][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_470;WeightsStore[8][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_471;WeightsStore[8][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_472;WeightsStore[8][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_473;WeightsStore[8][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_474;WeightsStore[8][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_475;WeightsStore[8][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_476;WeightsStore[8][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_477;WeightsStore[8][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_478;WeightsStore[8][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_479;WeightsStore[8][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_480;WeightsStore[8][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_481;WeightsStore[8][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_482;WeightsStore[8][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_483;WeightsStore[8][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_484;WeightsStore[8][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_485;WeightsStore[8][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_486;WeightsStore[8][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_487;WeightsStore[8][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_488;WeightsStore[8][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_489;WeightsStore[8][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_490;WeightsStore[8][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_491;WeightsStore[8][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_492;WeightsStore[8][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_493;WeightsStore[8][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_494;WeightsStore[8][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_495;WeightsStore[8][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_496;WeightsStore[8][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_497;WeightsStore[8][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_498;WeightsStore[8][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_499;WeightsStore[8][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_500;WeightsStore[8][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_501;WeightsStore[8][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_502;WeightsStore[8][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_503;WeightsStore[8][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_504;WeightsStore[8][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_505;WeightsStore[8][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_506;WeightsStore[8][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_507;WeightsStore[8][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_508;WeightsStore[8][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_509;WeightsStore[8][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_510;WeightsStore[8][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_511;WeightsStore[8][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_512;WeightsStore[8][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_513;WeightsStore[8][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_514;WeightsStore[8][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_515;WeightsStore[8][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_516;WeightsStore[8][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_517;WeightsStore[8][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_518;WeightsStore[8][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_519;WeightsStore[8][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_520;WeightsStore[8][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_521;WeightsStore[8][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_522;WeightsStore[8][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_523;WeightsStore[8][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_524;WeightsStore[8][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_525;WeightsStore[8][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_526;WeightsStore[8][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_527;WeightsStore[8][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_528;WeightsStore[8][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_529;WeightsStore[8][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_530;WeightsStore[8][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_531;WeightsStore[8][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_532;WeightsStore[8][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_533;WeightsStore[8][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_534;WeightsStore[8][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_535;WeightsStore[8][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_536;WeightsStore[8][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_537;WeightsStore[8][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_538;WeightsStore[8][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_539;WeightsStore[8][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_540;WeightsStore[8][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_541;WeightsStore[8][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_542;WeightsStore[8][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_543;WeightsStore[8][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_544;WeightsStore[8][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_545;WeightsStore[8][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_546;WeightsStore[8][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_547;WeightsStore[8][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_548;WeightsStore[8][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_549;WeightsStore[8][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_550;WeightsStore[8][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_551;WeightsStore[8][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_552;WeightsStore[8][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_553;WeightsStore[8][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_554;WeightsStore[8][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_555;WeightsStore[8][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_556;WeightsStore[8][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_557;WeightsStore[8][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_558;WeightsStore[8][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_559;WeightsStore[8][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_560;WeightsStore[8][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_561;WeightsStore[8][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_562;WeightsStore[8][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_563;WeightsStore[8][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_564;WeightsStore[8][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_565;WeightsStore[8][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_566;WeightsStore[8][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_567;WeightsStore[8][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_568;WeightsStore[8][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_569;WeightsStore[8][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_570;WeightsStore[8][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_571;WeightsStore[8][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_572;WeightsStore[8][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_573;WeightsStore[8][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_574;WeightsStore[8][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_575;WeightsStore[8][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_576;WeightsStore[8][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_577;WeightsStore[8][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_578;WeightsStore[8][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_579;WeightsStore[8][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_580;WeightsStore[8][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_581;WeightsStore[8][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_582;WeightsStore[8][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_583;WeightsStore[8][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_584;WeightsStore[8][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_585;WeightsStore[8][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_586;WeightsStore[8][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_587;WeightsStore[8][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_588;WeightsStore[8][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_589;WeightsStore[8][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_590;WeightsStore[8][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_591;WeightsStore[8][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_592;WeightsStore[8][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_593;WeightsStore[8][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_594;WeightsStore[8][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_595;WeightsStore[8][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_596;WeightsStore[8][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_597;WeightsStore[8][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_598;WeightsStore[8][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_599;WeightsStore[8][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_600;WeightsStore[8][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_601;WeightsStore[8][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_602;WeightsStore[8][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_603;WeightsStore[8][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_604;WeightsStore[8][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_605;WeightsStore[8][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_606;WeightsStore[8][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_607;WeightsStore[8][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_608;WeightsStore[8][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_609;WeightsStore[8][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_610;WeightsStore[8][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_611;WeightsStore[8][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_612;WeightsStore[8][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_613;WeightsStore[8][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_614;WeightsStore[8][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_615;WeightsStore[8][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_616;WeightsStore[8][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_617;WeightsStore[8][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_618;WeightsStore[8][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_619;WeightsStore[8][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_620;WeightsStore[8][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_621;WeightsStore[8][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_622;WeightsStore[8][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_623;WeightsStore[8][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_624;WeightsStore[8][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_625;WeightsStore[8][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_626;WeightsStore[8][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_627;WeightsStore[8][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_628;WeightsStore[8][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_629;WeightsStore[8][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_630;WeightsStore[8][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_631;WeightsStore[8][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_632;WeightsStore[8][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_633;WeightsStore[8][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_634;WeightsStore[8][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_635;WeightsStore[8][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_636;WeightsStore[8][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_637;WeightsStore[8][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_638;WeightsStore[8][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_639;WeightsStore[8][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_640;WeightsStore[8][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_641;WeightsStore[8][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_642;WeightsStore[8][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_643;WeightsStore[8][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_644;WeightsStore[8][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_645;WeightsStore[8][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_646;WeightsStore[8][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_647;WeightsStore[8][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_648;WeightsStore[8][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_649;WeightsStore[8][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_650;WeightsStore[8][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_651;WeightsStore[8][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_652;WeightsStore[8][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_653;WeightsStore[8][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_654;WeightsStore[8][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_655;WeightsStore[8][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_656;WeightsStore[8][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_657;WeightsStore[8][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_658;WeightsStore[8][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_659;WeightsStore[8][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_660;WeightsStore[8][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_661;WeightsStore[8][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_662;WeightsStore[8][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_663;WeightsStore[8][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_664;WeightsStore[8][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_665;WeightsStore[8][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_666;WeightsStore[8][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_667;WeightsStore[8][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_668;WeightsStore[8][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_669;WeightsStore[8][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_670;WeightsStore[8][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_671;WeightsStore[8][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_672;WeightsStore[8][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_673;WeightsStore[8][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_674;WeightsStore[8][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_675;WeightsStore[8][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_676;WeightsStore[8][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_677;WeightsStore[8][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_678;WeightsStore[8][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_679;WeightsStore[8][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_680;WeightsStore[8][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_681;WeightsStore[8][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_682;WeightsStore[8][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_683;WeightsStore[8][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_684;WeightsStore[8][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_685;WeightsStore[8][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_686;WeightsStore[8][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_687;WeightsStore[8][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_688;WeightsStore[8][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_689;WeightsStore[8][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_690;WeightsStore[8][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_691;WeightsStore[8][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_692;WeightsStore[8][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_693;WeightsStore[8][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_694;WeightsStore[8][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_695;WeightsStore[8][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_696;WeightsStore[8][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_697;WeightsStore[8][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_698;WeightsStore[8][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_699;WeightsStore[8][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_700;WeightsStore[8][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_701;WeightsStore[8][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_702;WeightsStore[8][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_703;WeightsStore[8][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_704;WeightsStore[8][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_705;WeightsStore[8][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_706;WeightsStore[8][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_707;WeightsStore[8][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_708;WeightsStore[8][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_709;WeightsStore[8][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_710;WeightsStore[8][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_711;WeightsStore[8][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_712;WeightsStore[8][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_713;WeightsStore[8][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_714;WeightsStore[8][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_715;WeightsStore[8][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_716;WeightsStore[8][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_717;WeightsStore[8][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_718;WeightsStore[8][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_719;WeightsStore[8][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_720;WeightsStore[8][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_721;WeightsStore[8][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_722;WeightsStore[8][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_723;WeightsStore[8][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_724;WeightsStore[8][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_725;WeightsStore[8][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_726;WeightsStore[8][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_727;WeightsStore[8][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_728;WeightsStore[8][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_729;WeightsStore[8][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_730;WeightsStore[8][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_731;WeightsStore[8][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_732;WeightsStore[8][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_733;WeightsStore[8][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_734;WeightsStore[8][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_735;WeightsStore[8][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_736;WeightsStore[8][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_737;WeightsStore[8][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_738;WeightsStore[8][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_739;WeightsStore[8][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_740;WeightsStore[8][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_741;WeightsStore[8][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_742;WeightsStore[8][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_743;WeightsStore[8][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_744;WeightsStore[8][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_745;WeightsStore[8][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_746;WeightsStore[8][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_747;WeightsStore[8][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_748;WeightsStore[8][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_749;WeightsStore[8][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_750;WeightsStore[8][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_751;WeightsStore[8][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_752;WeightsStore[8][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_753;WeightsStore[8][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_754;WeightsStore[8][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_755;WeightsStore[8][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_756;WeightsStore[8][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_757;WeightsStore[8][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_758;WeightsStore[8][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_759;WeightsStore[8][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_760;WeightsStore[8][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_761;WeightsStore[8][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_762;WeightsStore[8][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_763;WeightsStore[8][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_764;WeightsStore[8][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_765;WeightsStore[8][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_766;WeightsStore[8][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_767;WeightsStore[8][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_768;WeightsStore[8][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_769;WeightsStore[8][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_770;WeightsStore[8][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_771;WeightsStore[8][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_772;WeightsStore[8][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_773;WeightsStore[8][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_774;WeightsStore[8][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_775;WeightsStore[8][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_776;WeightsStore[8][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_777;WeightsStore[8][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_778;WeightsStore[8][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_779;WeightsStore[8][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_780;WeightsStore[8][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_781;WeightsStore[8][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_782;WeightsStore[8][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_783;WeightsStore[8][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_8_784;WeightsStore[9][0*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_0;WeightsStore[9][1*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_1;WeightsStore[9][2*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_2;WeightsStore[9][3*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_3;WeightsStore[9][4*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_4;WeightsStore[9][5*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_5;WeightsStore[9][6*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_6;WeightsStore[9][7*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_7;WeightsStore[9][8*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_8;WeightsStore[9][9*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_9;WeightsStore[9][10*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_10;WeightsStore[9][11*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_11;WeightsStore[9][12*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_12;WeightsStore[9][13*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_13;WeightsStore[9][14*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_14;WeightsStore[9][15*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_15;WeightsStore[9][16*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_16;WeightsStore[9][17*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_17;WeightsStore[9][18*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_18;WeightsStore[9][19*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_19;WeightsStore[9][20*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_20;WeightsStore[9][21*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_21;WeightsStore[9][22*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_22;WeightsStore[9][23*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_23;WeightsStore[9][24*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_24;WeightsStore[9][25*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_25;WeightsStore[9][26*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_26;WeightsStore[9][27*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_27;WeightsStore[9][28*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_28;WeightsStore[9][29*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_29;WeightsStore[9][30*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_30;WeightsStore[9][31*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_31;WeightsStore[9][32*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_32;WeightsStore[9][33*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_33;WeightsStore[9][34*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_34;WeightsStore[9][35*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_35;WeightsStore[9][36*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_36;WeightsStore[9][37*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_37;WeightsStore[9][38*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_38;WeightsStore[9][39*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_39;WeightsStore[9][40*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_40;WeightsStore[9][41*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_41;WeightsStore[9][42*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_42;WeightsStore[9][43*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_43;WeightsStore[9][44*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_44;WeightsStore[9][45*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_45;WeightsStore[9][46*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_46;WeightsStore[9][47*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_47;WeightsStore[9][48*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_48;WeightsStore[9][49*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_49;WeightsStore[9][50*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_50;WeightsStore[9][51*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_51;WeightsStore[9][52*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_52;WeightsStore[9][53*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_53;WeightsStore[9][54*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_54;WeightsStore[9][55*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_55;WeightsStore[9][56*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_56;WeightsStore[9][57*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_57;WeightsStore[9][58*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_58;WeightsStore[9][59*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_59;WeightsStore[9][60*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_60;WeightsStore[9][61*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_61;WeightsStore[9][62*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_62;WeightsStore[9][63*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_63;WeightsStore[9][64*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_64;WeightsStore[9][65*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_65;WeightsStore[9][66*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_66;WeightsStore[9][67*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_67;WeightsStore[9][68*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_68;WeightsStore[9][69*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_69;WeightsStore[9][70*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_70;WeightsStore[9][71*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_71;WeightsStore[9][72*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_72;WeightsStore[9][73*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_73;WeightsStore[9][74*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_74;WeightsStore[9][75*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_75;WeightsStore[9][76*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_76;WeightsStore[9][77*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_77;WeightsStore[9][78*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_78;WeightsStore[9][79*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_79;WeightsStore[9][80*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_80;WeightsStore[9][81*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_81;WeightsStore[9][82*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_82;WeightsStore[9][83*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_83;WeightsStore[9][84*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_84;WeightsStore[9][85*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_85;WeightsStore[9][86*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_86;WeightsStore[9][87*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_87;WeightsStore[9][88*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_88;WeightsStore[9][89*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_89;WeightsStore[9][90*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_90;WeightsStore[9][91*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_91;WeightsStore[9][92*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_92;WeightsStore[9][93*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_93;WeightsStore[9][94*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_94;WeightsStore[9][95*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_95;WeightsStore[9][96*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_96;WeightsStore[9][97*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_97;WeightsStore[9][98*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_98;WeightsStore[9][99*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_99;WeightsStore[9][100*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_100;WeightsStore[9][101*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_101;WeightsStore[9][102*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_102;WeightsStore[9][103*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_103;WeightsStore[9][104*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_104;WeightsStore[9][105*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_105;WeightsStore[9][106*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_106;WeightsStore[9][107*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_107;WeightsStore[9][108*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_108;WeightsStore[9][109*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_109;WeightsStore[9][110*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_110;WeightsStore[9][111*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_111;WeightsStore[9][112*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_112;WeightsStore[9][113*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_113;WeightsStore[9][114*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_114;WeightsStore[9][115*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_115;WeightsStore[9][116*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_116;WeightsStore[9][117*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_117;WeightsStore[9][118*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_118;WeightsStore[9][119*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_119;WeightsStore[9][120*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_120;WeightsStore[9][121*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_121;WeightsStore[9][122*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_122;WeightsStore[9][123*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_123;WeightsStore[9][124*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_124;WeightsStore[9][125*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_125;WeightsStore[9][126*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_126;WeightsStore[9][127*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_127;WeightsStore[9][128*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_128;WeightsStore[9][129*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_129;WeightsStore[9][130*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_130;WeightsStore[9][131*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_131;WeightsStore[9][132*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_132;WeightsStore[9][133*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_133;WeightsStore[9][134*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_134;WeightsStore[9][135*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_135;WeightsStore[9][136*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_136;WeightsStore[9][137*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_137;WeightsStore[9][138*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_138;WeightsStore[9][139*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_139;WeightsStore[9][140*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_140;WeightsStore[9][141*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_141;WeightsStore[9][142*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_142;WeightsStore[9][143*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_143;WeightsStore[9][144*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_144;WeightsStore[9][145*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_145;WeightsStore[9][146*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_146;WeightsStore[9][147*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_147;WeightsStore[9][148*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_148;WeightsStore[9][149*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_149;WeightsStore[9][150*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_150;WeightsStore[9][151*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_151;WeightsStore[9][152*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_152;WeightsStore[9][153*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_153;WeightsStore[9][154*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_154;WeightsStore[9][155*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_155;WeightsStore[9][156*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_156;WeightsStore[9][157*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_157;WeightsStore[9][158*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_158;WeightsStore[9][159*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_159;WeightsStore[9][160*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_160;WeightsStore[9][161*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_161;WeightsStore[9][162*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_162;WeightsStore[9][163*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_163;WeightsStore[9][164*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_164;WeightsStore[9][165*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_165;WeightsStore[9][166*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_166;WeightsStore[9][167*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_167;WeightsStore[9][168*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_168;WeightsStore[9][169*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_169;WeightsStore[9][170*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_170;WeightsStore[9][171*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_171;WeightsStore[9][172*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_172;WeightsStore[9][173*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_173;WeightsStore[9][174*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_174;WeightsStore[9][175*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_175;WeightsStore[9][176*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_176;WeightsStore[9][177*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_177;WeightsStore[9][178*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_178;WeightsStore[9][179*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_179;WeightsStore[9][180*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_180;WeightsStore[9][181*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_181;WeightsStore[9][182*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_182;WeightsStore[9][183*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_183;WeightsStore[9][184*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_184;WeightsStore[9][185*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_185;WeightsStore[9][186*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_186;WeightsStore[9][187*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_187;WeightsStore[9][188*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_188;WeightsStore[9][189*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_189;WeightsStore[9][190*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_190;WeightsStore[9][191*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_191;WeightsStore[9][192*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_192;WeightsStore[9][193*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_193;WeightsStore[9][194*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_194;WeightsStore[9][195*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_195;WeightsStore[9][196*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_196;WeightsStore[9][197*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_197;WeightsStore[9][198*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_198;WeightsStore[9][199*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_199;WeightsStore[9][200*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_200;WeightsStore[9][201*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_201;WeightsStore[9][202*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_202;WeightsStore[9][203*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_203;WeightsStore[9][204*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_204;WeightsStore[9][205*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_205;WeightsStore[9][206*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_206;WeightsStore[9][207*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_207;WeightsStore[9][208*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_208;WeightsStore[9][209*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_209;WeightsStore[9][210*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_210;WeightsStore[9][211*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_211;WeightsStore[9][212*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_212;WeightsStore[9][213*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_213;WeightsStore[9][214*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_214;WeightsStore[9][215*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_215;WeightsStore[9][216*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_216;WeightsStore[9][217*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_217;WeightsStore[9][218*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_218;WeightsStore[9][219*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_219;WeightsStore[9][220*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_220;WeightsStore[9][221*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_221;WeightsStore[9][222*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_222;WeightsStore[9][223*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_223;WeightsStore[9][224*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_224;WeightsStore[9][225*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_225;WeightsStore[9][226*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_226;WeightsStore[9][227*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_227;WeightsStore[9][228*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_228;WeightsStore[9][229*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_229;WeightsStore[9][230*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_230;WeightsStore[9][231*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_231;WeightsStore[9][232*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_232;WeightsStore[9][233*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_233;WeightsStore[9][234*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_234;WeightsStore[9][235*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_235;WeightsStore[9][236*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_236;WeightsStore[9][237*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_237;WeightsStore[9][238*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_238;WeightsStore[9][239*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_239;WeightsStore[9][240*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_240;WeightsStore[9][241*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_241;WeightsStore[9][242*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_242;WeightsStore[9][243*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_243;WeightsStore[9][244*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_244;WeightsStore[9][245*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_245;WeightsStore[9][246*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_246;WeightsStore[9][247*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_247;WeightsStore[9][248*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_248;WeightsStore[9][249*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_249;WeightsStore[9][250*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_250;WeightsStore[9][251*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_251;WeightsStore[9][252*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_252;WeightsStore[9][253*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_253;WeightsStore[9][254*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_254;WeightsStore[9][255*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_255;WeightsStore[9][256*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_256;WeightsStore[9][257*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_257;WeightsStore[9][258*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_258;WeightsStore[9][259*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_259;WeightsStore[9][260*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_260;WeightsStore[9][261*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_261;WeightsStore[9][262*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_262;WeightsStore[9][263*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_263;WeightsStore[9][264*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_264;WeightsStore[9][265*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_265;WeightsStore[9][266*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_266;WeightsStore[9][267*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_267;WeightsStore[9][268*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_268;WeightsStore[9][269*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_269;WeightsStore[9][270*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_270;WeightsStore[9][271*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_271;WeightsStore[9][272*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_272;WeightsStore[9][273*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_273;WeightsStore[9][274*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_274;WeightsStore[9][275*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_275;WeightsStore[9][276*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_276;WeightsStore[9][277*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_277;WeightsStore[9][278*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_278;WeightsStore[9][279*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_279;WeightsStore[9][280*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_280;WeightsStore[9][281*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_281;WeightsStore[9][282*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_282;WeightsStore[9][283*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_283;WeightsStore[9][284*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_284;WeightsStore[9][285*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_285;WeightsStore[9][286*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_286;WeightsStore[9][287*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_287;WeightsStore[9][288*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_288;WeightsStore[9][289*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_289;WeightsStore[9][290*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_290;WeightsStore[9][291*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_291;WeightsStore[9][292*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_292;WeightsStore[9][293*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_293;WeightsStore[9][294*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_294;WeightsStore[9][295*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_295;WeightsStore[9][296*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_296;WeightsStore[9][297*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_297;WeightsStore[9][298*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_298;WeightsStore[9][299*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_299;WeightsStore[9][300*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_300;WeightsStore[9][301*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_301;WeightsStore[9][302*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_302;WeightsStore[9][303*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_303;WeightsStore[9][304*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_304;WeightsStore[9][305*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_305;WeightsStore[9][306*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_306;WeightsStore[9][307*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_307;WeightsStore[9][308*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_308;WeightsStore[9][309*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_309;WeightsStore[9][310*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_310;WeightsStore[9][311*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_311;WeightsStore[9][312*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_312;WeightsStore[9][313*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_313;WeightsStore[9][314*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_314;WeightsStore[9][315*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_315;WeightsStore[9][316*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_316;WeightsStore[9][317*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_317;WeightsStore[9][318*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_318;WeightsStore[9][319*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_319;WeightsStore[9][320*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_320;WeightsStore[9][321*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_321;WeightsStore[9][322*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_322;WeightsStore[9][323*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_323;WeightsStore[9][324*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_324;WeightsStore[9][325*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_325;WeightsStore[9][326*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_326;WeightsStore[9][327*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_327;WeightsStore[9][328*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_328;WeightsStore[9][329*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_329;WeightsStore[9][330*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_330;WeightsStore[9][331*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_331;WeightsStore[9][332*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_332;WeightsStore[9][333*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_333;WeightsStore[9][334*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_334;WeightsStore[9][335*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_335;WeightsStore[9][336*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_336;WeightsStore[9][337*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_337;WeightsStore[9][338*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_338;WeightsStore[9][339*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_339;WeightsStore[9][340*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_340;WeightsStore[9][341*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_341;WeightsStore[9][342*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_342;WeightsStore[9][343*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_343;WeightsStore[9][344*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_344;WeightsStore[9][345*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_345;WeightsStore[9][346*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_346;WeightsStore[9][347*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_347;WeightsStore[9][348*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_348;WeightsStore[9][349*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_349;WeightsStore[9][350*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_350;WeightsStore[9][351*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_351;WeightsStore[9][352*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_352;WeightsStore[9][353*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_353;WeightsStore[9][354*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_354;WeightsStore[9][355*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_355;WeightsStore[9][356*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_356;WeightsStore[9][357*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_357;WeightsStore[9][358*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_358;WeightsStore[9][359*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_359;WeightsStore[9][360*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_360;WeightsStore[9][361*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_361;WeightsStore[9][362*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_362;WeightsStore[9][363*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_363;WeightsStore[9][364*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_364;WeightsStore[9][365*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_365;WeightsStore[9][366*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_366;WeightsStore[9][367*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_367;WeightsStore[9][368*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_368;WeightsStore[9][369*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_369;WeightsStore[9][370*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_370;WeightsStore[9][371*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_371;WeightsStore[9][372*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_372;WeightsStore[9][373*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_373;WeightsStore[9][374*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_374;WeightsStore[9][375*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_375;WeightsStore[9][376*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_376;WeightsStore[9][377*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_377;WeightsStore[9][378*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_378;WeightsStore[9][379*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_379;WeightsStore[9][380*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_380;WeightsStore[9][381*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_381;WeightsStore[9][382*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_382;WeightsStore[9][383*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_383;WeightsStore[9][384*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_384;WeightsStore[9][385*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_385;WeightsStore[9][386*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_386;WeightsStore[9][387*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_387;WeightsStore[9][388*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_388;WeightsStore[9][389*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_389;WeightsStore[9][390*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_390;WeightsStore[9][391*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_391;WeightsStore[9][392*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_392;WeightsStore[9][393*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_393;WeightsStore[9][394*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_394;WeightsStore[9][395*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_395;WeightsStore[9][396*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_396;WeightsStore[9][397*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_397;WeightsStore[9][398*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_398;WeightsStore[9][399*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_399;WeightsStore[9][400*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_400;WeightsStore[9][401*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_401;WeightsStore[9][402*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_402;WeightsStore[9][403*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_403;WeightsStore[9][404*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_404;WeightsStore[9][405*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_405;WeightsStore[9][406*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_406;WeightsStore[9][407*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_407;WeightsStore[9][408*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_408;WeightsStore[9][409*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_409;WeightsStore[9][410*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_410;WeightsStore[9][411*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_411;WeightsStore[9][412*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_412;WeightsStore[9][413*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_413;WeightsStore[9][414*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_414;WeightsStore[9][415*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_415;WeightsStore[9][416*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_416;WeightsStore[9][417*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_417;WeightsStore[9][418*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_418;WeightsStore[9][419*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_419;WeightsStore[9][420*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_420;WeightsStore[9][421*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_421;WeightsStore[9][422*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_422;WeightsStore[9][423*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_423;WeightsStore[9][424*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_424;WeightsStore[9][425*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_425;WeightsStore[9][426*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_426;WeightsStore[9][427*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_427;WeightsStore[9][428*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_428;WeightsStore[9][429*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_429;WeightsStore[9][430*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_430;WeightsStore[9][431*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_431;WeightsStore[9][432*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_432;WeightsStore[9][433*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_433;WeightsStore[9][434*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_434;WeightsStore[9][435*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_435;WeightsStore[9][436*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_436;WeightsStore[9][437*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_437;WeightsStore[9][438*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_438;WeightsStore[9][439*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_439;WeightsStore[9][440*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_440;WeightsStore[9][441*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_441;WeightsStore[9][442*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_442;WeightsStore[9][443*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_443;WeightsStore[9][444*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_444;WeightsStore[9][445*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_445;WeightsStore[9][446*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_446;WeightsStore[9][447*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_447;WeightsStore[9][448*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_448;WeightsStore[9][449*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_449;WeightsStore[9][450*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_450;WeightsStore[9][451*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_451;WeightsStore[9][452*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_452;WeightsStore[9][453*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_453;WeightsStore[9][454*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_454;WeightsStore[9][455*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_455;WeightsStore[9][456*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_456;WeightsStore[9][457*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_457;WeightsStore[9][458*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_458;WeightsStore[9][459*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_459;WeightsStore[9][460*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_460;WeightsStore[9][461*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_461;WeightsStore[9][462*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_462;WeightsStore[9][463*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_463;WeightsStore[9][464*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_464;WeightsStore[9][465*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_465;WeightsStore[9][466*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_466;WeightsStore[9][467*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_467;WeightsStore[9][468*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_468;WeightsStore[9][469*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_469;WeightsStore[9][470*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_470;WeightsStore[9][471*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_471;WeightsStore[9][472*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_472;WeightsStore[9][473*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_473;WeightsStore[9][474*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_474;WeightsStore[9][475*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_475;WeightsStore[9][476*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_476;WeightsStore[9][477*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_477;WeightsStore[9][478*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_478;WeightsStore[9][479*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_479;WeightsStore[9][480*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_480;WeightsStore[9][481*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_481;WeightsStore[9][482*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_482;WeightsStore[9][483*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_483;WeightsStore[9][484*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_484;WeightsStore[9][485*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_485;WeightsStore[9][486*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_486;WeightsStore[9][487*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_487;WeightsStore[9][488*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_488;WeightsStore[9][489*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_489;WeightsStore[9][490*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_490;WeightsStore[9][491*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_491;WeightsStore[9][492*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_492;WeightsStore[9][493*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_493;WeightsStore[9][494*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_494;WeightsStore[9][495*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_495;WeightsStore[9][496*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_496;WeightsStore[9][497*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_497;WeightsStore[9][498*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_498;WeightsStore[9][499*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_499;WeightsStore[9][500*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_500;WeightsStore[9][501*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_501;WeightsStore[9][502*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_502;WeightsStore[9][503*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_503;WeightsStore[9][504*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_504;WeightsStore[9][505*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_505;WeightsStore[9][506*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_506;WeightsStore[9][507*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_507;WeightsStore[9][508*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_508;WeightsStore[9][509*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_509;WeightsStore[9][510*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_510;WeightsStore[9][511*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_511;WeightsStore[9][512*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_512;WeightsStore[9][513*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_513;WeightsStore[9][514*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_514;WeightsStore[9][515*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_515;WeightsStore[9][516*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_516;WeightsStore[9][517*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_517;WeightsStore[9][518*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_518;WeightsStore[9][519*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_519;WeightsStore[9][520*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_520;WeightsStore[9][521*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_521;WeightsStore[9][522*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_522;WeightsStore[9][523*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_523;WeightsStore[9][524*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_524;WeightsStore[9][525*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_525;WeightsStore[9][526*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_526;WeightsStore[9][527*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_527;WeightsStore[9][528*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_528;WeightsStore[9][529*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_529;WeightsStore[9][530*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_530;WeightsStore[9][531*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_531;WeightsStore[9][532*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_532;WeightsStore[9][533*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_533;WeightsStore[9][534*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_534;WeightsStore[9][535*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_535;WeightsStore[9][536*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_536;WeightsStore[9][537*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_537;WeightsStore[9][538*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_538;WeightsStore[9][539*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_539;WeightsStore[9][540*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_540;WeightsStore[9][541*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_541;WeightsStore[9][542*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_542;WeightsStore[9][543*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_543;WeightsStore[9][544*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_544;WeightsStore[9][545*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_545;WeightsStore[9][546*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_546;WeightsStore[9][547*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_547;WeightsStore[9][548*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_548;WeightsStore[9][549*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_549;WeightsStore[9][550*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_550;WeightsStore[9][551*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_551;WeightsStore[9][552*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_552;WeightsStore[9][553*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_553;WeightsStore[9][554*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_554;WeightsStore[9][555*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_555;WeightsStore[9][556*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_556;WeightsStore[9][557*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_557;WeightsStore[9][558*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_558;WeightsStore[9][559*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_559;WeightsStore[9][560*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_560;WeightsStore[9][561*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_561;WeightsStore[9][562*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_562;WeightsStore[9][563*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_563;WeightsStore[9][564*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_564;WeightsStore[9][565*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_565;WeightsStore[9][566*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_566;WeightsStore[9][567*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_567;WeightsStore[9][568*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_568;WeightsStore[9][569*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_569;WeightsStore[9][570*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_570;WeightsStore[9][571*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_571;WeightsStore[9][572*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_572;WeightsStore[9][573*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_573;WeightsStore[9][574*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_574;WeightsStore[9][575*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_575;WeightsStore[9][576*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_576;WeightsStore[9][577*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_577;WeightsStore[9][578*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_578;WeightsStore[9][579*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_579;WeightsStore[9][580*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_580;WeightsStore[9][581*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_581;WeightsStore[9][582*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_582;WeightsStore[9][583*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_583;WeightsStore[9][584*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_584;WeightsStore[9][585*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_585;WeightsStore[9][586*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_586;WeightsStore[9][587*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_587;WeightsStore[9][588*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_588;WeightsStore[9][589*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_589;WeightsStore[9][590*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_590;WeightsStore[9][591*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_591;WeightsStore[9][592*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_592;WeightsStore[9][593*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_593;WeightsStore[9][594*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_594;WeightsStore[9][595*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_595;WeightsStore[9][596*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_596;WeightsStore[9][597*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_597;WeightsStore[9][598*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_598;WeightsStore[9][599*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_599;WeightsStore[9][600*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_600;WeightsStore[9][601*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_601;WeightsStore[9][602*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_602;WeightsStore[9][603*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_603;WeightsStore[9][604*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_604;WeightsStore[9][605*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_605;WeightsStore[9][606*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_606;WeightsStore[9][607*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_607;WeightsStore[9][608*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_608;WeightsStore[9][609*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_609;WeightsStore[9][610*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_610;WeightsStore[9][611*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_611;WeightsStore[9][612*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_612;WeightsStore[9][613*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_613;WeightsStore[9][614*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_614;WeightsStore[9][615*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_615;WeightsStore[9][616*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_616;WeightsStore[9][617*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_617;WeightsStore[9][618*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_618;WeightsStore[9][619*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_619;WeightsStore[9][620*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_620;WeightsStore[9][621*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_621;WeightsStore[9][622*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_622;WeightsStore[9][623*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_623;WeightsStore[9][624*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_624;WeightsStore[9][625*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_625;WeightsStore[9][626*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_626;WeightsStore[9][627*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_627;WeightsStore[9][628*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_628;WeightsStore[9][629*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_629;WeightsStore[9][630*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_630;WeightsStore[9][631*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_631;WeightsStore[9][632*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_632;WeightsStore[9][633*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_633;WeightsStore[9][634*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_634;WeightsStore[9][635*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_635;WeightsStore[9][636*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_636;WeightsStore[9][637*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_637;WeightsStore[9][638*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_638;WeightsStore[9][639*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_639;WeightsStore[9][640*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_640;WeightsStore[9][641*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_641;WeightsStore[9][642*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_642;WeightsStore[9][643*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_643;WeightsStore[9][644*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_644;WeightsStore[9][645*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_645;WeightsStore[9][646*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_646;WeightsStore[9][647*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_647;WeightsStore[9][648*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_648;WeightsStore[9][649*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_649;WeightsStore[9][650*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_650;WeightsStore[9][651*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_651;WeightsStore[9][652*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_652;WeightsStore[9][653*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_653;WeightsStore[9][654*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_654;WeightsStore[9][655*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_655;WeightsStore[9][656*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_656;WeightsStore[9][657*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_657;WeightsStore[9][658*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_658;WeightsStore[9][659*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_659;WeightsStore[9][660*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_660;WeightsStore[9][661*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_661;WeightsStore[9][662*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_662;WeightsStore[9][663*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_663;WeightsStore[9][664*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_664;WeightsStore[9][665*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_665;WeightsStore[9][666*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_666;WeightsStore[9][667*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_667;WeightsStore[9][668*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_668;WeightsStore[9][669*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_669;WeightsStore[9][670*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_670;WeightsStore[9][671*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_671;WeightsStore[9][672*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_672;WeightsStore[9][673*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_673;WeightsStore[9][674*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_674;WeightsStore[9][675*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_675;WeightsStore[9][676*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_676;WeightsStore[9][677*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_677;WeightsStore[9][678*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_678;WeightsStore[9][679*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_679;WeightsStore[9][680*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_680;WeightsStore[9][681*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_681;WeightsStore[9][682*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_682;WeightsStore[9][683*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_683;WeightsStore[9][684*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_684;WeightsStore[9][685*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_685;WeightsStore[9][686*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_686;WeightsStore[9][687*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_687;WeightsStore[9][688*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_688;WeightsStore[9][689*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_689;WeightsStore[9][690*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_690;WeightsStore[9][691*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_691;WeightsStore[9][692*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_692;WeightsStore[9][693*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_693;WeightsStore[9][694*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_694;WeightsStore[9][695*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_695;WeightsStore[9][696*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_696;WeightsStore[9][697*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_697;WeightsStore[9][698*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_698;WeightsStore[9][699*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_699;WeightsStore[9][700*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_700;WeightsStore[9][701*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_701;WeightsStore[9][702*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_702;WeightsStore[9][703*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_703;WeightsStore[9][704*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_704;WeightsStore[9][705*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_705;WeightsStore[9][706*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_706;WeightsStore[9][707*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_707;WeightsStore[9][708*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_708;WeightsStore[9][709*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_709;WeightsStore[9][710*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_710;WeightsStore[9][711*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_711;WeightsStore[9][712*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_712;WeightsStore[9][713*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_713;WeightsStore[9][714*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_714;WeightsStore[9][715*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_715;WeightsStore[9][716*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_716;WeightsStore[9][717*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_717;WeightsStore[9][718*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_718;WeightsStore[9][719*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_719;WeightsStore[9][720*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_720;WeightsStore[9][721*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_721;WeightsStore[9][722*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_722;WeightsStore[9][723*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_723;WeightsStore[9][724*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_724;WeightsStore[9][725*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_725;WeightsStore[9][726*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_726;WeightsStore[9][727*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_727;WeightsStore[9][728*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_728;WeightsStore[9][729*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_729;WeightsStore[9][730*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_730;WeightsStore[9][731*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_731;WeightsStore[9][732*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_732;WeightsStore[9][733*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_733;WeightsStore[9][734*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_734;WeightsStore[9][735*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_735;WeightsStore[9][736*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_736;WeightsStore[9][737*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_737;WeightsStore[9][738*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_738;WeightsStore[9][739*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_739;WeightsStore[9][740*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_740;WeightsStore[9][741*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_741;WeightsStore[9][742*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_742;WeightsStore[9][743*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_743;WeightsStore[9][744*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_744;WeightsStore[9][745*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_745;WeightsStore[9][746*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_746;WeightsStore[9][747*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_747;WeightsStore[9][748*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_748;WeightsStore[9][749*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_749;WeightsStore[9][750*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_750;WeightsStore[9][751*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_751;WeightsStore[9][752*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_752;WeightsStore[9][753*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_753;WeightsStore[9][754*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_754;WeightsStore[9][755*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_755;WeightsStore[9][756*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_756;WeightsStore[9][757*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_757;WeightsStore[9][758*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_758;WeightsStore[9][759*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_759;WeightsStore[9][760*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_760;WeightsStore[9][761*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_761;WeightsStore[9][762*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_762;WeightsStore[9][763*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_763;WeightsStore[9][764*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_764;WeightsStore[9][765*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_765;WeightsStore[9][766*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_766;WeightsStore[9][767*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_767;WeightsStore[9][768*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_768;WeightsStore[9][769*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_769;WeightsStore[9][770*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_770;WeightsStore[9][771*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_771;WeightsStore[9][772*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_772;WeightsStore[9][773*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_773;WeightsStore[9][774*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_774;WeightsStore[9][775*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_775;WeightsStore[9][776*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_776;WeightsStore[9][777*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_777;WeightsStore[9][778*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_778;WeightsStore[9][779*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_779;WeightsStore[9][780*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_780;WeightsStore[9][781*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_781;WeightsStore[9][782*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_782;WeightsStore[9][783*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_783;WeightsStore[9][784*WEIGHT_SIZE+:WEIGHT_SIZE]<=Wgt_9_784;
		flag <= 1;
	end
	else if(flag == 1) begin
		switchCounter <= 0;
        internalReset <= 1'b0;
		flag <= 0;
	end
	else begin
		PixelInput <= 0;
		if(switchCounter < 300) begin
			switchCounter <= switchCounter + 1;
		end
		else if(switchCounter==320) begin
			ready <= 1'b1;
			/*
			$display("9: %d %b.%b %h", switchCounter, value[259:252],value[251:234],value[259:234]);
			$display("8: %d %b.%b %h", switchCounter, value[233:226],value[225:208],value[233:208]);
			$display("7: %d %b.%b %h", switchCounter, value[207:200],value[199:182],value[207:182]);
			$display("6: %d %b.%b %h", switchCounter, value[181:174],value[173:156],value[181:156]);
			$display("5: %d %b.%b %h", switchCounter, value[155:148],value[147:130],value[155:130]);
			$display("4: %d %b.%b %h", switchCounter, value[129:122],value[121:104],value[129:104]);
			$display("3: %d %b.%b %h", switchCounter, value[103:96],value[95:78],value[103:78]);
			$display("2: %d %b.%b %h", switchCounter, value[77:70],value[69:52],value[77:52]);
			$display("1: %d %b.%b %h", switchCounter, value[51:44],value[43:26],value[51:26]);
			$display("0: %d %b.%b %h", switchCounter, value[25:18],value[17:0],value[25:0]);
			*/
			switchCounter <= switchCounter + 1;
			//$display("%h", PixelsStore);
		end

	end
end
endmodule
