module VectorMatrixProduct
#(parameter PIXEL_N = 784,
parameter WEIGHT_SIZE = 19,
parameter PIXEL_SIZE = 10)
(
input clk,
input GlobalReset,
input [PIXEL_N*PIXEL_SIZE-1:0] Pixels,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights0,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights1,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights2,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights3,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights4,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights5,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights6,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights7,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights8,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights9,
output [259:0] value
);

reg[9:0] PixelsStore[0:27];
reg[18:0] WeightsStore0[0:27];
reg[18:0] WeightsStore1[0:27];
reg[18:0] WeightsStore2[0:27];
reg[18:0] WeightsStore3[0:27];
reg[18:0] WeightsStore4[0:27];
reg[18:0] WeightsStore5[0:27];
reg[18:0] WeightsStore6[0:27];
reg[18:0] WeightsStore7[0:27];
reg[18:0] WeightsStore8[0:27];
reg[18:0] WeightsStore9[0:27];
reg[31:0] switchCounter;
wire[25:0] vals [0:9];

assign value[25:0] = vals[0];
assign value[51:26] = vals[1];
assign value[77:52] = vals[2];
assign value[103:78] = vals[3];
assign value[129:104] = vals[4];
assign value[155:130] = vals[5];
assign value[181:156] = vals[6];
assign value[207:182] = vals[7];
assign value[233:208] = vals[8];
assign value[259:234] = vals[9];
DotProduct784 DP0(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore0[0]),
	.Weight1(WeightsStore0[1]),
	.Weight2(WeightsStore0[2]),
	.Weight3(WeightsStore0[3]),
	.Weight4(WeightsStore0[4]),
	.Weight5(WeightsStore0[5]),
	.Weight6(WeightsStore0[6]),
	.Weight7(WeightsStore0[7]),
	.Weight8(WeightsStore0[8]),
	.Weight9(WeightsStore0[9]),
	.Weight10(WeightsStore0[10]),
	.Weight11(WeightsStore0[11]),
	.Weight12(WeightsStore0[12]),
	.Weight13(WeightsStore0[13]),
	.Weight14(WeightsStore0[14]),
	.Weight15(WeightsStore0[15]),
	.Weight16(WeightsStore0[16]),
	.Weight17(WeightsStore0[17]),
	.Weight18(WeightsStore0[18]),
	.Weight19(WeightsStore0[19]),
	.Weight20(WeightsStore0[20]),
	.Weight21(WeightsStore0[21]),
	.Weight22(WeightsStore0[22]),
	.Weight23(WeightsStore0[23]),
	.Weight24(WeightsStore0[24]),
	.Weight25(WeightsStore0[25]),
	.Weight26(WeightsStore0[26]),
	.Weight27(WeightsStore0[27]),
	.value(vals[0])
	);
DotProduct784 DP1(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore1[0]),
	.Weight1(WeightsStore1[1]),
	.Weight2(WeightsStore1[2]),
	.Weight3(WeightsStore1[3]),
	.Weight4(WeightsStore1[4]),
	.Weight5(WeightsStore1[5]),
	.Weight6(WeightsStore1[6]),
	.Weight7(WeightsStore1[7]),
	.Weight8(WeightsStore1[8]),
	.Weight9(WeightsStore1[9]),
	.Weight10(WeightsStore1[10]),
	.Weight11(WeightsStore1[11]),
	.Weight12(WeightsStore1[12]),
	.Weight13(WeightsStore1[13]),
	.Weight14(WeightsStore1[14]),
	.Weight15(WeightsStore1[15]),
	.Weight16(WeightsStore1[16]),
	.Weight17(WeightsStore1[17]),
	.Weight18(WeightsStore1[18]),
	.Weight19(WeightsStore1[19]),
	.Weight20(WeightsStore1[20]),
	.Weight21(WeightsStore1[21]),
	.Weight22(WeightsStore1[22]),
	.Weight23(WeightsStore1[23]),
	.Weight24(WeightsStore1[24]),
	.Weight25(WeightsStore1[25]),
	.Weight26(WeightsStore1[26]),
	.Weight27(WeightsStore1[27]),
	.value(vals[1])
	);
DotProduct784 DP2(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore2[0]),
	.Weight1(WeightsStore2[1]),
	.Weight2(WeightsStore2[2]),
	.Weight3(WeightsStore2[3]),
	.Weight4(WeightsStore2[4]),
	.Weight5(WeightsStore2[5]),
	.Weight6(WeightsStore2[6]),
	.Weight7(WeightsStore2[7]),
	.Weight8(WeightsStore2[8]),
	.Weight9(WeightsStore2[9]),
	.Weight10(WeightsStore2[10]),
	.Weight11(WeightsStore2[11]),
	.Weight12(WeightsStore2[12]),
	.Weight13(WeightsStore2[13]),
	.Weight14(WeightsStore2[14]),
	.Weight15(WeightsStore2[15]),
	.Weight16(WeightsStore2[16]),
	.Weight17(WeightsStore2[17]),
	.Weight18(WeightsStore2[18]),
	.Weight19(WeightsStore2[19]),
	.Weight20(WeightsStore2[20]),
	.Weight21(WeightsStore2[21]),
	.Weight22(WeightsStore2[22]),
	.Weight23(WeightsStore2[23]),
	.Weight24(WeightsStore2[24]),
	.Weight25(WeightsStore2[25]),
	.Weight26(WeightsStore2[26]),
	.Weight27(WeightsStore2[27]),
	.value(vals[2])
	);
DotProduct784 DP3(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore3[0]),
	.Weight1(WeightsStore3[1]),
	.Weight2(WeightsStore3[2]),
	.Weight3(WeightsStore3[3]),
	.Weight4(WeightsStore3[4]),
	.Weight5(WeightsStore3[5]),
	.Weight6(WeightsStore3[6]),
	.Weight7(WeightsStore3[7]),
	.Weight8(WeightsStore3[8]),
	.Weight9(WeightsStore3[9]),
	.Weight10(WeightsStore3[10]),
	.Weight11(WeightsStore3[11]),
	.Weight12(WeightsStore3[12]),
	.Weight13(WeightsStore3[13]),
	.Weight14(WeightsStore3[14]),
	.Weight15(WeightsStore3[15]),
	.Weight16(WeightsStore3[16]),
	.Weight17(WeightsStore3[17]),
	.Weight18(WeightsStore3[18]),
	.Weight19(WeightsStore3[19]),
	.Weight20(WeightsStore3[20]),
	.Weight21(WeightsStore3[21]),
	.Weight22(WeightsStore3[22]),
	.Weight23(WeightsStore3[23]),
	.Weight24(WeightsStore3[24]),
	.Weight25(WeightsStore3[25]),
	.Weight26(WeightsStore3[26]),
	.Weight27(WeightsStore3[27]),
	.value(vals[3])
	);
DotProduct784 DP4(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore4[0]),
	.Weight1(WeightsStore4[1]),
	.Weight2(WeightsStore4[2]),
	.Weight3(WeightsStore4[3]),
	.Weight4(WeightsStore4[4]),
	.Weight5(WeightsStore4[5]),
	.Weight6(WeightsStore4[6]),
	.Weight7(WeightsStore4[7]),
	.Weight8(WeightsStore4[8]),
	.Weight9(WeightsStore4[9]),
	.Weight10(WeightsStore4[10]),
	.Weight11(WeightsStore4[11]),
	.Weight12(WeightsStore4[12]),
	.Weight13(WeightsStore4[13]),
	.Weight14(WeightsStore4[14]),
	.Weight15(WeightsStore4[15]),
	.Weight16(WeightsStore4[16]),
	.Weight17(WeightsStore4[17]),
	.Weight18(WeightsStore4[18]),
	.Weight19(WeightsStore4[19]),
	.Weight20(WeightsStore4[20]),
	.Weight21(WeightsStore4[21]),
	.Weight22(WeightsStore4[22]),
	.Weight23(WeightsStore4[23]),
	.Weight24(WeightsStore4[24]),
	.Weight25(WeightsStore4[25]),
	.Weight26(WeightsStore4[26]),
	.Weight27(WeightsStore4[27]),
	.value(vals[4])
	);
DotProduct784 DP5(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore5[0]),
	.Weight1(WeightsStore5[1]),
	.Weight2(WeightsStore5[2]),
	.Weight3(WeightsStore5[3]),
	.Weight4(WeightsStore5[4]),
	.Weight5(WeightsStore5[5]),
	.Weight6(WeightsStore5[6]),
	.Weight7(WeightsStore5[7]),
	.Weight8(WeightsStore5[8]),
	.Weight9(WeightsStore5[9]),
	.Weight10(WeightsStore5[10]),
	.Weight11(WeightsStore5[11]),
	.Weight12(WeightsStore5[12]),
	.Weight13(WeightsStore5[13]),
	.Weight14(WeightsStore5[14]),
	.Weight15(WeightsStore5[15]),
	.Weight16(WeightsStore5[16]),
	.Weight17(WeightsStore5[17]),
	.Weight18(WeightsStore5[18]),
	.Weight19(WeightsStore5[19]),
	.Weight20(WeightsStore5[20]),
	.Weight21(WeightsStore5[21]),
	.Weight22(WeightsStore5[22]),
	.Weight23(WeightsStore5[23]),
	.Weight24(WeightsStore5[24]),
	.Weight25(WeightsStore5[25]),
	.Weight26(WeightsStore5[26]),
	.Weight27(WeightsStore5[27]),
	.value(vals[5])
	);
DotProduct784 DP6(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore6[0]),
	.Weight1(WeightsStore6[1]),
	.Weight2(WeightsStore6[2]),
	.Weight3(WeightsStore6[3]),
	.Weight4(WeightsStore6[4]),
	.Weight5(WeightsStore6[5]),
	.Weight6(WeightsStore6[6]),
	.Weight7(WeightsStore6[7]),
	.Weight8(WeightsStore6[8]),
	.Weight9(WeightsStore6[9]),
	.Weight10(WeightsStore6[10]),
	.Weight11(WeightsStore6[11]),
	.Weight12(WeightsStore6[12]),
	.Weight13(WeightsStore6[13]),
	.Weight14(WeightsStore6[14]),
	.Weight15(WeightsStore6[15]),
	.Weight16(WeightsStore6[16]),
	.Weight17(WeightsStore6[17]),
	.Weight18(WeightsStore6[18]),
	.Weight19(WeightsStore6[19]),
	.Weight20(WeightsStore6[20]),
	.Weight21(WeightsStore6[21]),
	.Weight22(WeightsStore6[22]),
	.Weight23(WeightsStore6[23]),
	.Weight24(WeightsStore6[24]),
	.Weight25(WeightsStore6[25]),
	.Weight26(WeightsStore6[26]),
	.Weight27(WeightsStore6[27]),
	.value(vals[6])
	);
DotProduct784 DP7(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore7[0]),
	.Weight1(WeightsStore7[1]),
	.Weight2(WeightsStore7[2]),
	.Weight3(WeightsStore7[3]),
	.Weight4(WeightsStore7[4]),
	.Weight5(WeightsStore7[5]),
	.Weight6(WeightsStore7[6]),
	.Weight7(WeightsStore7[7]),
	.Weight8(WeightsStore7[8]),
	.Weight9(WeightsStore7[9]),
	.Weight10(WeightsStore7[10]),
	.Weight11(WeightsStore7[11]),
	.Weight12(WeightsStore7[12]),
	.Weight13(WeightsStore7[13]),
	.Weight14(WeightsStore7[14]),
	.Weight15(WeightsStore7[15]),
	.Weight16(WeightsStore7[16]),
	.Weight17(WeightsStore7[17]),
	.Weight18(WeightsStore7[18]),
	.Weight19(WeightsStore7[19]),
	.Weight20(WeightsStore7[20]),
	.Weight21(WeightsStore7[21]),
	.Weight22(WeightsStore7[22]),
	.Weight23(WeightsStore7[23]),
	.Weight24(WeightsStore7[24]),
	.Weight25(WeightsStore7[25]),
	.Weight26(WeightsStore7[26]),
	.Weight27(WeightsStore7[27]),
	.value(vals[7])
	);
DotProduct784 DP8(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore8[0]),
	.Weight1(WeightsStore8[1]),
	.Weight2(WeightsStore8[2]),
	.Weight3(WeightsStore8[3]),
	.Weight4(WeightsStore8[4]),
	.Weight5(WeightsStore8[5]),
	.Weight6(WeightsStore8[6]),
	.Weight7(WeightsStore8[7]),
	.Weight8(WeightsStore8[8]),
	.Weight9(WeightsStore8[9]),
	.Weight10(WeightsStore8[10]),
	.Weight11(WeightsStore8[11]),
	.Weight12(WeightsStore8[12]),
	.Weight13(WeightsStore8[13]),
	.Weight14(WeightsStore8[14]),
	.Weight15(WeightsStore8[15]),
	.Weight16(WeightsStore8[16]),
	.Weight17(WeightsStore8[17]),
	.Weight18(WeightsStore8[18]),
	.Weight19(WeightsStore8[19]),
	.Weight20(WeightsStore8[20]),
	.Weight21(WeightsStore8[21]),
	.Weight22(WeightsStore8[22]),
	.Weight23(WeightsStore8[23]),
	.Weight24(WeightsStore8[24]),
	.Weight25(WeightsStore8[25]),
	.Weight26(WeightsStore8[26]),
	.Weight27(WeightsStore8[27]),
	.value(vals[8])
	);
DotProduct784 DP9(.clk(clk),
	.GlobalReset(GlobalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore9[0]),
	.Weight1(WeightsStore9[1]),
	.Weight2(WeightsStore9[2]),
	.Weight3(WeightsStore9[3]),
	.Weight4(WeightsStore9[4]),
	.Weight5(WeightsStore9[5]),
	.Weight6(WeightsStore9[6]),
	.Weight7(WeightsStore9[7]),
	.Weight8(WeightsStore9[8]),
	.Weight9(WeightsStore9[9]),
	.Weight10(WeightsStore9[10]),
	.Weight11(WeightsStore9[11]),
	.Weight12(WeightsStore9[12]),
	.Weight13(WeightsStore9[13]),
	.Weight14(WeightsStore9[14]),
	.Weight15(WeightsStore9[15]),
	.Weight16(WeightsStore9[16]),
	.Weight17(WeightsStore9[17]),
	.Weight18(WeightsStore9[18]),
	.Weight19(WeightsStore9[19]),
	.Weight20(WeightsStore9[20]),
	.Weight21(WeightsStore9[21]),
	.Weight22(WeightsStore9[22]),
	.Weight23(WeightsStore9[23]),
	.Weight24(WeightsStore9[24]),
	.Weight25(WeightsStore9[25]),
	.Weight26(WeightsStore9[26]),
	.Weight27(WeightsStore9[27]),
	.value(vals[9])
	);

always@(posedge clk)begin
	if(GlobalReset == 1'b1)begin
		switchCounter <= 32'd0;
		PixelsStore[0] <= 10'd0;
		PixelsStore[1] <= 10'd0;
		PixelsStore[2] <= 10'd0;
		PixelsStore[3] <= 10'd0;
		PixelsStore[4] <= 10'd0;
		PixelsStore[5] <= 10'd0;
		PixelsStore[6] <= 10'd0;
		PixelsStore[7] <= 10'd0;
		PixelsStore[8] <= 10'd0;
		PixelsStore[9] <= 10'd0;
		PixelsStore[10] <= 10'd0;
		PixelsStore[11] <= 10'd0;
		PixelsStore[12] <= 10'd0;
		PixelsStore[13] <= 10'd0;
		PixelsStore[14] <= 10'd0;
		PixelsStore[15] <= 10'd0;
		PixelsStore[16] <= 10'd0;
		PixelsStore[17] <= 10'd0;
		PixelsStore[18] <= 10'd0;
		PixelsStore[19] <= 10'd0;
		PixelsStore[20] <= 10'd0;
		PixelsStore[21] <= 10'd0;
		PixelsStore[22] <= 10'd0;
		PixelsStore[23] <= 10'd0;
		PixelsStore[24] <= 10'd0;
		PixelsStore[25] <= 10'd0;
		PixelsStore[26] <= 10'd0;
		PixelsStore[27] <= 10'd0;
		WeightsStore0[0] <= 19'd0;
		WeightsStore0[1] <= 19'd0;
		WeightsStore0[2] <= 19'd0;
		WeightsStore0[3] <= 19'd0;
		WeightsStore0[4] <= 19'd0;
		WeightsStore0[5] <= 19'd0;
		WeightsStore0[6] <= 19'd0;
		WeightsStore0[7] <= 19'd0;
		WeightsStore0[8] <= 19'd0;
		WeightsStore0[9] <= 19'd0;
		WeightsStore0[10] <= 19'd0;
		WeightsStore0[11] <= 19'd0;
		WeightsStore0[12] <= 19'd0;
		WeightsStore0[13] <= 19'd0;
		WeightsStore0[14] <= 19'd0;
		WeightsStore0[15] <= 19'd0;
		WeightsStore0[16] <= 19'd0;
		WeightsStore0[17] <= 19'd0;
		WeightsStore0[18] <= 19'd0;
		WeightsStore0[19] <= 19'd0;
		WeightsStore0[20] <= 19'd0;
		WeightsStore0[21] <= 19'd0;
		WeightsStore0[22] <= 19'd0;
		WeightsStore0[23] <= 19'd0;
		WeightsStore0[24] <= 19'd0;
		WeightsStore0[25] <= 19'd0;
		WeightsStore0[26] <= 19'd0;
		WeightsStore0[27] <= 19'd0;
		WeightsStore1[0] <= 19'd0;
		WeightsStore1[1] <= 19'd0;
		WeightsStore1[2] <= 19'd0;
		WeightsStore1[3] <= 19'd0;
		WeightsStore1[4] <= 19'd0;
		WeightsStore1[5] <= 19'd0;
		WeightsStore1[6] <= 19'd0;
		WeightsStore1[7] <= 19'd0;
		WeightsStore1[8] <= 19'd0;
		WeightsStore1[9] <= 19'd0;
		WeightsStore1[10] <= 19'd0;
		WeightsStore1[11] <= 19'd0;
		WeightsStore1[12] <= 19'd0;
		WeightsStore1[13] <= 19'd0;
		WeightsStore1[14] <= 19'd0;
		WeightsStore1[15] <= 19'd0;
		WeightsStore1[16] <= 19'd0;
		WeightsStore1[17] <= 19'd0;
		WeightsStore1[18] <= 19'd0;
		WeightsStore1[19] <= 19'd0;
		WeightsStore1[20] <= 19'd0;
		WeightsStore1[21] <= 19'd0;
		WeightsStore1[22] <= 19'd0;
		WeightsStore1[23] <= 19'd0;
		WeightsStore1[24] <= 19'd0;
		WeightsStore1[25] <= 19'd0;
		WeightsStore1[26] <= 19'd0;
		WeightsStore1[27] <= 19'd0;
		WeightsStore2[0] <= 19'd0;
		WeightsStore2[1] <= 19'd0;
		WeightsStore2[2] <= 19'd0;
		WeightsStore2[3] <= 19'd0;
		WeightsStore2[4] <= 19'd0;
		WeightsStore2[5] <= 19'd0;
		WeightsStore2[6] <= 19'd0;
		WeightsStore2[7] <= 19'd0;
		WeightsStore2[8] <= 19'd0;
		WeightsStore2[9] <= 19'd0;
		WeightsStore2[10] <= 19'd0;
		WeightsStore2[11] <= 19'd0;
		WeightsStore2[12] <= 19'd0;
		WeightsStore2[13] <= 19'd0;
		WeightsStore2[14] <= 19'd0;
		WeightsStore2[15] <= 19'd0;
		WeightsStore2[16] <= 19'd0;
		WeightsStore2[17] <= 19'd0;
		WeightsStore2[18] <= 19'd0;
		WeightsStore2[19] <= 19'd0;
		WeightsStore2[20] <= 19'd0;
		WeightsStore2[21] <= 19'd0;
		WeightsStore2[22] <= 19'd0;
		WeightsStore2[23] <= 19'd0;
		WeightsStore2[24] <= 19'd0;
		WeightsStore2[25] <= 19'd0;
		WeightsStore2[26] <= 19'd0;
		WeightsStore2[27] <= 19'd0;
		WeightsStore3[0] <= 19'd0;
		WeightsStore3[1] <= 19'd0;
		WeightsStore3[2] <= 19'd0;
		WeightsStore3[3] <= 19'd0;
		WeightsStore3[4] <= 19'd0;
		WeightsStore3[5] <= 19'd0;
		WeightsStore3[6] <= 19'd0;
		WeightsStore3[7] <= 19'd0;
		WeightsStore3[8] <= 19'd0;
		WeightsStore3[9] <= 19'd0;
		WeightsStore3[10] <= 19'd0;
		WeightsStore3[11] <= 19'd0;
		WeightsStore3[12] <= 19'd0;
		WeightsStore3[13] <= 19'd0;
		WeightsStore3[14] <= 19'd0;
		WeightsStore3[15] <= 19'd0;
		WeightsStore3[16] <= 19'd0;
		WeightsStore3[17] <= 19'd0;
		WeightsStore3[18] <= 19'd0;
		WeightsStore3[19] <= 19'd0;
		WeightsStore3[20] <= 19'd0;
		WeightsStore3[21] <= 19'd0;
		WeightsStore3[22] <= 19'd0;
		WeightsStore3[23] <= 19'd0;
		WeightsStore3[24] <= 19'd0;
		WeightsStore3[25] <= 19'd0;
		WeightsStore3[26] <= 19'd0;
		WeightsStore3[27] <= 19'd0;
		WeightsStore4[0] <= 19'd0;
		WeightsStore4[1] <= 19'd0;
		WeightsStore4[2] <= 19'd0;
		WeightsStore4[3] <= 19'd0;
		WeightsStore4[4] <= 19'd0;
		WeightsStore4[5] <= 19'd0;
		WeightsStore4[6] <= 19'd0;
		WeightsStore4[7] <= 19'd0;
		WeightsStore4[8] <= 19'd0;
		WeightsStore4[9] <= 19'd0;
		WeightsStore4[10] <= 19'd0;
		WeightsStore4[11] <= 19'd0;
		WeightsStore4[12] <= 19'd0;
		WeightsStore4[13] <= 19'd0;
		WeightsStore4[14] <= 19'd0;
		WeightsStore4[15] <= 19'd0;
		WeightsStore4[16] <= 19'd0;
		WeightsStore4[17] <= 19'd0;
		WeightsStore4[18] <= 19'd0;
		WeightsStore4[19] <= 19'd0;
		WeightsStore4[20] <= 19'd0;
		WeightsStore4[21] <= 19'd0;
		WeightsStore4[22] <= 19'd0;
		WeightsStore4[23] <= 19'd0;
		WeightsStore4[24] <= 19'd0;
		WeightsStore4[25] <= 19'd0;
		WeightsStore4[26] <= 19'd0;
		WeightsStore4[27] <= 19'd0;
		WeightsStore5[0] <= 19'd0;
		WeightsStore5[1] <= 19'd0;
		WeightsStore5[2] <= 19'd0;
		WeightsStore5[3] <= 19'd0;
		WeightsStore5[4] <= 19'd0;
		WeightsStore5[5] <= 19'd0;
		WeightsStore5[6] <= 19'd0;
		WeightsStore5[7] <= 19'd0;
		WeightsStore5[8] <= 19'd0;
		WeightsStore5[9] <= 19'd0;
		WeightsStore5[10] <= 19'd0;
		WeightsStore5[11] <= 19'd0;
		WeightsStore5[12] <= 19'd0;
		WeightsStore5[13] <= 19'd0;
		WeightsStore5[14] <= 19'd0;
		WeightsStore5[15] <= 19'd0;
		WeightsStore5[16] <= 19'd0;
		WeightsStore5[17] <= 19'd0;
		WeightsStore5[18] <= 19'd0;
		WeightsStore5[19] <= 19'd0;
		WeightsStore5[20] <= 19'd0;
		WeightsStore5[21] <= 19'd0;
		WeightsStore5[22] <= 19'd0;
		WeightsStore5[23] <= 19'd0;
		WeightsStore5[24] <= 19'd0;
		WeightsStore5[25] <= 19'd0;
		WeightsStore5[26] <= 19'd0;
		WeightsStore5[27] <= 19'd0;
		WeightsStore6[0] <= 19'd0;
		WeightsStore6[1] <= 19'd0;
		WeightsStore6[2] <= 19'd0;
		WeightsStore6[3] <= 19'd0;
		WeightsStore6[4] <= 19'd0;
		WeightsStore6[5] <= 19'd0;
		WeightsStore6[6] <= 19'd0;
		WeightsStore6[7] <= 19'd0;
		WeightsStore6[8] <= 19'd0;
		WeightsStore6[9] <= 19'd0;
		WeightsStore6[10] <= 19'd0;
		WeightsStore6[11] <= 19'd0;
		WeightsStore6[12] <= 19'd0;
		WeightsStore6[13] <= 19'd0;
		WeightsStore6[14] <= 19'd0;
		WeightsStore6[15] <= 19'd0;
		WeightsStore6[16] <= 19'd0;
		WeightsStore6[17] <= 19'd0;
		WeightsStore6[18] <= 19'd0;
		WeightsStore6[19] <= 19'd0;
		WeightsStore6[20] <= 19'd0;
		WeightsStore6[21] <= 19'd0;
		WeightsStore6[22] <= 19'd0;
		WeightsStore6[23] <= 19'd0;
		WeightsStore6[24] <= 19'd0;
		WeightsStore6[25] <= 19'd0;
		WeightsStore6[26] <= 19'd0;
		WeightsStore6[27] <= 19'd0;
		WeightsStore7[0] <= 19'd0;
		WeightsStore7[1] <= 19'd0;
		WeightsStore7[2] <= 19'd0;
		WeightsStore7[3] <= 19'd0;
		WeightsStore7[4] <= 19'd0;
		WeightsStore7[5] <= 19'd0;
		WeightsStore7[6] <= 19'd0;
		WeightsStore7[7] <= 19'd0;
		WeightsStore7[8] <= 19'd0;
		WeightsStore7[9] <= 19'd0;
		WeightsStore7[10] <= 19'd0;
		WeightsStore7[11] <= 19'd0;
		WeightsStore7[12] <= 19'd0;
		WeightsStore7[13] <= 19'd0;
		WeightsStore7[14] <= 19'd0;
		WeightsStore7[15] <= 19'd0;
		WeightsStore7[16] <= 19'd0;
		WeightsStore7[17] <= 19'd0;
		WeightsStore7[18] <= 19'd0;
		WeightsStore7[19] <= 19'd0;
		WeightsStore7[20] <= 19'd0;
		WeightsStore7[21] <= 19'd0;
		WeightsStore7[22] <= 19'd0;
		WeightsStore7[23] <= 19'd0;
		WeightsStore7[24] <= 19'd0;
		WeightsStore7[25] <= 19'd0;
		WeightsStore7[26] <= 19'd0;
		WeightsStore7[27] <= 19'd0;
		WeightsStore8[0] <= 19'd0;
		WeightsStore8[1] <= 19'd0;
		WeightsStore8[2] <= 19'd0;
		WeightsStore8[3] <= 19'd0;
		WeightsStore8[4] <= 19'd0;
		WeightsStore8[5] <= 19'd0;
		WeightsStore8[6] <= 19'd0;
		WeightsStore8[7] <= 19'd0;
		WeightsStore8[8] <= 19'd0;
		WeightsStore8[9] <= 19'd0;
		WeightsStore8[10] <= 19'd0;
		WeightsStore8[11] <= 19'd0;
		WeightsStore8[12] <= 19'd0;
		WeightsStore8[13] <= 19'd0;
		WeightsStore8[14] <= 19'd0;
		WeightsStore8[15] <= 19'd0;
		WeightsStore8[16] <= 19'd0;
		WeightsStore8[17] <= 19'd0;
		WeightsStore8[18] <= 19'd0;
		WeightsStore8[19] <= 19'd0;
		WeightsStore8[20] <= 19'd0;
		WeightsStore8[21] <= 19'd0;
		WeightsStore8[22] <= 19'd0;
		WeightsStore8[23] <= 19'd0;
		WeightsStore8[24] <= 19'd0;
		WeightsStore8[25] <= 19'd0;
		WeightsStore8[26] <= 19'd0;
		WeightsStore8[27] <= 19'd0;
		WeightsStore9[0] <= 19'd0;
		WeightsStore9[1] <= 19'd0;
		WeightsStore9[2] <= 19'd0;
		WeightsStore9[3] <= 19'd0;
		WeightsStore9[4] <= 19'd0;
		WeightsStore9[5] <= 19'd0;
		WeightsStore9[6] <= 19'd0;
		WeightsStore9[7] <= 19'd0;
		WeightsStore9[8] <= 19'd0;
		WeightsStore9[9] <= 19'd0;
		WeightsStore9[10] <= 19'd0;
		WeightsStore9[11] <= 19'd0;
		WeightsStore9[12] <= 19'd0;
		WeightsStore9[13] <= 19'd0;
		WeightsStore9[14] <= 19'd0;
		WeightsStore9[15] <= 19'd0;
		WeightsStore9[16] <= 19'd0;
		WeightsStore9[17] <= 19'd0;
		WeightsStore9[18] <= 19'd0;
		WeightsStore9[19] <= 19'd0;
		WeightsStore9[20] <= 19'd0;
		WeightsStore9[21] <= 19'd0;
		WeightsStore9[22] <= 19'd0;
		WeightsStore9[23] <= 19'd0;
		WeightsStore9[24] <= 19'd0;
		WeightsStore9[25] <= 19'd0;
		WeightsStore9[26] <= 19'd0;
		WeightsStore9[27] <= 19'd0;
	end else begin
		if(switchCounter == 32'd0)begin
			PixelsStore[0] <= Pixels[(32'd0+32'd1)*32'd10-1:32'd0*32'd10];
			PixelsStore[1] <= Pixels[(32'd1+32'd1)*32'd10-1:32'd1*32'd10];
			PixelsStore[2] <= Pixels[(32'd2+32'd1)*32'd10-1:32'd2*32'd10];
			PixelsStore[3] <= Pixels[(32'd3+32'd1)*32'd10-1:32'd3*32'd10];
			PixelsStore[4] <= Pixels[(32'd4+32'd1)*32'd10-1:32'd4*32'd10];
			PixelsStore[5] <= Pixels[(32'd5+32'd1)*32'd10-1:32'd5*32'd10];
			PixelsStore[6] <= Pixels[(32'd6+32'd1)*32'd10-1:32'd6*32'd10];
			PixelsStore[7] <= Pixels[(32'd7+32'd1)*32'd10-1:32'd7*32'd10];
			PixelsStore[8] <= Pixels[(32'd8+32'd1)*32'd10-1:32'd8*32'd10];
			PixelsStore[9] <= Pixels[(32'd9+32'd1)*32'd10-1:32'd9*32'd10];
			PixelsStore[10] <= Pixels[(32'd10+32'd1)*32'd10-1:32'd10*32'd10];
			PixelsStore[11] <= Pixels[(32'd11+32'd1)*32'd10-1:32'd11*32'd10];
			PixelsStore[12] <= Pixels[(32'd12+32'd1)*32'd10-1:32'd12*32'd10];
			PixelsStore[13] <= Pixels[(32'd13+32'd1)*32'd10-1:32'd13*32'd10];
			PixelsStore[14] <= Pixels[(32'd14+32'd1)*32'd10-1:32'd14*32'd10];
			PixelsStore[15] <= Pixels[(32'd15+32'd1)*32'd10-1:32'd15*32'd10];
			PixelsStore[16] <= Pixels[(32'd16+32'd1)*32'd10-1:32'd16*32'd10];
			PixelsStore[17] <= Pixels[(32'd17+32'd1)*32'd10-1:32'd17*32'd10];
			PixelsStore[18] <= Pixels[(32'd18+32'd1)*32'd10-1:32'd18*32'd10];
			PixelsStore[19] <= Pixels[(32'd19+32'd1)*32'd10-1:32'd19*32'd10];
			PixelsStore[20] <= Pixels[(32'd20+32'd1)*32'd10-1:32'd20*32'd10];
			PixelsStore[21] <= Pixels[(32'd21+32'd1)*32'd10-1:32'd21*32'd10];
			PixelsStore[22] <= Pixels[(32'd22+32'd1)*32'd10-1:32'd22*32'd10];
			PixelsStore[23] <= Pixels[(32'd23+32'd1)*32'd10-1:32'd23*32'd10];
			PixelsStore[24] <= Pixels[(32'd24+32'd1)*32'd10-1:32'd24*32'd10];
			PixelsStore[25] <= Pixels[(32'd25+32'd1)*32'd10-1:32'd25*32'd10];
			PixelsStore[26] <= Pixels[(32'd26+32'd1)*32'd10-1:32'd26*32'd10];
			PixelsStore[27] <= Pixels[(32'd27+32'd1)*32'd10-1:32'd27*32'd10];
			WeightsStore0[0] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[1] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[2] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[3] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[4] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[5] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[6] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[7] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[8] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[9] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[10] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[11] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[12] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[13] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[14] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[15] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[16] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[17] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[18] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[19] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[20] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[21] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[22] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[23] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[24] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[25] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[26] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore0[27] <= Weights0[(32'd0+32'd1)*32'd19-1:32'd0*32'd19];
			WeightsStore1[0] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[1] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[2] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[3] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[4] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[5] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[6] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[7] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[8] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[9] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[10] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[11] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[12] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[13] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[14] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[15] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[16] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[17] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[18] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[19] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[20] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[21] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[22] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[23] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[24] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[25] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[26] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore1[27] <= Weights1[(32'd1+32'd1)*32'd19-1:32'd1*32'd19];
			WeightsStore2[0] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[1] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[2] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[3] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[4] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[5] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[6] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[7] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[8] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[9] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[10] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[11] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[12] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[13] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[14] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[15] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[16] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[17] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[18] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[19] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[20] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[21] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[22] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[23] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[24] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[25] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[26] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore2[27] <= Weights2[(32'd2+32'd1)*32'd19-1:32'd2*32'd19];
			WeightsStore3[0] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[1] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[2] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[3] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[4] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[5] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[6] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[7] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[8] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[9] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[10] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[11] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[12] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[13] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[14] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[15] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[16] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[17] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[18] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[19] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[20] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[21] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[22] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[23] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[24] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[25] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[26] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore3[27] <= Weights3[(32'd3+32'd1)*32'd19-1:32'd3*32'd19];
			WeightsStore4[0] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[1] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[2] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[3] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[4] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[5] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[6] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[7] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[8] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[9] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[10] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[11] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[12] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[13] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[14] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[15] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[16] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[17] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[18] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[19] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[20] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[21] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[22] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[23] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[24] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[25] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[26] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore4[27] <= Weights4[(32'd4+32'd1)*32'd19-1:32'd4*32'd19];
			WeightsStore5[0] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[1] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[2] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[3] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[4] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[5] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[6] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[7] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[8] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[9] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[10] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[11] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[12] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[13] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[14] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[15] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[16] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[17] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[18] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[19] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[20] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[21] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[22] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[23] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[24] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[25] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[26] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore5[27] <= Weights5[(32'd5+32'd1)*32'd19-1:32'd5*32'd19];
			WeightsStore6[0] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[1] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[2] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[3] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[4] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[5] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[6] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[7] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[8] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[9] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[10] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[11] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[12] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[13] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[14] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[15] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[16] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[17] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[18] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[19] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[20] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[21] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[22] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[23] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[24] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[25] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[26] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore6[27] <= Weights6[(32'd6+32'd1)*32'd19-1:32'd6*32'd19];
			WeightsStore7[0] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[1] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[2] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[3] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[4] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[5] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[6] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[7] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[8] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[9] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[10] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[11] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[12] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[13] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[14] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[15] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[16] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[17] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[18] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[19] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[20] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[21] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[22] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[23] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[24] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[25] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[26] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore7[27] <= Weights7[(32'd7+32'd1)*32'd19-1:32'd7*32'd19];
			WeightsStore8[0] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[1] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[2] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[3] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[4] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[5] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[6] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[7] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[8] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[9] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[10] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[11] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[12] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[13] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[14] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[15] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[16] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[17] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[18] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[19] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[20] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[21] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[22] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[23] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[24] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[25] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[26] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore8[27] <= Weights8[(32'd8+32'd1)*32'd19-1:32'd8*32'd19];
			WeightsStore9[0] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[1] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[2] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[3] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[4] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[5] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[6] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[7] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[8] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[9] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[10] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[11] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[12] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[13] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[14] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[15] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[16] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[17] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[18] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[19] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[20] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[21] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[22] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[23] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[24] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[25] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[26] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
			WeightsStore9[27] <= Weights9[(32'd9+32'd1)*32'd19-1:32'd9*32'd19];
		end else if(switchCounter == 32'd1)begin
			PixelsStore[0] <= Pixels[(32'd28+32'd1)*32'd10-1:32'd28*32'd10];
			PixelsStore[1] <= Pixels[(32'd29+32'd1)*32'd10-1:32'd29*32'd10];
			PixelsStore[2] <= Pixels[(32'd30+32'd1)*32'd10-1:32'd30*32'd10];
			PixelsStore[3] <= Pixels[(32'd31+32'd1)*32'd10-1:32'd31*32'd10];
			PixelsStore[4] <= Pixels[(32'd32+32'd1)*32'd10-1:32'd32*32'd10];
			PixelsStore[5] <= Pixels[(32'd33+32'd1)*32'd10-1:32'd33*32'd10];
			PixelsStore[6] <= Pixels[(32'd34+32'd1)*32'd10-1:32'd34*32'd10];
			PixelsStore[7] <= Pixels[(32'd35+32'd1)*32'd10-1:32'd35*32'd10];
			PixelsStore[8] <= Pixels[(32'd36+32'd1)*32'd10-1:32'd36*32'd10];
			PixelsStore[9] <= Pixels[(32'd37+32'd1)*32'd10-1:32'd37*32'd10];
			PixelsStore[10] <= Pixels[(32'd38+32'd1)*32'd10-1:32'd38*32'd10];
			PixelsStore[11] <= Pixels[(32'd39+32'd1)*32'd10-1:32'd39*32'd10];
			PixelsStore[12] <= Pixels[(32'd40+32'd1)*32'd10-1:32'd40*32'd10];
			PixelsStore[13] <= Pixels[(32'd41+32'd1)*32'd10-1:32'd41*32'd10];
			PixelsStore[14] <= Pixels[(32'd42+32'd1)*32'd10-1:32'd42*32'd10];
			PixelsStore[15] <= Pixels[(32'd43+32'd1)*32'd10-1:32'd43*32'd10];
			PixelsStore[16] <= Pixels[(32'd44+32'd1)*32'd10-1:32'd44*32'd10];
			PixelsStore[17] <= Pixels[(32'd45+32'd1)*32'd10-1:32'd45*32'd10];
			PixelsStore[18] <= Pixels[(32'd46+32'd1)*32'd10-1:32'd46*32'd10];
			PixelsStore[19] <= Pixels[(32'd47+32'd1)*32'd10-1:32'd47*32'd10];
			PixelsStore[20] <= Pixels[(32'd48+32'd1)*32'd10-1:32'd48*32'd10];
			PixelsStore[21] <= Pixels[(32'd49+32'd1)*32'd10-1:32'd49*32'd10];
			PixelsStore[22] <= Pixels[(32'd50+32'd1)*32'd10-1:32'd50*32'd10];
			PixelsStore[23] <= Pixels[(32'd51+32'd1)*32'd10-1:32'd51*32'd10];
			PixelsStore[24] <= Pixels[(32'd52+32'd1)*32'd10-1:32'd52*32'd10];
			PixelsStore[25] <= Pixels[(32'd53+32'd1)*32'd10-1:32'd53*32'd10];
			PixelsStore[26] <= Pixels[(32'd54+32'd1)*32'd10-1:32'd54*32'd10];
			PixelsStore[27] <= Pixels[(32'd55+32'd1)*32'd10-1:32'd55*32'd10];
			WeightsStore0[0] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[1] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[2] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[3] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[4] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[5] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[6] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[7] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[8] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[9] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[10] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[11] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[12] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[13] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[14] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[15] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[16] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[17] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[18] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[19] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[20] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[21] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[22] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[23] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[24] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[25] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[26] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore0[27] <= Weights0[(32'd28+32'd1)*32'd19-1:32'd28*32'd19];
			WeightsStore1[0] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[1] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[2] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[3] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[4] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[5] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[6] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[7] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[8] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[9] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[10] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[11] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[12] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[13] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[14] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[15] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[16] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[17] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[18] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[19] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[20] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[21] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[22] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[23] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[24] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[25] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[26] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore1[27] <= Weights1[(32'd29+32'd1)*32'd19-1:32'd29*32'd19];
			WeightsStore2[0] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[1] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[2] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[3] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[4] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[5] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[6] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[7] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[8] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[9] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[10] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[11] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[12] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[13] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[14] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[15] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[16] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[17] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[18] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[19] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[20] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[21] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[22] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[23] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[24] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[25] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[26] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore2[27] <= Weights2[(32'd30+32'd1)*32'd19-1:32'd30*32'd19];
			WeightsStore3[0] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[1] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[2] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[3] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[4] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[5] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[6] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[7] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[8] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[9] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[10] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[11] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[12] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[13] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[14] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[15] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[16] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[17] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[18] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[19] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[20] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[21] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[22] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[23] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[24] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[25] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[26] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore3[27] <= Weights3[(32'd31+32'd1)*32'd19-1:32'd31*32'd19];
			WeightsStore4[0] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[1] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[2] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[3] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[4] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[5] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[6] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[7] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[8] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[9] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[10] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[11] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[12] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[13] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[14] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[15] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[16] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[17] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[18] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[19] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[20] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[21] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[22] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[23] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[24] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[25] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[26] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore4[27] <= Weights4[(32'd32+32'd1)*32'd19-1:32'd32*32'd19];
			WeightsStore5[0] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[1] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[2] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[3] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[4] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[5] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[6] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[7] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[8] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[9] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[10] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[11] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[12] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[13] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[14] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[15] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[16] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[17] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[18] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[19] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[20] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[21] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[22] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[23] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[24] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[25] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[26] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore5[27] <= Weights5[(32'd33+32'd1)*32'd19-1:32'd33*32'd19];
			WeightsStore6[0] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[1] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[2] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[3] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[4] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[5] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[6] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[7] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[8] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[9] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[10] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[11] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[12] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[13] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[14] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[15] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[16] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[17] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[18] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[19] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[20] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[21] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[22] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[23] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[24] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[25] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[26] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore6[27] <= Weights6[(32'd34+32'd1)*32'd19-1:32'd34*32'd19];
			WeightsStore7[0] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[1] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[2] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[3] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[4] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[5] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[6] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[7] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[8] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[9] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[10] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[11] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[12] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[13] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[14] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[15] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[16] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[17] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[18] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[19] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[20] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[21] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[22] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[23] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[24] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[25] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[26] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore7[27] <= Weights7[(32'd35+32'd1)*32'd19-1:32'd35*32'd19];
			WeightsStore8[0] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[1] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[2] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[3] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[4] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[5] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[6] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[7] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[8] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[9] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[10] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[11] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[12] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[13] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[14] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[15] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[16] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[17] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[18] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[19] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[20] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[21] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[22] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[23] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[24] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[25] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[26] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore8[27] <= Weights8[(32'd36+32'd1)*32'd19-1:32'd36*32'd19];
			WeightsStore9[0] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[1] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[2] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[3] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[4] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[5] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[6] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[7] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[8] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[9] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[10] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[11] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[12] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[13] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[14] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[15] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[16] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[17] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[18] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[19] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[20] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[21] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[22] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[23] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[24] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[25] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[26] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
			WeightsStore9[27] <= Weights9[(32'd37+32'd1)*32'd19-1:32'd37*32'd19];
		end else if(switchCounter == 32'd2)begin
			PixelsStore[0] <= Pixels[(32'd56+32'd1)*32'd10-1:32'd56*32'd10];
			PixelsStore[1] <= Pixels[(32'd57+32'd1)*32'd10-1:32'd57*32'd10];
			PixelsStore[2] <= Pixels[(32'd58+32'd1)*32'd10-1:32'd58*32'd10];
			PixelsStore[3] <= Pixels[(32'd59+32'd1)*32'd10-1:32'd59*32'd10];
			PixelsStore[4] <= Pixels[(32'd60+32'd1)*32'd10-1:32'd60*32'd10];
			PixelsStore[5] <= Pixels[(32'd61+32'd1)*32'd10-1:32'd61*32'd10];
			PixelsStore[6] <= Pixels[(32'd62+32'd1)*32'd10-1:32'd62*32'd10];
			PixelsStore[7] <= Pixels[(32'd63+32'd1)*32'd10-1:32'd63*32'd10];
			PixelsStore[8] <= Pixels[(32'd64+32'd1)*32'd10-1:32'd64*32'd10];
			PixelsStore[9] <= Pixels[(32'd65+32'd1)*32'd10-1:32'd65*32'd10];
			PixelsStore[10] <= Pixels[(32'd66+32'd1)*32'd10-1:32'd66*32'd10];
			PixelsStore[11] <= Pixels[(32'd67+32'd1)*32'd10-1:32'd67*32'd10];
			PixelsStore[12] <= Pixels[(32'd68+32'd1)*32'd10-1:32'd68*32'd10];
			PixelsStore[13] <= Pixels[(32'd69+32'd1)*32'd10-1:32'd69*32'd10];
			PixelsStore[14] <= Pixels[(32'd70+32'd1)*32'd10-1:32'd70*32'd10];
			PixelsStore[15] <= Pixels[(32'd71+32'd1)*32'd10-1:32'd71*32'd10];
			PixelsStore[16] <= Pixels[(32'd72+32'd1)*32'd10-1:32'd72*32'd10];
			PixelsStore[17] <= Pixels[(32'd73+32'd1)*32'd10-1:32'd73*32'd10];
			PixelsStore[18] <= Pixels[(32'd74+32'd1)*32'd10-1:32'd74*32'd10];
			PixelsStore[19] <= Pixels[(32'd75+32'd1)*32'd10-1:32'd75*32'd10];
			PixelsStore[20] <= Pixels[(32'd76+32'd1)*32'd10-1:32'd76*32'd10];
			PixelsStore[21] <= Pixels[(32'd77+32'd1)*32'd10-1:32'd77*32'd10];
			PixelsStore[22] <= Pixels[(32'd78+32'd1)*32'd10-1:32'd78*32'd10];
			PixelsStore[23] <= Pixels[(32'd79+32'd1)*32'd10-1:32'd79*32'd10];
			PixelsStore[24] <= Pixels[(32'd80+32'd1)*32'd10-1:32'd80*32'd10];
			PixelsStore[25] <= Pixels[(32'd81+32'd1)*32'd10-1:32'd81*32'd10];
			PixelsStore[26] <= Pixels[(32'd82+32'd1)*32'd10-1:32'd82*32'd10];
			PixelsStore[27] <= Pixels[(32'd83+32'd1)*32'd10-1:32'd83*32'd10];
			WeightsStore0[0] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[1] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[2] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[3] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[4] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[5] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[6] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[7] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[8] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[9] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[10] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[11] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[12] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[13] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[14] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[15] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[16] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[17] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[18] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[19] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[20] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[21] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[22] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[23] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[24] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[25] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[26] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore0[27] <= Weights0[(32'd56+32'd1)*32'd19-1:32'd56*32'd19];
			WeightsStore1[0] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[1] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[2] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[3] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[4] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[5] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[6] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[7] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[8] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[9] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[10] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[11] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[12] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[13] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[14] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[15] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[16] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[17] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[18] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[19] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[20] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[21] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[22] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[23] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[24] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[25] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[26] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore1[27] <= Weights1[(32'd57+32'd1)*32'd19-1:32'd57*32'd19];
			WeightsStore2[0] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[1] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[2] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[3] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[4] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[5] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[6] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[7] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[8] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[9] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[10] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[11] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[12] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[13] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[14] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[15] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[16] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[17] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[18] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[19] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[20] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[21] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[22] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[23] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[24] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[25] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[26] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore2[27] <= Weights2[(32'd58+32'd1)*32'd19-1:32'd58*32'd19];
			WeightsStore3[0] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[1] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[2] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[3] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[4] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[5] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[6] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[7] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[8] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[9] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[10] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[11] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[12] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[13] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[14] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[15] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[16] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[17] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[18] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[19] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[20] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[21] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[22] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[23] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[24] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[25] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[26] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore3[27] <= Weights3[(32'd59+32'd1)*32'd19-1:32'd59*32'd19];
			WeightsStore4[0] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[1] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[2] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[3] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[4] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[5] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[6] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[7] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[8] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[9] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[10] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[11] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[12] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[13] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[14] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[15] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[16] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[17] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[18] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[19] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[20] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[21] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[22] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[23] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[24] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[25] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[26] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore4[27] <= Weights4[(32'd60+32'd1)*32'd19-1:32'd60*32'd19];
			WeightsStore5[0] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[1] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[2] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[3] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[4] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[5] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[6] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[7] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[8] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[9] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[10] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[11] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[12] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[13] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[14] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[15] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[16] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[17] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[18] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[19] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[20] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[21] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[22] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[23] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[24] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[25] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[26] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore5[27] <= Weights5[(32'd61+32'd1)*32'd19-1:32'd61*32'd19];
			WeightsStore6[0] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[1] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[2] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[3] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[4] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[5] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[6] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[7] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[8] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[9] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[10] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[11] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[12] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[13] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[14] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[15] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[16] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[17] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[18] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[19] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[20] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[21] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[22] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[23] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[24] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[25] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[26] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore6[27] <= Weights6[(32'd62+32'd1)*32'd19-1:32'd62*32'd19];
			WeightsStore7[0] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[1] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[2] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[3] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[4] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[5] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[6] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[7] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[8] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[9] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[10] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[11] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[12] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[13] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[14] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[15] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[16] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[17] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[18] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[19] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[20] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[21] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[22] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[23] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[24] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[25] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[26] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore7[27] <= Weights7[(32'd63+32'd1)*32'd19-1:32'd63*32'd19];
			WeightsStore8[0] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[1] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[2] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[3] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[4] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[5] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[6] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[7] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[8] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[9] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[10] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[11] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[12] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[13] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[14] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[15] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[16] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[17] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[18] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[19] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[20] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[21] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[22] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[23] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[24] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[25] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[26] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore8[27] <= Weights8[(32'd64+32'd1)*32'd19-1:32'd64*32'd19];
			WeightsStore9[0] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[1] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[2] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[3] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[4] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[5] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[6] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[7] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[8] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[9] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[10] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[11] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[12] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[13] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[14] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[15] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[16] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[17] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[18] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[19] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[20] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[21] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[22] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[23] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[24] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[25] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[26] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
			WeightsStore9[27] <= Weights9[(32'd65+32'd1)*32'd19-1:32'd65*32'd19];
		end else if(switchCounter == 32'd3)begin
			PixelsStore[0] <= Pixels[(32'd84+32'd1)*32'd10-1:32'd84*32'd10];
			PixelsStore[1] <= Pixels[(32'd85+32'd1)*32'd10-1:32'd85*32'd10];
			PixelsStore[2] <= Pixels[(32'd86+32'd1)*32'd10-1:32'd86*32'd10];
			PixelsStore[3] <= Pixels[(32'd87+32'd1)*32'd10-1:32'd87*32'd10];
			PixelsStore[4] <= Pixels[(32'd88+32'd1)*32'd10-1:32'd88*32'd10];
			PixelsStore[5] <= Pixels[(32'd89+32'd1)*32'd10-1:32'd89*32'd10];
			PixelsStore[6] <= Pixels[(32'd90+32'd1)*32'd10-1:32'd90*32'd10];
			PixelsStore[7] <= Pixels[(32'd91+32'd1)*32'd10-1:32'd91*32'd10];
			PixelsStore[8] <= Pixels[(32'd92+32'd1)*32'd10-1:32'd92*32'd10];
			PixelsStore[9] <= Pixels[(32'd93+32'd1)*32'd10-1:32'd93*32'd10];
			PixelsStore[10] <= Pixels[(32'd94+32'd1)*32'd10-1:32'd94*32'd10];
			PixelsStore[11] <= Pixels[(32'd95+32'd1)*32'd10-1:32'd95*32'd10];
			PixelsStore[12] <= Pixels[(32'd96+32'd1)*32'd10-1:32'd96*32'd10];
			PixelsStore[13] <= Pixels[(32'd97+32'd1)*32'd10-1:32'd97*32'd10];
			PixelsStore[14] <= Pixels[(32'd98+32'd1)*32'd10-1:32'd98*32'd10];
			PixelsStore[15] <= Pixels[(32'd99+32'd1)*32'd10-1:32'd99*32'd10];
			PixelsStore[16] <= Pixels[(32'd100+32'd1)*32'd10-1:32'd100*32'd10];
			PixelsStore[17] <= Pixels[(32'd101+32'd1)*32'd10-1:32'd101*32'd10];
			PixelsStore[18] <= Pixels[(32'd102+32'd1)*32'd10-1:32'd102*32'd10];
			PixelsStore[19] <= Pixels[(32'd103+32'd1)*32'd10-1:32'd103*32'd10];
			PixelsStore[20] <= Pixels[(32'd104+32'd1)*32'd10-1:32'd104*32'd10];
			PixelsStore[21] <= Pixels[(32'd105+32'd1)*32'd10-1:32'd105*32'd10];
			PixelsStore[22] <= Pixels[(32'd106+32'd1)*32'd10-1:32'd106*32'd10];
			PixelsStore[23] <= Pixels[(32'd107+32'd1)*32'd10-1:32'd107*32'd10];
			PixelsStore[24] <= Pixels[(32'd108+32'd1)*32'd10-1:32'd108*32'd10];
			PixelsStore[25] <= Pixels[(32'd109+32'd1)*32'd10-1:32'd109*32'd10];
			PixelsStore[26] <= Pixels[(32'd110+32'd1)*32'd10-1:32'd110*32'd10];
			PixelsStore[27] <= Pixels[(32'd111+32'd1)*32'd10-1:32'd111*32'd10];
			WeightsStore0[0] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[1] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[2] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[3] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[4] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[5] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[6] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[7] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[8] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[9] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[10] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[11] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[12] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[13] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[14] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[15] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[16] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[17] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[18] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[19] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[20] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[21] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[22] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[23] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[24] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[25] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[26] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore0[27] <= Weights0[(32'd84+32'd1)*32'd19-1:32'd84*32'd19];
			WeightsStore1[0] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[1] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[2] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[3] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[4] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[5] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[6] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[7] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[8] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[9] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[10] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[11] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[12] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[13] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[14] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[15] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[16] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[17] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[18] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[19] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[20] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[21] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[22] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[23] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[24] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[25] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[26] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore1[27] <= Weights1[(32'd85+32'd1)*32'd19-1:32'd85*32'd19];
			WeightsStore2[0] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[1] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[2] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[3] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[4] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[5] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[6] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[7] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[8] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[9] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[10] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[11] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[12] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[13] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[14] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[15] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[16] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[17] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[18] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[19] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[20] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[21] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[22] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[23] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[24] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[25] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[26] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore2[27] <= Weights2[(32'd86+32'd1)*32'd19-1:32'd86*32'd19];
			WeightsStore3[0] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[1] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[2] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[3] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[4] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[5] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[6] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[7] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[8] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[9] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[10] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[11] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[12] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[13] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[14] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[15] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[16] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[17] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[18] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[19] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[20] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[21] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[22] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[23] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[24] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[25] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[26] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore3[27] <= Weights3[(32'd87+32'd1)*32'd19-1:32'd87*32'd19];
			WeightsStore4[0] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[1] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[2] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[3] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[4] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[5] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[6] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[7] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[8] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[9] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[10] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[11] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[12] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[13] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[14] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[15] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[16] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[17] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[18] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[19] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[20] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[21] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[22] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[23] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[24] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[25] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[26] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore4[27] <= Weights4[(32'd88+32'd1)*32'd19-1:32'd88*32'd19];
			WeightsStore5[0] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[1] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[2] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[3] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[4] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[5] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[6] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[7] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[8] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[9] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[10] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[11] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[12] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[13] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[14] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[15] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[16] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[17] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[18] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[19] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[20] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[21] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[22] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[23] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[24] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[25] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[26] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore5[27] <= Weights5[(32'd89+32'd1)*32'd19-1:32'd89*32'd19];
			WeightsStore6[0] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[1] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[2] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[3] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[4] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[5] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[6] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[7] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[8] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[9] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[10] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[11] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[12] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[13] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[14] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[15] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[16] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[17] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[18] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[19] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[20] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[21] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[22] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[23] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[24] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[25] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[26] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore6[27] <= Weights6[(32'd90+32'd1)*32'd19-1:32'd90*32'd19];
			WeightsStore7[0] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[1] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[2] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[3] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[4] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[5] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[6] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[7] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[8] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[9] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[10] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[11] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[12] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[13] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[14] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[15] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[16] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[17] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[18] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[19] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[20] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[21] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[22] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[23] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[24] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[25] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[26] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore7[27] <= Weights7[(32'd91+32'd1)*32'd19-1:32'd91*32'd19];
			WeightsStore8[0] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[1] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[2] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[3] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[4] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[5] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[6] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[7] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[8] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[9] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[10] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[11] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[12] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[13] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[14] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[15] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[16] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[17] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[18] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[19] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[20] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[21] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[22] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[23] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[24] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[25] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[26] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore8[27] <= Weights8[(32'd92+32'd1)*32'd19-1:32'd92*32'd19];
			WeightsStore9[0] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[1] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[2] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[3] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[4] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[5] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[6] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[7] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[8] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[9] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[10] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[11] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[12] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[13] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[14] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[15] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[16] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[17] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[18] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[19] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[20] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[21] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[22] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[23] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[24] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[25] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[26] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
			WeightsStore9[27] <= Weights9[(32'd93+32'd1)*32'd19-1:32'd93*32'd19];
		end else if(switchCounter == 32'd4)begin
			PixelsStore[0] <= Pixels[(32'd112+32'd1)*32'd10-1:32'd112*32'd10];
			PixelsStore[1] <= Pixels[(32'd113+32'd1)*32'd10-1:32'd113*32'd10];
			PixelsStore[2] <= Pixels[(32'd114+32'd1)*32'd10-1:32'd114*32'd10];
			PixelsStore[3] <= Pixels[(32'd115+32'd1)*32'd10-1:32'd115*32'd10];
			PixelsStore[4] <= Pixels[(32'd116+32'd1)*32'd10-1:32'd116*32'd10];
			PixelsStore[5] <= Pixels[(32'd117+32'd1)*32'd10-1:32'd117*32'd10];
			PixelsStore[6] <= Pixels[(32'd118+32'd1)*32'd10-1:32'd118*32'd10];
			PixelsStore[7] <= Pixels[(32'd119+32'd1)*32'd10-1:32'd119*32'd10];
			PixelsStore[8] <= Pixels[(32'd120+32'd1)*32'd10-1:32'd120*32'd10];
			PixelsStore[9] <= Pixels[(32'd121+32'd1)*32'd10-1:32'd121*32'd10];
			PixelsStore[10] <= Pixels[(32'd122+32'd1)*32'd10-1:32'd122*32'd10];
			PixelsStore[11] <= Pixels[(32'd123+32'd1)*32'd10-1:32'd123*32'd10];
			PixelsStore[12] <= Pixels[(32'd124+32'd1)*32'd10-1:32'd124*32'd10];
			PixelsStore[13] <= Pixels[(32'd125+32'd1)*32'd10-1:32'd125*32'd10];
			PixelsStore[14] <= Pixels[(32'd126+32'd1)*32'd10-1:32'd126*32'd10];
			PixelsStore[15] <= Pixels[(32'd127+32'd1)*32'd10-1:32'd127*32'd10];
			PixelsStore[16] <= Pixels[(32'd128+32'd1)*32'd10-1:32'd128*32'd10];
			PixelsStore[17] <= Pixels[(32'd129+32'd1)*32'd10-1:32'd129*32'd10];
			PixelsStore[18] <= Pixels[(32'd130+32'd1)*32'd10-1:32'd130*32'd10];
			PixelsStore[19] <= Pixels[(32'd131+32'd1)*32'd10-1:32'd131*32'd10];
			PixelsStore[20] <= Pixels[(32'd132+32'd1)*32'd10-1:32'd132*32'd10];
			PixelsStore[21] <= Pixels[(32'd133+32'd1)*32'd10-1:32'd133*32'd10];
			PixelsStore[22] <= Pixels[(32'd134+32'd1)*32'd10-1:32'd134*32'd10];
			PixelsStore[23] <= Pixels[(32'd135+32'd1)*32'd10-1:32'd135*32'd10];
			PixelsStore[24] <= Pixels[(32'd136+32'd1)*32'd10-1:32'd136*32'd10];
			PixelsStore[25] <= Pixels[(32'd137+32'd1)*32'd10-1:32'd137*32'd10];
			PixelsStore[26] <= Pixels[(32'd138+32'd1)*32'd10-1:32'd138*32'd10];
			PixelsStore[27] <= Pixels[(32'd139+32'd1)*32'd10-1:32'd139*32'd10];
			WeightsStore0[0] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[1] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[2] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[3] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[4] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[5] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[6] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[7] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[8] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[9] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[10] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[11] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[12] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[13] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[14] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[15] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[16] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[17] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[18] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[19] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[20] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[21] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[22] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[23] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[24] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[25] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[26] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore0[27] <= Weights0[(32'd112+32'd1)*32'd19-1:32'd112*32'd19];
			WeightsStore1[0] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[1] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[2] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[3] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[4] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[5] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[6] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[7] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[8] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[9] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[10] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[11] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[12] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[13] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[14] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[15] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[16] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[17] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[18] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[19] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[20] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[21] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[22] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[23] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[24] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[25] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[26] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore1[27] <= Weights1[(32'd113+32'd1)*32'd19-1:32'd113*32'd19];
			WeightsStore2[0] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[1] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[2] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[3] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[4] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[5] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[6] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[7] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[8] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[9] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[10] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[11] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[12] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[13] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[14] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[15] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[16] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[17] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[18] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[19] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[20] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[21] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[22] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[23] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[24] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[25] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[26] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore2[27] <= Weights2[(32'd114+32'd1)*32'd19-1:32'd114*32'd19];
			WeightsStore3[0] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[1] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[2] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[3] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[4] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[5] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[6] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[7] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[8] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[9] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[10] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[11] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[12] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[13] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[14] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[15] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[16] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[17] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[18] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[19] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[20] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[21] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[22] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[23] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[24] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[25] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[26] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore3[27] <= Weights3[(32'd115+32'd1)*32'd19-1:32'd115*32'd19];
			WeightsStore4[0] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[1] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[2] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[3] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[4] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[5] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[6] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[7] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[8] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[9] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[10] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[11] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[12] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[13] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[14] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[15] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[16] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[17] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[18] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[19] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[20] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[21] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[22] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[23] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[24] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[25] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[26] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore4[27] <= Weights4[(32'd116+32'd1)*32'd19-1:32'd116*32'd19];
			WeightsStore5[0] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[1] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[2] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[3] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[4] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[5] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[6] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[7] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[8] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[9] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[10] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[11] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[12] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[13] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[14] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[15] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[16] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[17] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[18] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[19] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[20] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[21] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[22] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[23] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[24] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[25] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[26] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore5[27] <= Weights5[(32'd117+32'd1)*32'd19-1:32'd117*32'd19];
			WeightsStore6[0] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[1] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[2] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[3] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[4] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[5] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[6] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[7] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[8] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[9] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[10] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[11] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[12] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[13] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[14] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[15] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[16] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[17] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[18] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[19] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[20] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[21] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[22] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[23] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[24] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[25] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[26] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore6[27] <= Weights6[(32'd118+32'd1)*32'd19-1:32'd118*32'd19];
			WeightsStore7[0] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[1] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[2] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[3] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[4] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[5] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[6] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[7] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[8] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[9] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[10] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[11] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[12] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[13] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[14] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[15] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[16] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[17] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[18] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[19] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[20] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[21] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[22] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[23] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[24] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[25] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[26] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore7[27] <= Weights7[(32'd119+32'd1)*32'd19-1:32'd119*32'd19];
			WeightsStore8[0] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[1] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[2] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[3] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[4] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[5] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[6] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[7] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[8] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[9] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[10] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[11] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[12] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[13] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[14] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[15] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[16] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[17] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[18] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[19] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[20] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[21] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[22] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[23] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[24] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[25] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[26] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore8[27] <= Weights8[(32'd120+32'd1)*32'd19-1:32'd120*32'd19];
			WeightsStore9[0] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[1] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[2] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[3] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[4] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[5] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[6] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[7] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[8] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[9] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[10] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[11] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[12] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[13] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[14] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[15] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[16] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[17] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[18] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[19] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[20] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[21] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[22] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[23] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[24] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[25] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[26] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
			WeightsStore9[27] <= Weights9[(32'd121+32'd1)*32'd19-1:32'd121*32'd19];
		end else if(switchCounter == 32'd5)begin
			PixelsStore[0] <= Pixels[(32'd140+32'd1)*32'd10-1:32'd140*32'd10];
			PixelsStore[1] <= Pixels[(32'd141+32'd1)*32'd10-1:32'd141*32'd10];
			PixelsStore[2] <= Pixels[(32'd142+32'd1)*32'd10-1:32'd142*32'd10];
			PixelsStore[3] <= Pixels[(32'd143+32'd1)*32'd10-1:32'd143*32'd10];
			PixelsStore[4] <= Pixels[(32'd144+32'd1)*32'd10-1:32'd144*32'd10];
			PixelsStore[5] <= Pixels[(32'd145+32'd1)*32'd10-1:32'd145*32'd10];
			PixelsStore[6] <= Pixels[(32'd146+32'd1)*32'd10-1:32'd146*32'd10];
			PixelsStore[7] <= Pixels[(32'd147+32'd1)*32'd10-1:32'd147*32'd10];
			PixelsStore[8] <= Pixels[(32'd148+32'd1)*32'd10-1:32'd148*32'd10];
			PixelsStore[9] <= Pixels[(32'd149+32'd1)*32'd10-1:32'd149*32'd10];
			PixelsStore[10] <= Pixels[(32'd150+32'd1)*32'd10-1:32'd150*32'd10];
			PixelsStore[11] <= Pixels[(32'd151+32'd1)*32'd10-1:32'd151*32'd10];
			PixelsStore[12] <= Pixels[(32'd152+32'd1)*32'd10-1:32'd152*32'd10];
			PixelsStore[13] <= Pixels[(32'd153+32'd1)*32'd10-1:32'd153*32'd10];
			PixelsStore[14] <= Pixels[(32'd154+32'd1)*32'd10-1:32'd154*32'd10];
			PixelsStore[15] <= Pixels[(32'd155+32'd1)*32'd10-1:32'd155*32'd10];
			PixelsStore[16] <= Pixels[(32'd156+32'd1)*32'd10-1:32'd156*32'd10];
			PixelsStore[17] <= Pixels[(32'd157+32'd1)*32'd10-1:32'd157*32'd10];
			PixelsStore[18] <= Pixels[(32'd158+32'd1)*32'd10-1:32'd158*32'd10];
			PixelsStore[19] <= Pixels[(32'd159+32'd1)*32'd10-1:32'd159*32'd10];
			PixelsStore[20] <= Pixels[(32'd160+32'd1)*32'd10-1:32'd160*32'd10];
			PixelsStore[21] <= Pixels[(32'd161+32'd1)*32'd10-1:32'd161*32'd10];
			PixelsStore[22] <= Pixels[(32'd162+32'd1)*32'd10-1:32'd162*32'd10];
			PixelsStore[23] <= Pixels[(32'd163+32'd1)*32'd10-1:32'd163*32'd10];
			PixelsStore[24] <= Pixels[(32'd164+32'd1)*32'd10-1:32'd164*32'd10];
			PixelsStore[25] <= Pixels[(32'd165+32'd1)*32'd10-1:32'd165*32'd10];
			PixelsStore[26] <= Pixels[(32'd166+32'd1)*32'd10-1:32'd166*32'd10];
			PixelsStore[27] <= Pixels[(32'd167+32'd1)*32'd10-1:32'd167*32'd10];
			WeightsStore0[0] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[1] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[2] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[3] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[4] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[5] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[6] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[7] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[8] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[9] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[10] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[11] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[12] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[13] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[14] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[15] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[16] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[17] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[18] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[19] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[20] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[21] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[22] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[23] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[24] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[25] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[26] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore0[27] <= Weights0[(32'd140+32'd1)*32'd19-1:32'd140*32'd19];
			WeightsStore1[0] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[1] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[2] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[3] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[4] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[5] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[6] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[7] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[8] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[9] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[10] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[11] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[12] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[13] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[14] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[15] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[16] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[17] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[18] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[19] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[20] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[21] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[22] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[23] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[24] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[25] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[26] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore1[27] <= Weights1[(32'd141+32'd1)*32'd19-1:32'd141*32'd19];
			WeightsStore2[0] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[1] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[2] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[3] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[4] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[5] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[6] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[7] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[8] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[9] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[10] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[11] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[12] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[13] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[14] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[15] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[16] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[17] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[18] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[19] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[20] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[21] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[22] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[23] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[24] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[25] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[26] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore2[27] <= Weights2[(32'd142+32'd1)*32'd19-1:32'd142*32'd19];
			WeightsStore3[0] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[1] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[2] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[3] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[4] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[5] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[6] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[7] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[8] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[9] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[10] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[11] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[12] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[13] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[14] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[15] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[16] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[17] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[18] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[19] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[20] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[21] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[22] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[23] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[24] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[25] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[26] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore3[27] <= Weights3[(32'd143+32'd1)*32'd19-1:32'd143*32'd19];
			WeightsStore4[0] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[1] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[2] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[3] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[4] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[5] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[6] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[7] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[8] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[9] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[10] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[11] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[12] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[13] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[14] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[15] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[16] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[17] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[18] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[19] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[20] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[21] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[22] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[23] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[24] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[25] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[26] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore4[27] <= Weights4[(32'd144+32'd1)*32'd19-1:32'd144*32'd19];
			WeightsStore5[0] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[1] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[2] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[3] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[4] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[5] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[6] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[7] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[8] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[9] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[10] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[11] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[12] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[13] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[14] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[15] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[16] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[17] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[18] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[19] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[20] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[21] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[22] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[23] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[24] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[25] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[26] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore5[27] <= Weights5[(32'd145+32'd1)*32'd19-1:32'd145*32'd19];
			WeightsStore6[0] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[1] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[2] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[3] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[4] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[5] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[6] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[7] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[8] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[9] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[10] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[11] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[12] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[13] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[14] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[15] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[16] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[17] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[18] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[19] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[20] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[21] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[22] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[23] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[24] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[25] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[26] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore6[27] <= Weights6[(32'd146+32'd1)*32'd19-1:32'd146*32'd19];
			WeightsStore7[0] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[1] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[2] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[3] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[4] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[5] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[6] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[7] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[8] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[9] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[10] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[11] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[12] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[13] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[14] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[15] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[16] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[17] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[18] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[19] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[20] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[21] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[22] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[23] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[24] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[25] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[26] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore7[27] <= Weights7[(32'd147+32'd1)*32'd19-1:32'd147*32'd19];
			WeightsStore8[0] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[1] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[2] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[3] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[4] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[5] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[6] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[7] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[8] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[9] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[10] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[11] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[12] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[13] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[14] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[15] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[16] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[17] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[18] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[19] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[20] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[21] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[22] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[23] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[24] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[25] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[26] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore8[27] <= Weights8[(32'd148+32'd1)*32'd19-1:32'd148*32'd19];
			WeightsStore9[0] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[1] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[2] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[3] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[4] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[5] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[6] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[7] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[8] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[9] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[10] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[11] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[12] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[13] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[14] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[15] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[16] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[17] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[18] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[19] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[20] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[21] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[22] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[23] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[24] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[25] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[26] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
			WeightsStore9[27] <= Weights9[(32'd149+32'd1)*32'd19-1:32'd149*32'd19];
		end else if(switchCounter == 32'd6)begin
			PixelsStore[0] <= Pixels[(32'd168+32'd1)*32'd10-1:32'd168*32'd10];
			PixelsStore[1] <= Pixels[(32'd169+32'd1)*32'd10-1:32'd169*32'd10];
			PixelsStore[2] <= Pixels[(32'd170+32'd1)*32'd10-1:32'd170*32'd10];
			PixelsStore[3] <= Pixels[(32'd171+32'd1)*32'd10-1:32'd171*32'd10];
			PixelsStore[4] <= Pixels[(32'd172+32'd1)*32'd10-1:32'd172*32'd10];
			PixelsStore[5] <= Pixels[(32'd173+32'd1)*32'd10-1:32'd173*32'd10];
			PixelsStore[6] <= Pixels[(32'd174+32'd1)*32'd10-1:32'd174*32'd10];
			PixelsStore[7] <= Pixels[(32'd175+32'd1)*32'd10-1:32'd175*32'd10];
			PixelsStore[8] <= Pixels[(32'd176+32'd1)*32'd10-1:32'd176*32'd10];
			PixelsStore[9] <= Pixels[(32'd177+32'd1)*32'd10-1:32'd177*32'd10];
			PixelsStore[10] <= Pixels[(32'd178+32'd1)*32'd10-1:32'd178*32'd10];
			PixelsStore[11] <= Pixels[(32'd179+32'd1)*32'd10-1:32'd179*32'd10];
			PixelsStore[12] <= Pixels[(32'd180+32'd1)*32'd10-1:32'd180*32'd10];
			PixelsStore[13] <= Pixels[(32'd181+32'd1)*32'd10-1:32'd181*32'd10];
			PixelsStore[14] <= Pixels[(32'd182+32'd1)*32'd10-1:32'd182*32'd10];
			PixelsStore[15] <= Pixels[(32'd183+32'd1)*32'd10-1:32'd183*32'd10];
			PixelsStore[16] <= Pixels[(32'd184+32'd1)*32'd10-1:32'd184*32'd10];
			PixelsStore[17] <= Pixels[(32'd185+32'd1)*32'd10-1:32'd185*32'd10];
			PixelsStore[18] <= Pixels[(32'd186+32'd1)*32'd10-1:32'd186*32'd10];
			PixelsStore[19] <= Pixels[(32'd187+32'd1)*32'd10-1:32'd187*32'd10];
			PixelsStore[20] <= Pixels[(32'd188+32'd1)*32'd10-1:32'd188*32'd10];
			PixelsStore[21] <= Pixels[(32'd189+32'd1)*32'd10-1:32'd189*32'd10];
			PixelsStore[22] <= Pixels[(32'd190+32'd1)*32'd10-1:32'd190*32'd10];
			PixelsStore[23] <= Pixels[(32'd191+32'd1)*32'd10-1:32'd191*32'd10];
			PixelsStore[24] <= Pixels[(32'd192+32'd1)*32'd10-1:32'd192*32'd10];
			PixelsStore[25] <= Pixels[(32'd193+32'd1)*32'd10-1:32'd193*32'd10];
			PixelsStore[26] <= Pixels[(32'd194+32'd1)*32'd10-1:32'd194*32'd10];
			PixelsStore[27] <= Pixels[(32'd195+32'd1)*32'd10-1:32'd195*32'd10];
			WeightsStore0[0] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[1] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[2] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[3] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[4] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[5] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[6] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[7] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[8] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[9] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[10] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[11] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[12] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[13] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[14] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[15] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[16] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[17] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[18] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[19] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[20] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[21] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[22] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[23] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[24] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[25] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[26] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore0[27] <= Weights0[(32'd168+32'd1)*32'd19-1:32'd168*32'd19];
			WeightsStore1[0] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[1] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[2] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[3] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[4] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[5] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[6] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[7] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[8] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[9] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[10] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[11] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[12] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[13] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[14] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[15] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[16] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[17] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[18] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[19] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[20] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[21] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[22] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[23] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[24] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[25] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[26] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore1[27] <= Weights1[(32'd169+32'd1)*32'd19-1:32'd169*32'd19];
			WeightsStore2[0] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[1] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[2] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[3] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[4] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[5] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[6] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[7] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[8] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[9] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[10] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[11] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[12] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[13] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[14] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[15] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[16] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[17] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[18] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[19] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[20] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[21] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[22] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[23] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[24] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[25] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[26] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore2[27] <= Weights2[(32'd170+32'd1)*32'd19-1:32'd170*32'd19];
			WeightsStore3[0] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[1] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[2] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[3] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[4] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[5] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[6] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[7] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[8] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[9] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[10] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[11] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[12] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[13] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[14] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[15] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[16] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[17] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[18] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[19] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[20] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[21] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[22] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[23] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[24] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[25] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[26] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore3[27] <= Weights3[(32'd171+32'd1)*32'd19-1:32'd171*32'd19];
			WeightsStore4[0] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[1] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[2] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[3] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[4] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[5] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[6] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[7] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[8] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[9] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[10] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[11] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[12] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[13] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[14] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[15] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[16] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[17] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[18] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[19] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[20] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[21] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[22] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[23] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[24] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[25] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[26] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore4[27] <= Weights4[(32'd172+32'd1)*32'd19-1:32'd172*32'd19];
			WeightsStore5[0] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[1] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[2] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[3] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[4] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[5] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[6] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[7] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[8] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[9] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[10] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[11] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[12] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[13] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[14] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[15] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[16] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[17] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[18] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[19] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[20] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[21] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[22] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[23] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[24] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[25] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[26] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore5[27] <= Weights5[(32'd173+32'd1)*32'd19-1:32'd173*32'd19];
			WeightsStore6[0] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[1] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[2] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[3] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[4] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[5] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[6] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[7] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[8] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[9] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[10] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[11] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[12] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[13] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[14] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[15] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[16] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[17] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[18] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[19] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[20] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[21] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[22] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[23] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[24] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[25] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[26] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore6[27] <= Weights6[(32'd174+32'd1)*32'd19-1:32'd174*32'd19];
			WeightsStore7[0] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[1] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[2] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[3] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[4] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[5] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[6] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[7] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[8] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[9] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[10] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[11] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[12] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[13] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[14] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[15] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[16] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[17] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[18] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[19] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[20] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[21] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[22] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[23] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[24] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[25] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[26] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore7[27] <= Weights7[(32'd175+32'd1)*32'd19-1:32'd175*32'd19];
			WeightsStore8[0] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[1] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[2] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[3] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[4] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[5] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[6] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[7] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[8] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[9] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[10] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[11] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[12] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[13] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[14] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[15] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[16] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[17] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[18] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[19] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[20] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[21] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[22] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[23] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[24] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[25] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[26] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore8[27] <= Weights8[(32'd176+32'd1)*32'd19-1:32'd176*32'd19];
			WeightsStore9[0] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[1] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[2] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[3] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[4] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[5] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[6] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[7] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[8] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[9] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[10] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[11] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[12] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[13] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[14] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[15] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[16] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[17] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[18] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[19] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[20] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[21] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[22] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[23] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[24] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[25] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[26] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
			WeightsStore9[27] <= Weights9[(32'd177+32'd1)*32'd19-1:32'd177*32'd19];
		end else if(switchCounter == 32'd7)begin
			PixelsStore[0] <= Pixels[(32'd196+32'd1)*32'd10-1:32'd196*32'd10];
			PixelsStore[1] <= Pixels[(32'd197+32'd1)*32'd10-1:32'd197*32'd10];
			PixelsStore[2] <= Pixels[(32'd198+32'd1)*32'd10-1:32'd198*32'd10];
			PixelsStore[3] <= Pixels[(32'd199+32'd1)*32'd10-1:32'd199*32'd10];
			PixelsStore[4] <= Pixels[(32'd200+32'd1)*32'd10-1:32'd200*32'd10];
			PixelsStore[5] <= Pixels[(32'd201+32'd1)*32'd10-1:32'd201*32'd10];
			PixelsStore[6] <= Pixels[(32'd202+32'd1)*32'd10-1:32'd202*32'd10];
			PixelsStore[7] <= Pixels[(32'd203+32'd1)*32'd10-1:32'd203*32'd10];
			PixelsStore[8] <= Pixels[(32'd204+32'd1)*32'd10-1:32'd204*32'd10];
			PixelsStore[9] <= Pixels[(32'd205+32'd1)*32'd10-1:32'd205*32'd10];
			PixelsStore[10] <= Pixels[(32'd206+32'd1)*32'd10-1:32'd206*32'd10];
			PixelsStore[11] <= Pixels[(32'd207+32'd1)*32'd10-1:32'd207*32'd10];
			PixelsStore[12] <= Pixels[(32'd208+32'd1)*32'd10-1:32'd208*32'd10];
			PixelsStore[13] <= Pixels[(32'd209+32'd1)*32'd10-1:32'd209*32'd10];
			PixelsStore[14] <= Pixels[(32'd210+32'd1)*32'd10-1:32'd210*32'd10];
			PixelsStore[15] <= Pixels[(32'd211+32'd1)*32'd10-1:32'd211*32'd10];
			PixelsStore[16] <= Pixels[(32'd212+32'd1)*32'd10-1:32'd212*32'd10];
			PixelsStore[17] <= Pixels[(32'd213+32'd1)*32'd10-1:32'd213*32'd10];
			PixelsStore[18] <= Pixels[(32'd214+32'd1)*32'd10-1:32'd214*32'd10];
			PixelsStore[19] <= Pixels[(32'd215+32'd1)*32'd10-1:32'd215*32'd10];
			PixelsStore[20] <= Pixels[(32'd216+32'd1)*32'd10-1:32'd216*32'd10];
			PixelsStore[21] <= Pixels[(32'd217+32'd1)*32'd10-1:32'd217*32'd10];
			PixelsStore[22] <= Pixels[(32'd218+32'd1)*32'd10-1:32'd218*32'd10];
			PixelsStore[23] <= Pixels[(32'd219+32'd1)*32'd10-1:32'd219*32'd10];
			PixelsStore[24] <= Pixels[(32'd220+32'd1)*32'd10-1:32'd220*32'd10];
			PixelsStore[25] <= Pixels[(32'd221+32'd1)*32'd10-1:32'd221*32'd10];
			PixelsStore[26] <= Pixels[(32'd222+32'd1)*32'd10-1:32'd222*32'd10];
			PixelsStore[27] <= Pixels[(32'd223+32'd1)*32'd10-1:32'd223*32'd10];
			WeightsStore0[0] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[1] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[2] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[3] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[4] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[5] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[6] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[7] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[8] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[9] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[10] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[11] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[12] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[13] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[14] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[15] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[16] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[17] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[18] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[19] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[20] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[21] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[22] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[23] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[24] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[25] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[26] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore0[27] <= Weights0[(32'd196+32'd1)*32'd19-1:32'd196*32'd19];
			WeightsStore1[0] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[1] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[2] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[3] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[4] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[5] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[6] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[7] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[8] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[9] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[10] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[11] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[12] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[13] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[14] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[15] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[16] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[17] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[18] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[19] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[20] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[21] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[22] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[23] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[24] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[25] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[26] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore1[27] <= Weights1[(32'd197+32'd1)*32'd19-1:32'd197*32'd19];
			WeightsStore2[0] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[1] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[2] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[3] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[4] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[5] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[6] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[7] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[8] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[9] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[10] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[11] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[12] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[13] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[14] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[15] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[16] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[17] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[18] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[19] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[20] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[21] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[22] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[23] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[24] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[25] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[26] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore2[27] <= Weights2[(32'd198+32'd1)*32'd19-1:32'd198*32'd19];
			WeightsStore3[0] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[1] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[2] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[3] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[4] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[5] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[6] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[7] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[8] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[9] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[10] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[11] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[12] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[13] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[14] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[15] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[16] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[17] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[18] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[19] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[20] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[21] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[22] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[23] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[24] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[25] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[26] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore3[27] <= Weights3[(32'd199+32'd1)*32'd19-1:32'd199*32'd19];
			WeightsStore4[0] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[1] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[2] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[3] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[4] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[5] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[6] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[7] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[8] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[9] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[10] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[11] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[12] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[13] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[14] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[15] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[16] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[17] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[18] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[19] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[20] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[21] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[22] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[23] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[24] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[25] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[26] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore4[27] <= Weights4[(32'd200+32'd1)*32'd19-1:32'd200*32'd19];
			WeightsStore5[0] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[1] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[2] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[3] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[4] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[5] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[6] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[7] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[8] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[9] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[10] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[11] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[12] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[13] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[14] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[15] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[16] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[17] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[18] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[19] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[20] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[21] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[22] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[23] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[24] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[25] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[26] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore5[27] <= Weights5[(32'd201+32'd1)*32'd19-1:32'd201*32'd19];
			WeightsStore6[0] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[1] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[2] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[3] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[4] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[5] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[6] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[7] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[8] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[9] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[10] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[11] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[12] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[13] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[14] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[15] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[16] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[17] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[18] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[19] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[20] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[21] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[22] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[23] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[24] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[25] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[26] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore6[27] <= Weights6[(32'd202+32'd1)*32'd19-1:32'd202*32'd19];
			WeightsStore7[0] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[1] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[2] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[3] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[4] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[5] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[6] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[7] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[8] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[9] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[10] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[11] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[12] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[13] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[14] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[15] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[16] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[17] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[18] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[19] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[20] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[21] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[22] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[23] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[24] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[25] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[26] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore7[27] <= Weights7[(32'd203+32'd1)*32'd19-1:32'd203*32'd19];
			WeightsStore8[0] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[1] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[2] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[3] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[4] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[5] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[6] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[7] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[8] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[9] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[10] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[11] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[12] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[13] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[14] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[15] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[16] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[17] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[18] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[19] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[20] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[21] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[22] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[23] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[24] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[25] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[26] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore8[27] <= Weights8[(32'd204+32'd1)*32'd19-1:32'd204*32'd19];
			WeightsStore9[0] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[1] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[2] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[3] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[4] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[5] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[6] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[7] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[8] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[9] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[10] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[11] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[12] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[13] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[14] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[15] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[16] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[17] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[18] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[19] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[20] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[21] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[22] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[23] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[24] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[25] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[26] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
			WeightsStore9[27] <= Weights9[(32'd205+32'd1)*32'd19-1:32'd205*32'd19];
		end else if(switchCounter == 32'd8)begin
			PixelsStore[0] <= Pixels[(32'd224+32'd1)*32'd10-1:32'd224*32'd10];
			PixelsStore[1] <= Pixels[(32'd225+32'd1)*32'd10-1:32'd225*32'd10];
			PixelsStore[2] <= Pixels[(32'd226+32'd1)*32'd10-1:32'd226*32'd10];
			PixelsStore[3] <= Pixels[(32'd227+32'd1)*32'd10-1:32'd227*32'd10];
			PixelsStore[4] <= Pixels[(32'd228+32'd1)*32'd10-1:32'd228*32'd10];
			PixelsStore[5] <= Pixels[(32'd229+32'd1)*32'd10-1:32'd229*32'd10];
			PixelsStore[6] <= Pixels[(32'd230+32'd1)*32'd10-1:32'd230*32'd10];
			PixelsStore[7] <= Pixels[(32'd231+32'd1)*32'd10-1:32'd231*32'd10];
			PixelsStore[8] <= Pixels[(32'd232+32'd1)*32'd10-1:32'd232*32'd10];
			PixelsStore[9] <= Pixels[(32'd233+32'd1)*32'd10-1:32'd233*32'd10];
			PixelsStore[10] <= Pixels[(32'd234+32'd1)*32'd10-1:32'd234*32'd10];
			PixelsStore[11] <= Pixels[(32'd235+32'd1)*32'd10-1:32'd235*32'd10];
			PixelsStore[12] <= Pixels[(32'd236+32'd1)*32'd10-1:32'd236*32'd10];
			PixelsStore[13] <= Pixels[(32'd237+32'd1)*32'd10-1:32'd237*32'd10];
			PixelsStore[14] <= Pixels[(32'd238+32'd1)*32'd10-1:32'd238*32'd10];
			PixelsStore[15] <= Pixels[(32'd239+32'd1)*32'd10-1:32'd239*32'd10];
			PixelsStore[16] <= Pixels[(32'd240+32'd1)*32'd10-1:32'd240*32'd10];
			PixelsStore[17] <= Pixels[(32'd241+32'd1)*32'd10-1:32'd241*32'd10];
			PixelsStore[18] <= Pixels[(32'd242+32'd1)*32'd10-1:32'd242*32'd10];
			PixelsStore[19] <= Pixels[(32'd243+32'd1)*32'd10-1:32'd243*32'd10];
			PixelsStore[20] <= Pixels[(32'd244+32'd1)*32'd10-1:32'd244*32'd10];
			PixelsStore[21] <= Pixels[(32'd245+32'd1)*32'd10-1:32'd245*32'd10];
			PixelsStore[22] <= Pixels[(32'd246+32'd1)*32'd10-1:32'd246*32'd10];
			PixelsStore[23] <= Pixels[(32'd247+32'd1)*32'd10-1:32'd247*32'd10];
			PixelsStore[24] <= Pixels[(32'd248+32'd1)*32'd10-1:32'd248*32'd10];
			PixelsStore[25] <= Pixels[(32'd249+32'd1)*32'd10-1:32'd249*32'd10];
			PixelsStore[26] <= Pixels[(32'd250+32'd1)*32'd10-1:32'd250*32'd10];
			PixelsStore[27] <= Pixels[(32'd251+32'd1)*32'd10-1:32'd251*32'd10];
			WeightsStore0[0] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[1] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[2] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[3] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[4] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[5] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[6] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[7] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[8] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[9] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[10] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[11] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[12] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[13] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[14] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[15] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[16] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[17] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[18] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[19] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[20] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[21] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[22] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[23] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[24] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[25] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[26] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore0[27] <= Weights0[(32'd224+32'd1)*32'd19-1:32'd224*32'd19];
			WeightsStore1[0] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[1] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[2] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[3] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[4] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[5] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[6] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[7] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[8] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[9] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[10] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[11] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[12] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[13] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[14] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[15] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[16] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[17] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[18] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[19] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[20] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[21] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[22] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[23] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[24] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[25] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[26] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore1[27] <= Weights1[(32'd225+32'd1)*32'd19-1:32'd225*32'd19];
			WeightsStore2[0] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[1] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[2] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[3] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[4] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[5] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[6] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[7] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[8] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[9] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[10] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[11] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[12] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[13] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[14] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[15] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[16] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[17] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[18] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[19] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[20] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[21] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[22] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[23] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[24] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[25] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[26] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore2[27] <= Weights2[(32'd226+32'd1)*32'd19-1:32'd226*32'd19];
			WeightsStore3[0] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[1] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[2] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[3] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[4] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[5] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[6] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[7] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[8] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[9] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[10] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[11] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[12] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[13] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[14] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[15] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[16] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[17] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[18] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[19] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[20] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[21] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[22] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[23] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[24] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[25] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[26] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore3[27] <= Weights3[(32'd227+32'd1)*32'd19-1:32'd227*32'd19];
			WeightsStore4[0] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[1] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[2] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[3] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[4] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[5] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[6] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[7] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[8] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[9] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[10] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[11] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[12] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[13] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[14] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[15] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[16] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[17] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[18] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[19] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[20] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[21] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[22] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[23] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[24] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[25] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[26] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore4[27] <= Weights4[(32'd228+32'd1)*32'd19-1:32'd228*32'd19];
			WeightsStore5[0] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[1] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[2] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[3] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[4] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[5] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[6] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[7] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[8] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[9] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[10] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[11] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[12] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[13] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[14] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[15] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[16] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[17] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[18] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[19] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[20] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[21] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[22] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[23] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[24] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[25] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[26] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore5[27] <= Weights5[(32'd229+32'd1)*32'd19-1:32'd229*32'd19];
			WeightsStore6[0] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[1] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[2] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[3] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[4] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[5] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[6] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[7] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[8] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[9] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[10] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[11] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[12] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[13] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[14] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[15] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[16] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[17] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[18] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[19] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[20] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[21] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[22] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[23] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[24] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[25] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[26] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore6[27] <= Weights6[(32'd230+32'd1)*32'd19-1:32'd230*32'd19];
			WeightsStore7[0] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[1] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[2] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[3] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[4] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[5] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[6] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[7] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[8] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[9] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[10] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[11] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[12] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[13] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[14] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[15] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[16] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[17] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[18] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[19] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[20] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[21] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[22] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[23] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[24] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[25] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[26] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore7[27] <= Weights7[(32'd231+32'd1)*32'd19-1:32'd231*32'd19];
			WeightsStore8[0] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[1] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[2] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[3] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[4] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[5] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[6] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[7] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[8] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[9] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[10] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[11] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[12] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[13] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[14] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[15] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[16] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[17] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[18] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[19] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[20] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[21] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[22] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[23] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[24] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[25] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[26] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore8[27] <= Weights8[(32'd232+32'd1)*32'd19-1:32'd232*32'd19];
			WeightsStore9[0] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[1] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[2] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[3] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[4] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[5] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[6] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[7] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[8] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[9] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[10] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[11] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[12] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[13] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[14] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[15] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[16] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[17] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[18] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[19] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[20] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[21] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[22] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[23] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[24] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[25] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[26] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
			WeightsStore9[27] <= Weights9[(32'd233+32'd1)*32'd19-1:32'd233*32'd19];
		end else if(switchCounter == 32'd9)begin
			PixelsStore[0] <= Pixels[(32'd252+32'd1)*32'd10-1:32'd252*32'd10];
			PixelsStore[1] <= Pixels[(32'd253+32'd1)*32'd10-1:32'd253*32'd10];
			PixelsStore[2] <= Pixels[(32'd254+32'd1)*32'd10-1:32'd254*32'd10];
			PixelsStore[3] <= Pixels[(32'd255+32'd1)*32'd10-1:32'd255*32'd10];
			PixelsStore[4] <= Pixels[(32'd256+32'd1)*32'd10-1:32'd256*32'd10];
			PixelsStore[5] <= Pixels[(32'd257+32'd1)*32'd10-1:32'd257*32'd10];
			PixelsStore[6] <= Pixels[(32'd258+32'd1)*32'd10-1:32'd258*32'd10];
			PixelsStore[7] <= Pixels[(32'd259+32'd1)*32'd10-1:32'd259*32'd10];
			PixelsStore[8] <= Pixels[(32'd260+32'd1)*32'd10-1:32'd260*32'd10];
			PixelsStore[9] <= Pixels[(32'd261+32'd1)*32'd10-1:32'd261*32'd10];
			PixelsStore[10] <= Pixels[(32'd262+32'd1)*32'd10-1:32'd262*32'd10];
			PixelsStore[11] <= Pixels[(32'd263+32'd1)*32'd10-1:32'd263*32'd10];
			PixelsStore[12] <= Pixels[(32'd264+32'd1)*32'd10-1:32'd264*32'd10];
			PixelsStore[13] <= Pixels[(32'd265+32'd1)*32'd10-1:32'd265*32'd10];
			PixelsStore[14] <= Pixels[(32'd266+32'd1)*32'd10-1:32'd266*32'd10];
			PixelsStore[15] <= Pixels[(32'd267+32'd1)*32'd10-1:32'd267*32'd10];
			PixelsStore[16] <= Pixels[(32'd268+32'd1)*32'd10-1:32'd268*32'd10];
			PixelsStore[17] <= Pixels[(32'd269+32'd1)*32'd10-1:32'd269*32'd10];
			PixelsStore[18] <= Pixels[(32'd270+32'd1)*32'd10-1:32'd270*32'd10];
			PixelsStore[19] <= Pixels[(32'd271+32'd1)*32'd10-1:32'd271*32'd10];
			PixelsStore[20] <= Pixels[(32'd272+32'd1)*32'd10-1:32'd272*32'd10];
			PixelsStore[21] <= Pixels[(32'd273+32'd1)*32'd10-1:32'd273*32'd10];
			PixelsStore[22] <= Pixels[(32'd274+32'd1)*32'd10-1:32'd274*32'd10];
			PixelsStore[23] <= Pixels[(32'd275+32'd1)*32'd10-1:32'd275*32'd10];
			PixelsStore[24] <= Pixels[(32'd276+32'd1)*32'd10-1:32'd276*32'd10];
			PixelsStore[25] <= Pixels[(32'd277+32'd1)*32'd10-1:32'd277*32'd10];
			PixelsStore[26] <= Pixels[(32'd278+32'd1)*32'd10-1:32'd278*32'd10];
			PixelsStore[27] <= Pixels[(32'd279+32'd1)*32'd10-1:32'd279*32'd10];
			WeightsStore0[0] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[1] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[2] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[3] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[4] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[5] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[6] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[7] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[8] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[9] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[10] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[11] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[12] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[13] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[14] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[15] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[16] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[17] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[18] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[19] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[20] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[21] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[22] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[23] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[24] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[25] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[26] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore0[27] <= Weights0[(32'd252+32'd1)*32'd19-1:32'd252*32'd19];
			WeightsStore1[0] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[1] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[2] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[3] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[4] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[5] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[6] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[7] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[8] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[9] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[10] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[11] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[12] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[13] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[14] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[15] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[16] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[17] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[18] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[19] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[20] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[21] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[22] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[23] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[24] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[25] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[26] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore1[27] <= Weights1[(32'd253+32'd1)*32'd19-1:32'd253*32'd19];
			WeightsStore2[0] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[1] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[2] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[3] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[4] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[5] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[6] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[7] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[8] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[9] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[10] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[11] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[12] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[13] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[14] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[15] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[16] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[17] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[18] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[19] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[20] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[21] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[22] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[23] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[24] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[25] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[26] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore2[27] <= Weights2[(32'd254+32'd1)*32'd19-1:32'd254*32'd19];
			WeightsStore3[0] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[1] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[2] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[3] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[4] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[5] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[6] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[7] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[8] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[9] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[10] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[11] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[12] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[13] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[14] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[15] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[16] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[17] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[18] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[19] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[20] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[21] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[22] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[23] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[24] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[25] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[26] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore3[27] <= Weights3[(32'd255+32'd1)*32'd19-1:32'd255*32'd19];
			WeightsStore4[0] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[1] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[2] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[3] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[4] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[5] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[6] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[7] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[8] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[9] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[10] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[11] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[12] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[13] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[14] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[15] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[16] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[17] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[18] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[19] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[20] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[21] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[22] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[23] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[24] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[25] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[26] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore4[27] <= Weights4[(32'd256+32'd1)*32'd19-1:32'd256*32'd19];
			WeightsStore5[0] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[1] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[2] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[3] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[4] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[5] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[6] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[7] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[8] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[9] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[10] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[11] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[12] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[13] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[14] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[15] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[16] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[17] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[18] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[19] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[20] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[21] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[22] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[23] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[24] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[25] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[26] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore5[27] <= Weights5[(32'd257+32'd1)*32'd19-1:32'd257*32'd19];
			WeightsStore6[0] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[1] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[2] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[3] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[4] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[5] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[6] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[7] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[8] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[9] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[10] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[11] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[12] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[13] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[14] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[15] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[16] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[17] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[18] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[19] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[20] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[21] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[22] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[23] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[24] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[25] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[26] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore6[27] <= Weights6[(32'd258+32'd1)*32'd19-1:32'd258*32'd19];
			WeightsStore7[0] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[1] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[2] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[3] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[4] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[5] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[6] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[7] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[8] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[9] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[10] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[11] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[12] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[13] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[14] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[15] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[16] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[17] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[18] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[19] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[20] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[21] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[22] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[23] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[24] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[25] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[26] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore7[27] <= Weights7[(32'd259+32'd1)*32'd19-1:32'd259*32'd19];
			WeightsStore8[0] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[1] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[2] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[3] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[4] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[5] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[6] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[7] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[8] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[9] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[10] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[11] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[12] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[13] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[14] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[15] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[16] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[17] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[18] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[19] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[20] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[21] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[22] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[23] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[24] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[25] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[26] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore8[27] <= Weights8[(32'd260+32'd1)*32'd19-1:32'd260*32'd19];
			WeightsStore9[0] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[1] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[2] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[3] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[4] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[5] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[6] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[7] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[8] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[9] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[10] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[11] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[12] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[13] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[14] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[15] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[16] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[17] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[18] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[19] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[20] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[21] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[22] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[23] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[24] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[25] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[26] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
			WeightsStore9[27] <= Weights9[(32'd261+32'd1)*32'd19-1:32'd261*32'd19];
		end else if(switchCounter == 32'd10)begin
			PixelsStore[0] <= Pixels[(32'd280+32'd1)*32'd10-1:32'd280*32'd10];
			PixelsStore[1] <= Pixels[(32'd281+32'd1)*32'd10-1:32'd281*32'd10];
			PixelsStore[2] <= Pixels[(32'd282+32'd1)*32'd10-1:32'd282*32'd10];
			PixelsStore[3] <= Pixels[(32'd283+32'd1)*32'd10-1:32'd283*32'd10];
			PixelsStore[4] <= Pixels[(32'd284+32'd1)*32'd10-1:32'd284*32'd10];
			PixelsStore[5] <= Pixels[(32'd285+32'd1)*32'd10-1:32'd285*32'd10];
			PixelsStore[6] <= Pixels[(32'd286+32'd1)*32'd10-1:32'd286*32'd10];
			PixelsStore[7] <= Pixels[(32'd287+32'd1)*32'd10-1:32'd287*32'd10];
			PixelsStore[8] <= Pixels[(32'd288+32'd1)*32'd10-1:32'd288*32'd10];
			PixelsStore[9] <= Pixels[(32'd289+32'd1)*32'd10-1:32'd289*32'd10];
			PixelsStore[10] <= Pixels[(32'd290+32'd1)*32'd10-1:32'd290*32'd10];
			PixelsStore[11] <= Pixels[(32'd291+32'd1)*32'd10-1:32'd291*32'd10];
			PixelsStore[12] <= Pixels[(32'd292+32'd1)*32'd10-1:32'd292*32'd10];
			PixelsStore[13] <= Pixels[(32'd293+32'd1)*32'd10-1:32'd293*32'd10];
			PixelsStore[14] <= Pixels[(32'd294+32'd1)*32'd10-1:32'd294*32'd10];
			PixelsStore[15] <= Pixels[(32'd295+32'd1)*32'd10-1:32'd295*32'd10];
			PixelsStore[16] <= Pixels[(32'd296+32'd1)*32'd10-1:32'd296*32'd10];
			PixelsStore[17] <= Pixels[(32'd297+32'd1)*32'd10-1:32'd297*32'd10];
			PixelsStore[18] <= Pixels[(32'd298+32'd1)*32'd10-1:32'd298*32'd10];
			PixelsStore[19] <= Pixels[(32'd299+32'd1)*32'd10-1:32'd299*32'd10];
			PixelsStore[20] <= Pixels[(32'd300+32'd1)*32'd10-1:32'd300*32'd10];
			PixelsStore[21] <= Pixels[(32'd301+32'd1)*32'd10-1:32'd301*32'd10];
			PixelsStore[22] <= Pixels[(32'd302+32'd1)*32'd10-1:32'd302*32'd10];
			PixelsStore[23] <= Pixels[(32'd303+32'd1)*32'd10-1:32'd303*32'd10];
			PixelsStore[24] <= Pixels[(32'd304+32'd1)*32'd10-1:32'd304*32'd10];
			PixelsStore[25] <= Pixels[(32'd305+32'd1)*32'd10-1:32'd305*32'd10];
			PixelsStore[26] <= Pixels[(32'd306+32'd1)*32'd10-1:32'd306*32'd10];
			PixelsStore[27] <= Pixels[(32'd307+32'd1)*32'd10-1:32'd307*32'd10];
			WeightsStore0[0] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[1] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[2] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[3] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[4] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[5] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[6] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[7] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[8] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[9] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[10] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[11] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[12] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[13] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[14] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[15] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[16] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[17] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[18] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[19] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[20] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[21] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[22] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[23] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[24] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[25] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[26] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore0[27] <= Weights0[(32'd280+32'd1)*32'd19-1:32'd280*32'd19];
			WeightsStore1[0] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[1] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[2] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[3] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[4] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[5] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[6] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[7] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[8] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[9] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[10] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[11] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[12] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[13] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[14] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[15] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[16] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[17] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[18] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[19] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[20] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[21] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[22] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[23] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[24] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[25] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[26] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore1[27] <= Weights1[(32'd281+32'd1)*32'd19-1:32'd281*32'd19];
			WeightsStore2[0] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[1] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[2] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[3] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[4] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[5] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[6] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[7] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[8] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[9] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[10] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[11] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[12] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[13] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[14] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[15] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[16] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[17] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[18] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[19] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[20] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[21] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[22] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[23] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[24] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[25] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[26] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore2[27] <= Weights2[(32'd282+32'd1)*32'd19-1:32'd282*32'd19];
			WeightsStore3[0] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[1] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[2] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[3] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[4] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[5] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[6] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[7] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[8] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[9] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[10] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[11] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[12] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[13] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[14] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[15] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[16] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[17] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[18] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[19] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[20] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[21] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[22] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[23] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[24] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[25] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[26] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore3[27] <= Weights3[(32'd283+32'd1)*32'd19-1:32'd283*32'd19];
			WeightsStore4[0] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[1] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[2] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[3] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[4] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[5] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[6] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[7] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[8] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[9] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[10] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[11] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[12] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[13] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[14] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[15] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[16] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[17] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[18] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[19] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[20] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[21] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[22] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[23] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[24] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[25] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[26] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore4[27] <= Weights4[(32'd284+32'd1)*32'd19-1:32'd284*32'd19];
			WeightsStore5[0] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[1] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[2] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[3] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[4] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[5] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[6] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[7] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[8] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[9] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[10] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[11] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[12] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[13] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[14] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[15] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[16] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[17] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[18] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[19] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[20] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[21] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[22] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[23] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[24] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[25] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[26] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore5[27] <= Weights5[(32'd285+32'd1)*32'd19-1:32'd285*32'd19];
			WeightsStore6[0] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[1] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[2] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[3] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[4] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[5] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[6] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[7] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[8] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[9] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[10] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[11] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[12] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[13] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[14] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[15] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[16] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[17] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[18] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[19] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[20] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[21] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[22] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[23] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[24] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[25] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[26] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore6[27] <= Weights6[(32'd286+32'd1)*32'd19-1:32'd286*32'd19];
			WeightsStore7[0] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[1] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[2] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[3] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[4] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[5] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[6] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[7] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[8] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[9] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[10] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[11] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[12] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[13] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[14] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[15] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[16] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[17] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[18] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[19] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[20] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[21] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[22] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[23] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[24] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[25] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[26] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore7[27] <= Weights7[(32'd287+32'd1)*32'd19-1:32'd287*32'd19];
			WeightsStore8[0] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[1] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[2] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[3] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[4] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[5] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[6] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[7] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[8] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[9] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[10] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[11] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[12] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[13] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[14] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[15] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[16] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[17] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[18] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[19] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[20] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[21] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[22] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[23] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[24] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[25] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[26] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore8[27] <= Weights8[(32'd288+32'd1)*32'd19-1:32'd288*32'd19];
			WeightsStore9[0] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[1] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[2] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[3] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[4] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[5] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[6] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[7] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[8] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[9] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[10] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[11] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[12] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[13] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[14] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[15] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[16] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[17] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[18] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[19] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[20] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[21] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[22] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[23] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[24] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[25] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[26] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
			WeightsStore9[27] <= Weights9[(32'd289+32'd1)*32'd19-1:32'd289*32'd19];
		end else if(switchCounter == 32'd11)begin
			PixelsStore[0] <= Pixels[(32'd308+32'd1)*32'd10-1:32'd308*32'd10];
			PixelsStore[1] <= Pixels[(32'd309+32'd1)*32'd10-1:32'd309*32'd10];
			PixelsStore[2] <= Pixels[(32'd310+32'd1)*32'd10-1:32'd310*32'd10];
			PixelsStore[3] <= Pixels[(32'd311+32'd1)*32'd10-1:32'd311*32'd10];
			PixelsStore[4] <= Pixels[(32'd312+32'd1)*32'd10-1:32'd312*32'd10];
			PixelsStore[5] <= Pixels[(32'd313+32'd1)*32'd10-1:32'd313*32'd10];
			PixelsStore[6] <= Pixels[(32'd314+32'd1)*32'd10-1:32'd314*32'd10];
			PixelsStore[7] <= Pixels[(32'd315+32'd1)*32'd10-1:32'd315*32'd10];
			PixelsStore[8] <= Pixels[(32'd316+32'd1)*32'd10-1:32'd316*32'd10];
			PixelsStore[9] <= Pixels[(32'd317+32'd1)*32'd10-1:32'd317*32'd10];
			PixelsStore[10] <= Pixels[(32'd318+32'd1)*32'd10-1:32'd318*32'd10];
			PixelsStore[11] <= Pixels[(32'd319+32'd1)*32'd10-1:32'd319*32'd10];
			PixelsStore[12] <= Pixels[(32'd320+32'd1)*32'd10-1:32'd320*32'd10];
			PixelsStore[13] <= Pixels[(32'd321+32'd1)*32'd10-1:32'd321*32'd10];
			PixelsStore[14] <= Pixels[(32'd322+32'd1)*32'd10-1:32'd322*32'd10];
			PixelsStore[15] <= Pixels[(32'd323+32'd1)*32'd10-1:32'd323*32'd10];
			PixelsStore[16] <= Pixels[(32'd324+32'd1)*32'd10-1:32'd324*32'd10];
			PixelsStore[17] <= Pixels[(32'd325+32'd1)*32'd10-1:32'd325*32'd10];
			PixelsStore[18] <= Pixels[(32'd326+32'd1)*32'd10-1:32'd326*32'd10];
			PixelsStore[19] <= Pixels[(32'd327+32'd1)*32'd10-1:32'd327*32'd10];
			PixelsStore[20] <= Pixels[(32'd328+32'd1)*32'd10-1:32'd328*32'd10];
			PixelsStore[21] <= Pixels[(32'd329+32'd1)*32'd10-1:32'd329*32'd10];
			PixelsStore[22] <= Pixels[(32'd330+32'd1)*32'd10-1:32'd330*32'd10];
			PixelsStore[23] <= Pixels[(32'd331+32'd1)*32'd10-1:32'd331*32'd10];
			PixelsStore[24] <= Pixels[(32'd332+32'd1)*32'd10-1:32'd332*32'd10];
			PixelsStore[25] <= Pixels[(32'd333+32'd1)*32'd10-1:32'd333*32'd10];
			PixelsStore[26] <= Pixels[(32'd334+32'd1)*32'd10-1:32'd334*32'd10];
			PixelsStore[27] <= Pixels[(32'd335+32'd1)*32'd10-1:32'd335*32'd10];
			WeightsStore0[0] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[1] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[2] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[3] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[4] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[5] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[6] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[7] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[8] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[9] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[10] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[11] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[12] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[13] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[14] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[15] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[16] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[17] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[18] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[19] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[20] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[21] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[22] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[23] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[24] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[25] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[26] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore0[27] <= Weights0[(32'd308+32'd1)*32'd19-1:32'd308*32'd19];
			WeightsStore1[0] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[1] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[2] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[3] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[4] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[5] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[6] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[7] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[8] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[9] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[10] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[11] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[12] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[13] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[14] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[15] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[16] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[17] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[18] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[19] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[20] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[21] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[22] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[23] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[24] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[25] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[26] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore1[27] <= Weights1[(32'd309+32'd1)*32'd19-1:32'd309*32'd19];
			WeightsStore2[0] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[1] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[2] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[3] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[4] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[5] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[6] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[7] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[8] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[9] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[10] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[11] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[12] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[13] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[14] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[15] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[16] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[17] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[18] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[19] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[20] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[21] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[22] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[23] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[24] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[25] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[26] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore2[27] <= Weights2[(32'd310+32'd1)*32'd19-1:32'd310*32'd19];
			WeightsStore3[0] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[1] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[2] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[3] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[4] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[5] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[6] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[7] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[8] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[9] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[10] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[11] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[12] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[13] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[14] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[15] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[16] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[17] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[18] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[19] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[20] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[21] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[22] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[23] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[24] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[25] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[26] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore3[27] <= Weights3[(32'd311+32'd1)*32'd19-1:32'd311*32'd19];
			WeightsStore4[0] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[1] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[2] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[3] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[4] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[5] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[6] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[7] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[8] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[9] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[10] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[11] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[12] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[13] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[14] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[15] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[16] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[17] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[18] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[19] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[20] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[21] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[22] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[23] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[24] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[25] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[26] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore4[27] <= Weights4[(32'd312+32'd1)*32'd19-1:32'd312*32'd19];
			WeightsStore5[0] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[1] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[2] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[3] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[4] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[5] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[6] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[7] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[8] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[9] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[10] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[11] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[12] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[13] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[14] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[15] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[16] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[17] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[18] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[19] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[20] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[21] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[22] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[23] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[24] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[25] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[26] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore5[27] <= Weights5[(32'd313+32'd1)*32'd19-1:32'd313*32'd19];
			WeightsStore6[0] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[1] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[2] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[3] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[4] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[5] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[6] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[7] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[8] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[9] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[10] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[11] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[12] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[13] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[14] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[15] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[16] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[17] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[18] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[19] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[20] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[21] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[22] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[23] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[24] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[25] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[26] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore6[27] <= Weights6[(32'd314+32'd1)*32'd19-1:32'd314*32'd19];
			WeightsStore7[0] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[1] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[2] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[3] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[4] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[5] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[6] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[7] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[8] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[9] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[10] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[11] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[12] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[13] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[14] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[15] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[16] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[17] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[18] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[19] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[20] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[21] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[22] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[23] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[24] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[25] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[26] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore7[27] <= Weights7[(32'd315+32'd1)*32'd19-1:32'd315*32'd19];
			WeightsStore8[0] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[1] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[2] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[3] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[4] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[5] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[6] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[7] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[8] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[9] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[10] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[11] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[12] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[13] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[14] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[15] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[16] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[17] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[18] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[19] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[20] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[21] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[22] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[23] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[24] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[25] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[26] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore8[27] <= Weights8[(32'd316+32'd1)*32'd19-1:32'd316*32'd19];
			WeightsStore9[0] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[1] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[2] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[3] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[4] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[5] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[6] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[7] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[8] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[9] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[10] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[11] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[12] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[13] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[14] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[15] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[16] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[17] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[18] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[19] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[20] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[21] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[22] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[23] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[24] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[25] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[26] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
			WeightsStore9[27] <= Weights9[(32'd317+32'd1)*32'd19-1:32'd317*32'd19];
		end else if(switchCounter == 32'd12)begin
			PixelsStore[0] <= Pixels[(32'd336+32'd1)*32'd10-1:32'd336*32'd10];
			PixelsStore[1] <= Pixels[(32'd337+32'd1)*32'd10-1:32'd337*32'd10];
			PixelsStore[2] <= Pixels[(32'd338+32'd1)*32'd10-1:32'd338*32'd10];
			PixelsStore[3] <= Pixels[(32'd339+32'd1)*32'd10-1:32'd339*32'd10];
			PixelsStore[4] <= Pixels[(32'd340+32'd1)*32'd10-1:32'd340*32'd10];
			PixelsStore[5] <= Pixels[(32'd341+32'd1)*32'd10-1:32'd341*32'd10];
			PixelsStore[6] <= Pixels[(32'd342+32'd1)*32'd10-1:32'd342*32'd10];
			PixelsStore[7] <= Pixels[(32'd343+32'd1)*32'd10-1:32'd343*32'd10];
			PixelsStore[8] <= Pixels[(32'd344+32'd1)*32'd10-1:32'd344*32'd10];
			PixelsStore[9] <= Pixels[(32'd345+32'd1)*32'd10-1:32'd345*32'd10];
			PixelsStore[10] <= Pixels[(32'd346+32'd1)*32'd10-1:32'd346*32'd10];
			PixelsStore[11] <= Pixels[(32'd347+32'd1)*32'd10-1:32'd347*32'd10];
			PixelsStore[12] <= Pixels[(32'd348+32'd1)*32'd10-1:32'd348*32'd10];
			PixelsStore[13] <= Pixels[(32'd349+32'd1)*32'd10-1:32'd349*32'd10];
			PixelsStore[14] <= Pixels[(32'd350+32'd1)*32'd10-1:32'd350*32'd10];
			PixelsStore[15] <= Pixels[(32'd351+32'd1)*32'd10-1:32'd351*32'd10];
			PixelsStore[16] <= Pixels[(32'd352+32'd1)*32'd10-1:32'd352*32'd10];
			PixelsStore[17] <= Pixels[(32'd353+32'd1)*32'd10-1:32'd353*32'd10];
			PixelsStore[18] <= Pixels[(32'd354+32'd1)*32'd10-1:32'd354*32'd10];
			PixelsStore[19] <= Pixels[(32'd355+32'd1)*32'd10-1:32'd355*32'd10];
			PixelsStore[20] <= Pixels[(32'd356+32'd1)*32'd10-1:32'd356*32'd10];
			PixelsStore[21] <= Pixels[(32'd357+32'd1)*32'd10-1:32'd357*32'd10];
			PixelsStore[22] <= Pixels[(32'd358+32'd1)*32'd10-1:32'd358*32'd10];
			PixelsStore[23] <= Pixels[(32'd359+32'd1)*32'd10-1:32'd359*32'd10];
			PixelsStore[24] <= Pixels[(32'd360+32'd1)*32'd10-1:32'd360*32'd10];
			PixelsStore[25] <= Pixels[(32'd361+32'd1)*32'd10-1:32'd361*32'd10];
			PixelsStore[26] <= Pixels[(32'd362+32'd1)*32'd10-1:32'd362*32'd10];
			PixelsStore[27] <= Pixels[(32'd363+32'd1)*32'd10-1:32'd363*32'd10];
			WeightsStore0[0] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[1] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[2] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[3] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[4] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[5] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[6] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[7] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[8] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[9] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[10] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[11] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[12] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[13] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[14] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[15] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[16] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[17] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[18] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[19] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[20] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[21] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[22] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[23] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[24] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[25] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[26] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore0[27] <= Weights0[(32'd336+32'd1)*32'd19-1:32'd336*32'd19];
			WeightsStore1[0] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[1] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[2] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[3] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[4] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[5] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[6] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[7] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[8] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[9] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[10] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[11] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[12] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[13] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[14] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[15] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[16] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[17] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[18] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[19] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[20] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[21] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[22] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[23] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[24] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[25] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[26] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore1[27] <= Weights1[(32'd337+32'd1)*32'd19-1:32'd337*32'd19];
			WeightsStore2[0] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[1] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[2] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[3] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[4] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[5] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[6] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[7] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[8] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[9] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[10] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[11] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[12] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[13] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[14] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[15] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[16] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[17] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[18] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[19] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[20] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[21] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[22] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[23] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[24] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[25] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[26] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore2[27] <= Weights2[(32'd338+32'd1)*32'd19-1:32'd338*32'd19];
			WeightsStore3[0] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[1] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[2] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[3] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[4] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[5] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[6] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[7] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[8] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[9] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[10] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[11] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[12] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[13] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[14] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[15] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[16] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[17] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[18] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[19] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[20] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[21] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[22] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[23] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[24] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[25] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[26] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore3[27] <= Weights3[(32'd339+32'd1)*32'd19-1:32'd339*32'd19];
			WeightsStore4[0] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[1] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[2] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[3] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[4] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[5] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[6] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[7] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[8] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[9] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[10] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[11] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[12] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[13] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[14] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[15] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[16] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[17] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[18] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[19] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[20] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[21] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[22] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[23] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[24] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[25] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[26] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore4[27] <= Weights4[(32'd340+32'd1)*32'd19-1:32'd340*32'd19];
			WeightsStore5[0] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[1] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[2] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[3] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[4] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[5] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[6] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[7] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[8] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[9] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[10] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[11] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[12] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[13] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[14] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[15] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[16] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[17] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[18] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[19] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[20] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[21] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[22] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[23] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[24] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[25] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[26] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore5[27] <= Weights5[(32'd341+32'd1)*32'd19-1:32'd341*32'd19];
			WeightsStore6[0] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[1] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[2] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[3] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[4] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[5] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[6] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[7] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[8] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[9] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[10] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[11] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[12] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[13] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[14] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[15] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[16] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[17] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[18] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[19] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[20] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[21] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[22] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[23] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[24] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[25] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[26] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore6[27] <= Weights6[(32'd342+32'd1)*32'd19-1:32'd342*32'd19];
			WeightsStore7[0] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[1] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[2] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[3] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[4] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[5] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[6] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[7] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[8] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[9] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[10] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[11] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[12] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[13] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[14] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[15] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[16] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[17] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[18] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[19] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[20] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[21] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[22] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[23] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[24] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[25] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[26] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore7[27] <= Weights7[(32'd343+32'd1)*32'd19-1:32'd343*32'd19];
			WeightsStore8[0] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[1] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[2] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[3] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[4] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[5] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[6] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[7] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[8] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[9] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[10] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[11] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[12] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[13] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[14] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[15] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[16] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[17] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[18] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[19] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[20] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[21] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[22] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[23] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[24] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[25] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[26] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore8[27] <= Weights8[(32'd344+32'd1)*32'd19-1:32'd344*32'd19];
			WeightsStore9[0] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[1] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[2] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[3] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[4] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[5] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[6] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[7] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[8] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[9] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[10] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[11] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[12] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[13] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[14] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[15] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[16] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[17] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[18] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[19] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[20] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[21] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[22] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[23] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[24] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[25] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[26] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
			WeightsStore9[27] <= Weights9[(32'd345+32'd1)*32'd19-1:32'd345*32'd19];
		end else if(switchCounter == 32'd13)begin
			PixelsStore[0] <= Pixels[(32'd364+32'd1)*32'd10-1:32'd364*32'd10];
			PixelsStore[1] <= Pixels[(32'd365+32'd1)*32'd10-1:32'd365*32'd10];
			PixelsStore[2] <= Pixels[(32'd366+32'd1)*32'd10-1:32'd366*32'd10];
			PixelsStore[3] <= Pixels[(32'd367+32'd1)*32'd10-1:32'd367*32'd10];
			PixelsStore[4] <= Pixels[(32'd368+32'd1)*32'd10-1:32'd368*32'd10];
			PixelsStore[5] <= Pixels[(32'd369+32'd1)*32'd10-1:32'd369*32'd10];
			PixelsStore[6] <= Pixels[(32'd370+32'd1)*32'd10-1:32'd370*32'd10];
			PixelsStore[7] <= Pixels[(32'd371+32'd1)*32'd10-1:32'd371*32'd10];
			PixelsStore[8] <= Pixels[(32'd372+32'd1)*32'd10-1:32'd372*32'd10];
			PixelsStore[9] <= Pixels[(32'd373+32'd1)*32'd10-1:32'd373*32'd10];
			PixelsStore[10] <= Pixels[(32'd374+32'd1)*32'd10-1:32'd374*32'd10];
			PixelsStore[11] <= Pixels[(32'd375+32'd1)*32'd10-1:32'd375*32'd10];
			PixelsStore[12] <= Pixels[(32'd376+32'd1)*32'd10-1:32'd376*32'd10];
			PixelsStore[13] <= Pixels[(32'd377+32'd1)*32'd10-1:32'd377*32'd10];
			PixelsStore[14] <= Pixels[(32'd378+32'd1)*32'd10-1:32'd378*32'd10];
			PixelsStore[15] <= Pixels[(32'd379+32'd1)*32'd10-1:32'd379*32'd10];
			PixelsStore[16] <= Pixels[(32'd380+32'd1)*32'd10-1:32'd380*32'd10];
			PixelsStore[17] <= Pixels[(32'd381+32'd1)*32'd10-1:32'd381*32'd10];
			PixelsStore[18] <= Pixels[(32'd382+32'd1)*32'd10-1:32'd382*32'd10];
			PixelsStore[19] <= Pixels[(32'd383+32'd1)*32'd10-1:32'd383*32'd10];
			PixelsStore[20] <= Pixels[(32'd384+32'd1)*32'd10-1:32'd384*32'd10];
			PixelsStore[21] <= Pixels[(32'd385+32'd1)*32'd10-1:32'd385*32'd10];
			PixelsStore[22] <= Pixels[(32'd386+32'd1)*32'd10-1:32'd386*32'd10];
			PixelsStore[23] <= Pixels[(32'd387+32'd1)*32'd10-1:32'd387*32'd10];
			PixelsStore[24] <= Pixels[(32'd388+32'd1)*32'd10-1:32'd388*32'd10];
			PixelsStore[25] <= Pixels[(32'd389+32'd1)*32'd10-1:32'd389*32'd10];
			PixelsStore[26] <= Pixels[(32'd390+32'd1)*32'd10-1:32'd390*32'd10];
			PixelsStore[27] <= Pixels[(32'd391+32'd1)*32'd10-1:32'd391*32'd10];
			WeightsStore0[0] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[1] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[2] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[3] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[4] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[5] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[6] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[7] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[8] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[9] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[10] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[11] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[12] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[13] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[14] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[15] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[16] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[17] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[18] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[19] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[20] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[21] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[22] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[23] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[24] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[25] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[26] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore0[27] <= Weights0[(32'd364+32'd1)*32'd19-1:32'd364*32'd19];
			WeightsStore1[0] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[1] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[2] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[3] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[4] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[5] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[6] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[7] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[8] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[9] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[10] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[11] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[12] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[13] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[14] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[15] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[16] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[17] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[18] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[19] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[20] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[21] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[22] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[23] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[24] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[25] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[26] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore1[27] <= Weights1[(32'd365+32'd1)*32'd19-1:32'd365*32'd19];
			WeightsStore2[0] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[1] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[2] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[3] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[4] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[5] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[6] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[7] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[8] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[9] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[10] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[11] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[12] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[13] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[14] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[15] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[16] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[17] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[18] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[19] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[20] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[21] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[22] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[23] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[24] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[25] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[26] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore2[27] <= Weights2[(32'd366+32'd1)*32'd19-1:32'd366*32'd19];
			WeightsStore3[0] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[1] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[2] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[3] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[4] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[5] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[6] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[7] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[8] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[9] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[10] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[11] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[12] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[13] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[14] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[15] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[16] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[17] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[18] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[19] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[20] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[21] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[22] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[23] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[24] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[25] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[26] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore3[27] <= Weights3[(32'd367+32'd1)*32'd19-1:32'd367*32'd19];
			WeightsStore4[0] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[1] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[2] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[3] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[4] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[5] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[6] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[7] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[8] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[9] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[10] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[11] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[12] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[13] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[14] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[15] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[16] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[17] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[18] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[19] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[20] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[21] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[22] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[23] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[24] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[25] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[26] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore4[27] <= Weights4[(32'd368+32'd1)*32'd19-1:32'd368*32'd19];
			WeightsStore5[0] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[1] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[2] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[3] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[4] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[5] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[6] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[7] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[8] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[9] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[10] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[11] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[12] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[13] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[14] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[15] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[16] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[17] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[18] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[19] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[20] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[21] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[22] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[23] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[24] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[25] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[26] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore5[27] <= Weights5[(32'd369+32'd1)*32'd19-1:32'd369*32'd19];
			WeightsStore6[0] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[1] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[2] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[3] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[4] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[5] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[6] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[7] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[8] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[9] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[10] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[11] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[12] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[13] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[14] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[15] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[16] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[17] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[18] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[19] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[20] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[21] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[22] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[23] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[24] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[25] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[26] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore6[27] <= Weights6[(32'd370+32'd1)*32'd19-1:32'd370*32'd19];
			WeightsStore7[0] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[1] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[2] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[3] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[4] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[5] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[6] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[7] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[8] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[9] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[10] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[11] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[12] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[13] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[14] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[15] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[16] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[17] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[18] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[19] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[20] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[21] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[22] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[23] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[24] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[25] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[26] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore7[27] <= Weights7[(32'd371+32'd1)*32'd19-1:32'd371*32'd19];
			WeightsStore8[0] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[1] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[2] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[3] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[4] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[5] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[6] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[7] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[8] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[9] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[10] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[11] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[12] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[13] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[14] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[15] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[16] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[17] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[18] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[19] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[20] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[21] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[22] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[23] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[24] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[25] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[26] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore8[27] <= Weights8[(32'd372+32'd1)*32'd19-1:32'd372*32'd19];
			WeightsStore9[0] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[1] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[2] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[3] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[4] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[5] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[6] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[7] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[8] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[9] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[10] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[11] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[12] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[13] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[14] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[15] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[16] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[17] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[18] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[19] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[20] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[21] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[22] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[23] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[24] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[25] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[26] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
			WeightsStore9[27] <= Weights9[(32'd373+32'd1)*32'd19-1:32'd373*32'd19];
		end else if(switchCounter == 32'd14)begin
			PixelsStore[0] <= Pixels[(32'd392+32'd1)*32'd10-1:32'd392*32'd10];
			PixelsStore[1] <= Pixels[(32'd393+32'd1)*32'd10-1:32'd393*32'd10];
			PixelsStore[2] <= Pixels[(32'd394+32'd1)*32'd10-1:32'd394*32'd10];
			PixelsStore[3] <= Pixels[(32'd395+32'd1)*32'd10-1:32'd395*32'd10];
			PixelsStore[4] <= Pixels[(32'd396+32'd1)*32'd10-1:32'd396*32'd10];
			PixelsStore[5] <= Pixels[(32'd397+32'd1)*32'd10-1:32'd397*32'd10];
			PixelsStore[6] <= Pixels[(32'd398+32'd1)*32'd10-1:32'd398*32'd10];
			PixelsStore[7] <= Pixels[(32'd399+32'd1)*32'd10-1:32'd399*32'd10];
			PixelsStore[8] <= Pixels[(32'd400+32'd1)*32'd10-1:32'd400*32'd10];
			PixelsStore[9] <= Pixels[(32'd401+32'd1)*32'd10-1:32'd401*32'd10];
			PixelsStore[10] <= Pixels[(32'd402+32'd1)*32'd10-1:32'd402*32'd10];
			PixelsStore[11] <= Pixels[(32'd403+32'd1)*32'd10-1:32'd403*32'd10];
			PixelsStore[12] <= Pixels[(32'd404+32'd1)*32'd10-1:32'd404*32'd10];
			PixelsStore[13] <= Pixels[(32'd405+32'd1)*32'd10-1:32'd405*32'd10];
			PixelsStore[14] <= Pixels[(32'd406+32'd1)*32'd10-1:32'd406*32'd10];
			PixelsStore[15] <= Pixels[(32'd407+32'd1)*32'd10-1:32'd407*32'd10];
			PixelsStore[16] <= Pixels[(32'd408+32'd1)*32'd10-1:32'd408*32'd10];
			PixelsStore[17] <= Pixels[(32'd409+32'd1)*32'd10-1:32'd409*32'd10];
			PixelsStore[18] <= Pixels[(32'd410+32'd1)*32'd10-1:32'd410*32'd10];
			PixelsStore[19] <= Pixels[(32'd411+32'd1)*32'd10-1:32'd411*32'd10];
			PixelsStore[20] <= Pixels[(32'd412+32'd1)*32'd10-1:32'd412*32'd10];
			PixelsStore[21] <= Pixels[(32'd413+32'd1)*32'd10-1:32'd413*32'd10];
			PixelsStore[22] <= Pixels[(32'd414+32'd1)*32'd10-1:32'd414*32'd10];
			PixelsStore[23] <= Pixels[(32'd415+32'd1)*32'd10-1:32'd415*32'd10];
			PixelsStore[24] <= Pixels[(32'd416+32'd1)*32'd10-1:32'd416*32'd10];
			PixelsStore[25] <= Pixels[(32'd417+32'd1)*32'd10-1:32'd417*32'd10];
			PixelsStore[26] <= Pixels[(32'd418+32'd1)*32'd10-1:32'd418*32'd10];
			PixelsStore[27] <= Pixels[(32'd419+32'd1)*32'd10-1:32'd419*32'd10];
			WeightsStore0[0] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[1] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[2] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[3] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[4] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[5] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[6] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[7] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[8] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[9] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[10] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[11] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[12] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[13] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[14] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[15] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[16] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[17] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[18] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[19] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[20] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[21] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[22] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[23] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[24] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[25] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[26] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore0[27] <= Weights0[(32'd392+32'd1)*32'd19-1:32'd392*32'd19];
			WeightsStore1[0] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[1] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[2] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[3] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[4] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[5] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[6] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[7] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[8] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[9] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[10] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[11] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[12] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[13] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[14] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[15] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[16] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[17] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[18] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[19] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[20] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[21] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[22] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[23] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[24] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[25] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[26] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore1[27] <= Weights1[(32'd393+32'd1)*32'd19-1:32'd393*32'd19];
			WeightsStore2[0] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[1] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[2] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[3] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[4] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[5] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[6] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[7] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[8] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[9] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[10] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[11] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[12] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[13] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[14] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[15] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[16] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[17] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[18] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[19] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[20] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[21] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[22] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[23] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[24] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[25] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[26] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore2[27] <= Weights2[(32'd394+32'd1)*32'd19-1:32'd394*32'd19];
			WeightsStore3[0] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[1] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[2] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[3] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[4] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[5] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[6] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[7] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[8] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[9] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[10] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[11] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[12] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[13] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[14] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[15] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[16] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[17] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[18] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[19] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[20] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[21] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[22] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[23] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[24] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[25] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[26] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore3[27] <= Weights3[(32'd395+32'd1)*32'd19-1:32'd395*32'd19];
			WeightsStore4[0] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[1] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[2] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[3] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[4] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[5] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[6] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[7] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[8] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[9] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[10] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[11] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[12] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[13] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[14] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[15] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[16] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[17] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[18] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[19] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[20] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[21] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[22] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[23] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[24] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[25] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[26] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore4[27] <= Weights4[(32'd396+32'd1)*32'd19-1:32'd396*32'd19];
			WeightsStore5[0] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[1] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[2] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[3] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[4] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[5] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[6] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[7] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[8] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[9] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[10] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[11] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[12] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[13] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[14] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[15] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[16] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[17] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[18] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[19] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[20] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[21] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[22] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[23] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[24] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[25] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[26] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore5[27] <= Weights5[(32'd397+32'd1)*32'd19-1:32'd397*32'd19];
			WeightsStore6[0] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[1] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[2] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[3] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[4] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[5] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[6] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[7] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[8] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[9] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[10] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[11] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[12] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[13] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[14] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[15] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[16] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[17] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[18] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[19] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[20] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[21] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[22] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[23] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[24] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[25] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[26] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore6[27] <= Weights6[(32'd398+32'd1)*32'd19-1:32'd398*32'd19];
			WeightsStore7[0] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[1] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[2] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[3] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[4] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[5] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[6] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[7] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[8] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[9] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[10] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[11] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[12] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[13] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[14] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[15] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[16] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[17] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[18] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[19] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[20] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[21] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[22] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[23] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[24] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[25] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[26] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore7[27] <= Weights7[(32'd399+32'd1)*32'd19-1:32'd399*32'd19];
			WeightsStore8[0] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[1] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[2] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[3] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[4] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[5] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[6] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[7] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[8] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[9] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[10] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[11] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[12] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[13] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[14] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[15] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[16] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[17] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[18] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[19] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[20] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[21] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[22] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[23] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[24] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[25] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[26] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore8[27] <= Weights8[(32'd400+32'd1)*32'd19-1:32'd400*32'd19];
			WeightsStore9[0] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[1] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[2] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[3] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[4] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[5] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[6] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[7] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[8] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[9] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[10] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[11] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[12] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[13] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[14] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[15] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[16] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[17] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[18] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[19] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[20] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[21] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[22] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[23] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[24] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[25] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[26] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
			WeightsStore9[27] <= Weights9[(32'd401+32'd1)*32'd19-1:32'd401*32'd19];
		end else if(switchCounter == 32'd15)begin
			PixelsStore[0] <= Pixels[(32'd420+32'd1)*32'd10-1:32'd420*32'd10];
			PixelsStore[1] <= Pixels[(32'd421+32'd1)*32'd10-1:32'd421*32'd10];
			PixelsStore[2] <= Pixels[(32'd422+32'd1)*32'd10-1:32'd422*32'd10];
			PixelsStore[3] <= Pixels[(32'd423+32'd1)*32'd10-1:32'd423*32'd10];
			PixelsStore[4] <= Pixels[(32'd424+32'd1)*32'd10-1:32'd424*32'd10];
			PixelsStore[5] <= Pixels[(32'd425+32'd1)*32'd10-1:32'd425*32'd10];
			PixelsStore[6] <= Pixels[(32'd426+32'd1)*32'd10-1:32'd426*32'd10];
			PixelsStore[7] <= Pixels[(32'd427+32'd1)*32'd10-1:32'd427*32'd10];
			PixelsStore[8] <= Pixels[(32'd428+32'd1)*32'd10-1:32'd428*32'd10];
			PixelsStore[9] <= Pixels[(32'd429+32'd1)*32'd10-1:32'd429*32'd10];
			PixelsStore[10] <= Pixels[(32'd430+32'd1)*32'd10-1:32'd430*32'd10];
			PixelsStore[11] <= Pixels[(32'd431+32'd1)*32'd10-1:32'd431*32'd10];
			PixelsStore[12] <= Pixels[(32'd432+32'd1)*32'd10-1:32'd432*32'd10];
			PixelsStore[13] <= Pixels[(32'd433+32'd1)*32'd10-1:32'd433*32'd10];
			PixelsStore[14] <= Pixels[(32'd434+32'd1)*32'd10-1:32'd434*32'd10];
			PixelsStore[15] <= Pixels[(32'd435+32'd1)*32'd10-1:32'd435*32'd10];
			PixelsStore[16] <= Pixels[(32'd436+32'd1)*32'd10-1:32'd436*32'd10];
			PixelsStore[17] <= Pixels[(32'd437+32'd1)*32'd10-1:32'd437*32'd10];
			PixelsStore[18] <= Pixels[(32'd438+32'd1)*32'd10-1:32'd438*32'd10];
			PixelsStore[19] <= Pixels[(32'd439+32'd1)*32'd10-1:32'd439*32'd10];
			PixelsStore[20] <= Pixels[(32'd440+32'd1)*32'd10-1:32'd440*32'd10];
			PixelsStore[21] <= Pixels[(32'd441+32'd1)*32'd10-1:32'd441*32'd10];
			PixelsStore[22] <= Pixels[(32'd442+32'd1)*32'd10-1:32'd442*32'd10];
			PixelsStore[23] <= Pixels[(32'd443+32'd1)*32'd10-1:32'd443*32'd10];
			PixelsStore[24] <= Pixels[(32'd444+32'd1)*32'd10-1:32'd444*32'd10];
			PixelsStore[25] <= Pixels[(32'd445+32'd1)*32'd10-1:32'd445*32'd10];
			PixelsStore[26] <= Pixels[(32'd446+32'd1)*32'd10-1:32'd446*32'd10];
			PixelsStore[27] <= Pixels[(32'd447+32'd1)*32'd10-1:32'd447*32'd10];
			WeightsStore0[0] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[1] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[2] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[3] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[4] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[5] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[6] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[7] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[8] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[9] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[10] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[11] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[12] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[13] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[14] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[15] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[16] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[17] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[18] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[19] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[20] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[21] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[22] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[23] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[24] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[25] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[26] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore0[27] <= Weights0[(32'd420+32'd1)*32'd19-1:32'd420*32'd19];
			WeightsStore1[0] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[1] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[2] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[3] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[4] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[5] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[6] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[7] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[8] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[9] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[10] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[11] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[12] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[13] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[14] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[15] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[16] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[17] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[18] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[19] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[20] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[21] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[22] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[23] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[24] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[25] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[26] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore1[27] <= Weights1[(32'd421+32'd1)*32'd19-1:32'd421*32'd19];
			WeightsStore2[0] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[1] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[2] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[3] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[4] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[5] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[6] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[7] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[8] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[9] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[10] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[11] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[12] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[13] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[14] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[15] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[16] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[17] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[18] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[19] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[20] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[21] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[22] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[23] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[24] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[25] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[26] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore2[27] <= Weights2[(32'd422+32'd1)*32'd19-1:32'd422*32'd19];
			WeightsStore3[0] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[1] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[2] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[3] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[4] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[5] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[6] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[7] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[8] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[9] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[10] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[11] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[12] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[13] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[14] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[15] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[16] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[17] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[18] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[19] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[20] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[21] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[22] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[23] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[24] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[25] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[26] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore3[27] <= Weights3[(32'd423+32'd1)*32'd19-1:32'd423*32'd19];
			WeightsStore4[0] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[1] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[2] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[3] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[4] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[5] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[6] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[7] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[8] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[9] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[10] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[11] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[12] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[13] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[14] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[15] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[16] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[17] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[18] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[19] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[20] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[21] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[22] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[23] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[24] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[25] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[26] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore4[27] <= Weights4[(32'd424+32'd1)*32'd19-1:32'd424*32'd19];
			WeightsStore5[0] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[1] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[2] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[3] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[4] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[5] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[6] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[7] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[8] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[9] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[10] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[11] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[12] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[13] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[14] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[15] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[16] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[17] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[18] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[19] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[20] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[21] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[22] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[23] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[24] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[25] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[26] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore5[27] <= Weights5[(32'd425+32'd1)*32'd19-1:32'd425*32'd19];
			WeightsStore6[0] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[1] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[2] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[3] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[4] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[5] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[6] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[7] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[8] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[9] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[10] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[11] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[12] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[13] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[14] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[15] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[16] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[17] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[18] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[19] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[20] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[21] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[22] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[23] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[24] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[25] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[26] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore6[27] <= Weights6[(32'd426+32'd1)*32'd19-1:32'd426*32'd19];
			WeightsStore7[0] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[1] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[2] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[3] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[4] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[5] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[6] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[7] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[8] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[9] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[10] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[11] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[12] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[13] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[14] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[15] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[16] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[17] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[18] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[19] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[20] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[21] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[22] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[23] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[24] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[25] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[26] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore7[27] <= Weights7[(32'd427+32'd1)*32'd19-1:32'd427*32'd19];
			WeightsStore8[0] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[1] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[2] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[3] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[4] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[5] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[6] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[7] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[8] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[9] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[10] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[11] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[12] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[13] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[14] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[15] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[16] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[17] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[18] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[19] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[20] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[21] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[22] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[23] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[24] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[25] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[26] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore8[27] <= Weights8[(32'd428+32'd1)*32'd19-1:32'd428*32'd19];
			WeightsStore9[0] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[1] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[2] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[3] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[4] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[5] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[6] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[7] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[8] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[9] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[10] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[11] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[12] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[13] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[14] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[15] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[16] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[17] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[18] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[19] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[20] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[21] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[22] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[23] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[24] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[25] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[26] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
			WeightsStore9[27] <= Weights9[(32'd429+32'd1)*32'd19-1:32'd429*32'd19];
		end else if(switchCounter == 32'd16)begin
			PixelsStore[0] <= Pixels[(32'd448+32'd1)*32'd10-1:32'd448*32'd10];
			PixelsStore[1] <= Pixels[(32'd449+32'd1)*32'd10-1:32'd449*32'd10];
			PixelsStore[2] <= Pixels[(32'd450+32'd1)*32'd10-1:32'd450*32'd10];
			PixelsStore[3] <= Pixels[(32'd451+32'd1)*32'd10-1:32'd451*32'd10];
			PixelsStore[4] <= Pixels[(32'd452+32'd1)*32'd10-1:32'd452*32'd10];
			PixelsStore[5] <= Pixels[(32'd453+32'd1)*32'd10-1:32'd453*32'd10];
			PixelsStore[6] <= Pixels[(32'd454+32'd1)*32'd10-1:32'd454*32'd10];
			PixelsStore[7] <= Pixels[(32'd455+32'd1)*32'd10-1:32'd455*32'd10];
			PixelsStore[8] <= Pixels[(32'd456+32'd1)*32'd10-1:32'd456*32'd10];
			PixelsStore[9] <= Pixels[(32'd457+32'd1)*32'd10-1:32'd457*32'd10];
			PixelsStore[10] <= Pixels[(32'd458+32'd1)*32'd10-1:32'd458*32'd10];
			PixelsStore[11] <= Pixels[(32'd459+32'd1)*32'd10-1:32'd459*32'd10];
			PixelsStore[12] <= Pixels[(32'd460+32'd1)*32'd10-1:32'd460*32'd10];
			PixelsStore[13] <= Pixels[(32'd461+32'd1)*32'd10-1:32'd461*32'd10];
			PixelsStore[14] <= Pixels[(32'd462+32'd1)*32'd10-1:32'd462*32'd10];
			PixelsStore[15] <= Pixels[(32'd463+32'd1)*32'd10-1:32'd463*32'd10];
			PixelsStore[16] <= Pixels[(32'd464+32'd1)*32'd10-1:32'd464*32'd10];
			PixelsStore[17] <= Pixels[(32'd465+32'd1)*32'd10-1:32'd465*32'd10];
			PixelsStore[18] <= Pixels[(32'd466+32'd1)*32'd10-1:32'd466*32'd10];
			PixelsStore[19] <= Pixels[(32'd467+32'd1)*32'd10-1:32'd467*32'd10];
			PixelsStore[20] <= Pixels[(32'd468+32'd1)*32'd10-1:32'd468*32'd10];
			PixelsStore[21] <= Pixels[(32'd469+32'd1)*32'd10-1:32'd469*32'd10];
			PixelsStore[22] <= Pixels[(32'd470+32'd1)*32'd10-1:32'd470*32'd10];
			PixelsStore[23] <= Pixels[(32'd471+32'd1)*32'd10-1:32'd471*32'd10];
			PixelsStore[24] <= Pixels[(32'd472+32'd1)*32'd10-1:32'd472*32'd10];
			PixelsStore[25] <= Pixels[(32'd473+32'd1)*32'd10-1:32'd473*32'd10];
			PixelsStore[26] <= Pixels[(32'd474+32'd1)*32'd10-1:32'd474*32'd10];
			PixelsStore[27] <= Pixels[(32'd475+32'd1)*32'd10-1:32'd475*32'd10];
			WeightsStore0[0] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[1] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[2] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[3] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[4] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[5] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[6] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[7] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[8] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[9] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[10] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[11] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[12] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[13] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[14] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[15] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[16] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[17] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[18] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[19] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[20] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[21] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[22] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[23] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[24] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[25] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[26] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore0[27] <= Weights0[(32'd448+32'd1)*32'd19-1:32'd448*32'd19];
			WeightsStore1[0] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[1] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[2] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[3] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[4] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[5] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[6] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[7] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[8] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[9] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[10] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[11] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[12] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[13] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[14] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[15] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[16] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[17] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[18] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[19] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[20] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[21] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[22] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[23] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[24] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[25] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[26] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore1[27] <= Weights1[(32'd449+32'd1)*32'd19-1:32'd449*32'd19];
			WeightsStore2[0] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[1] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[2] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[3] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[4] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[5] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[6] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[7] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[8] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[9] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[10] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[11] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[12] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[13] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[14] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[15] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[16] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[17] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[18] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[19] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[20] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[21] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[22] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[23] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[24] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[25] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[26] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore2[27] <= Weights2[(32'd450+32'd1)*32'd19-1:32'd450*32'd19];
			WeightsStore3[0] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[1] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[2] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[3] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[4] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[5] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[6] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[7] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[8] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[9] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[10] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[11] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[12] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[13] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[14] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[15] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[16] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[17] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[18] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[19] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[20] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[21] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[22] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[23] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[24] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[25] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[26] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore3[27] <= Weights3[(32'd451+32'd1)*32'd19-1:32'd451*32'd19];
			WeightsStore4[0] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[1] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[2] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[3] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[4] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[5] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[6] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[7] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[8] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[9] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[10] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[11] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[12] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[13] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[14] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[15] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[16] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[17] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[18] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[19] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[20] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[21] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[22] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[23] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[24] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[25] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[26] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore4[27] <= Weights4[(32'd452+32'd1)*32'd19-1:32'd452*32'd19];
			WeightsStore5[0] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[1] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[2] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[3] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[4] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[5] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[6] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[7] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[8] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[9] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[10] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[11] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[12] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[13] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[14] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[15] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[16] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[17] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[18] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[19] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[20] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[21] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[22] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[23] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[24] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[25] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[26] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore5[27] <= Weights5[(32'd453+32'd1)*32'd19-1:32'd453*32'd19];
			WeightsStore6[0] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[1] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[2] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[3] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[4] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[5] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[6] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[7] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[8] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[9] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[10] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[11] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[12] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[13] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[14] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[15] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[16] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[17] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[18] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[19] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[20] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[21] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[22] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[23] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[24] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[25] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[26] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore6[27] <= Weights6[(32'd454+32'd1)*32'd19-1:32'd454*32'd19];
			WeightsStore7[0] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[1] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[2] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[3] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[4] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[5] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[6] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[7] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[8] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[9] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[10] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[11] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[12] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[13] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[14] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[15] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[16] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[17] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[18] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[19] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[20] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[21] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[22] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[23] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[24] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[25] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[26] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore7[27] <= Weights7[(32'd455+32'd1)*32'd19-1:32'd455*32'd19];
			WeightsStore8[0] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[1] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[2] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[3] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[4] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[5] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[6] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[7] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[8] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[9] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[10] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[11] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[12] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[13] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[14] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[15] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[16] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[17] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[18] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[19] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[20] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[21] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[22] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[23] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[24] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[25] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[26] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore8[27] <= Weights8[(32'd456+32'd1)*32'd19-1:32'd456*32'd19];
			WeightsStore9[0] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[1] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[2] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[3] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[4] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[5] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[6] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[7] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[8] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[9] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[10] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[11] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[12] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[13] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[14] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[15] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[16] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[17] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[18] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[19] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[20] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[21] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[22] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[23] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[24] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[25] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[26] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
			WeightsStore9[27] <= Weights9[(32'd457+32'd1)*32'd19-1:32'd457*32'd19];
		end else if(switchCounter == 32'd17)begin
			PixelsStore[0] <= Pixels[(32'd476+32'd1)*32'd10-1:32'd476*32'd10];
			PixelsStore[1] <= Pixels[(32'd477+32'd1)*32'd10-1:32'd477*32'd10];
			PixelsStore[2] <= Pixels[(32'd478+32'd1)*32'd10-1:32'd478*32'd10];
			PixelsStore[3] <= Pixels[(32'd479+32'd1)*32'd10-1:32'd479*32'd10];
			PixelsStore[4] <= Pixels[(32'd480+32'd1)*32'd10-1:32'd480*32'd10];
			PixelsStore[5] <= Pixels[(32'd481+32'd1)*32'd10-1:32'd481*32'd10];
			PixelsStore[6] <= Pixels[(32'd482+32'd1)*32'd10-1:32'd482*32'd10];
			PixelsStore[7] <= Pixels[(32'd483+32'd1)*32'd10-1:32'd483*32'd10];
			PixelsStore[8] <= Pixels[(32'd484+32'd1)*32'd10-1:32'd484*32'd10];
			PixelsStore[9] <= Pixels[(32'd485+32'd1)*32'd10-1:32'd485*32'd10];
			PixelsStore[10] <= Pixels[(32'd486+32'd1)*32'd10-1:32'd486*32'd10];
			PixelsStore[11] <= Pixels[(32'd487+32'd1)*32'd10-1:32'd487*32'd10];
			PixelsStore[12] <= Pixels[(32'd488+32'd1)*32'd10-1:32'd488*32'd10];
			PixelsStore[13] <= Pixels[(32'd489+32'd1)*32'd10-1:32'd489*32'd10];
			PixelsStore[14] <= Pixels[(32'd490+32'd1)*32'd10-1:32'd490*32'd10];
			PixelsStore[15] <= Pixels[(32'd491+32'd1)*32'd10-1:32'd491*32'd10];
			PixelsStore[16] <= Pixels[(32'd492+32'd1)*32'd10-1:32'd492*32'd10];
			PixelsStore[17] <= Pixels[(32'd493+32'd1)*32'd10-1:32'd493*32'd10];
			PixelsStore[18] <= Pixels[(32'd494+32'd1)*32'd10-1:32'd494*32'd10];
			PixelsStore[19] <= Pixels[(32'd495+32'd1)*32'd10-1:32'd495*32'd10];
			PixelsStore[20] <= Pixels[(32'd496+32'd1)*32'd10-1:32'd496*32'd10];
			PixelsStore[21] <= Pixels[(32'd497+32'd1)*32'd10-1:32'd497*32'd10];
			PixelsStore[22] <= Pixels[(32'd498+32'd1)*32'd10-1:32'd498*32'd10];
			PixelsStore[23] <= Pixels[(32'd499+32'd1)*32'd10-1:32'd499*32'd10];
			PixelsStore[24] <= Pixels[(32'd500+32'd1)*32'd10-1:32'd500*32'd10];
			PixelsStore[25] <= Pixels[(32'd501+32'd1)*32'd10-1:32'd501*32'd10];
			PixelsStore[26] <= Pixels[(32'd502+32'd1)*32'd10-1:32'd502*32'd10];
			PixelsStore[27] <= Pixels[(32'd503+32'd1)*32'd10-1:32'd503*32'd10];
			WeightsStore0[0] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[1] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[2] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[3] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[4] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[5] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[6] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[7] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[8] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[9] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[10] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[11] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[12] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[13] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[14] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[15] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[16] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[17] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[18] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[19] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[20] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[21] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[22] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[23] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[24] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[25] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[26] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore0[27] <= Weights0[(32'd476+32'd1)*32'd19-1:32'd476*32'd19];
			WeightsStore1[0] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[1] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[2] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[3] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[4] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[5] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[6] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[7] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[8] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[9] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[10] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[11] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[12] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[13] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[14] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[15] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[16] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[17] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[18] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[19] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[20] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[21] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[22] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[23] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[24] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[25] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[26] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore1[27] <= Weights1[(32'd477+32'd1)*32'd19-1:32'd477*32'd19];
			WeightsStore2[0] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[1] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[2] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[3] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[4] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[5] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[6] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[7] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[8] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[9] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[10] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[11] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[12] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[13] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[14] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[15] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[16] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[17] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[18] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[19] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[20] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[21] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[22] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[23] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[24] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[25] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[26] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore2[27] <= Weights2[(32'd478+32'd1)*32'd19-1:32'd478*32'd19];
			WeightsStore3[0] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[1] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[2] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[3] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[4] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[5] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[6] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[7] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[8] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[9] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[10] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[11] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[12] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[13] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[14] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[15] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[16] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[17] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[18] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[19] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[20] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[21] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[22] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[23] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[24] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[25] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[26] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore3[27] <= Weights3[(32'd479+32'd1)*32'd19-1:32'd479*32'd19];
			WeightsStore4[0] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[1] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[2] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[3] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[4] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[5] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[6] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[7] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[8] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[9] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[10] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[11] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[12] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[13] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[14] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[15] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[16] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[17] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[18] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[19] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[20] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[21] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[22] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[23] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[24] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[25] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[26] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore4[27] <= Weights4[(32'd480+32'd1)*32'd19-1:32'd480*32'd19];
			WeightsStore5[0] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[1] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[2] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[3] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[4] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[5] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[6] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[7] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[8] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[9] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[10] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[11] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[12] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[13] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[14] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[15] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[16] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[17] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[18] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[19] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[20] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[21] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[22] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[23] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[24] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[25] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[26] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore5[27] <= Weights5[(32'd481+32'd1)*32'd19-1:32'd481*32'd19];
			WeightsStore6[0] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[1] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[2] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[3] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[4] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[5] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[6] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[7] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[8] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[9] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[10] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[11] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[12] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[13] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[14] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[15] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[16] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[17] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[18] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[19] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[20] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[21] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[22] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[23] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[24] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[25] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[26] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore6[27] <= Weights6[(32'd482+32'd1)*32'd19-1:32'd482*32'd19];
			WeightsStore7[0] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[1] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[2] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[3] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[4] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[5] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[6] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[7] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[8] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[9] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[10] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[11] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[12] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[13] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[14] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[15] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[16] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[17] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[18] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[19] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[20] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[21] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[22] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[23] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[24] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[25] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[26] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore7[27] <= Weights7[(32'd483+32'd1)*32'd19-1:32'd483*32'd19];
			WeightsStore8[0] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[1] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[2] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[3] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[4] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[5] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[6] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[7] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[8] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[9] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[10] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[11] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[12] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[13] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[14] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[15] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[16] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[17] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[18] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[19] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[20] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[21] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[22] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[23] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[24] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[25] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[26] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore8[27] <= Weights8[(32'd484+32'd1)*32'd19-1:32'd484*32'd19];
			WeightsStore9[0] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[1] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[2] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[3] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[4] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[5] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[6] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[7] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[8] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[9] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[10] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[11] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[12] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[13] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[14] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[15] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[16] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[17] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[18] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[19] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[20] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[21] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[22] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[23] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[24] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[25] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[26] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
			WeightsStore9[27] <= Weights9[(32'd485+32'd1)*32'd19-1:32'd485*32'd19];
		end else if(switchCounter == 32'd18)begin
			PixelsStore[0] <= Pixels[(32'd504+32'd1)*32'd10-1:32'd504*32'd10];
			PixelsStore[1] <= Pixels[(32'd505+32'd1)*32'd10-1:32'd505*32'd10];
			PixelsStore[2] <= Pixels[(32'd506+32'd1)*32'd10-1:32'd506*32'd10];
			PixelsStore[3] <= Pixels[(32'd507+32'd1)*32'd10-1:32'd507*32'd10];
			PixelsStore[4] <= Pixels[(32'd508+32'd1)*32'd10-1:32'd508*32'd10];
			PixelsStore[5] <= Pixels[(32'd509+32'd1)*32'd10-1:32'd509*32'd10];
			PixelsStore[6] <= Pixels[(32'd510+32'd1)*32'd10-1:32'd510*32'd10];
			PixelsStore[7] <= Pixels[(32'd511+32'd1)*32'd10-1:32'd511*32'd10];
			PixelsStore[8] <= Pixels[(32'd512+32'd1)*32'd10-1:32'd512*32'd10];
			PixelsStore[9] <= Pixels[(32'd513+32'd1)*32'd10-1:32'd513*32'd10];
			PixelsStore[10] <= Pixels[(32'd514+32'd1)*32'd10-1:32'd514*32'd10];
			PixelsStore[11] <= Pixels[(32'd515+32'd1)*32'd10-1:32'd515*32'd10];
			PixelsStore[12] <= Pixels[(32'd516+32'd1)*32'd10-1:32'd516*32'd10];
			PixelsStore[13] <= Pixels[(32'd517+32'd1)*32'd10-1:32'd517*32'd10];
			PixelsStore[14] <= Pixels[(32'd518+32'd1)*32'd10-1:32'd518*32'd10];
			PixelsStore[15] <= Pixels[(32'd519+32'd1)*32'd10-1:32'd519*32'd10];
			PixelsStore[16] <= Pixels[(32'd520+32'd1)*32'd10-1:32'd520*32'd10];
			PixelsStore[17] <= Pixels[(32'd521+32'd1)*32'd10-1:32'd521*32'd10];
			PixelsStore[18] <= Pixels[(32'd522+32'd1)*32'd10-1:32'd522*32'd10];
			PixelsStore[19] <= Pixels[(32'd523+32'd1)*32'd10-1:32'd523*32'd10];
			PixelsStore[20] <= Pixels[(32'd524+32'd1)*32'd10-1:32'd524*32'd10];
			PixelsStore[21] <= Pixels[(32'd525+32'd1)*32'd10-1:32'd525*32'd10];
			PixelsStore[22] <= Pixels[(32'd526+32'd1)*32'd10-1:32'd526*32'd10];
			PixelsStore[23] <= Pixels[(32'd527+32'd1)*32'd10-1:32'd527*32'd10];
			PixelsStore[24] <= Pixels[(32'd528+32'd1)*32'd10-1:32'd528*32'd10];
			PixelsStore[25] <= Pixels[(32'd529+32'd1)*32'd10-1:32'd529*32'd10];
			PixelsStore[26] <= Pixels[(32'd530+32'd1)*32'd10-1:32'd530*32'd10];
			PixelsStore[27] <= Pixels[(32'd531+32'd1)*32'd10-1:32'd531*32'd10];
			WeightsStore0[0] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[1] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[2] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[3] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[4] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[5] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[6] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[7] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[8] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[9] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[10] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[11] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[12] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[13] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[14] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[15] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[16] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[17] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[18] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[19] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[20] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[21] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[22] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[23] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[24] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[25] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[26] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore0[27] <= Weights0[(32'd504+32'd1)*32'd19-1:32'd504*32'd19];
			WeightsStore1[0] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[1] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[2] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[3] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[4] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[5] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[6] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[7] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[8] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[9] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[10] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[11] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[12] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[13] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[14] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[15] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[16] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[17] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[18] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[19] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[20] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[21] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[22] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[23] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[24] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[25] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[26] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore1[27] <= Weights1[(32'd505+32'd1)*32'd19-1:32'd505*32'd19];
			WeightsStore2[0] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[1] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[2] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[3] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[4] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[5] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[6] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[7] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[8] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[9] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[10] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[11] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[12] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[13] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[14] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[15] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[16] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[17] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[18] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[19] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[20] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[21] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[22] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[23] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[24] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[25] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[26] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore2[27] <= Weights2[(32'd506+32'd1)*32'd19-1:32'd506*32'd19];
			WeightsStore3[0] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[1] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[2] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[3] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[4] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[5] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[6] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[7] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[8] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[9] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[10] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[11] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[12] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[13] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[14] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[15] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[16] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[17] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[18] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[19] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[20] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[21] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[22] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[23] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[24] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[25] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[26] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore3[27] <= Weights3[(32'd507+32'd1)*32'd19-1:32'd507*32'd19];
			WeightsStore4[0] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[1] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[2] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[3] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[4] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[5] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[6] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[7] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[8] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[9] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[10] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[11] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[12] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[13] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[14] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[15] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[16] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[17] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[18] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[19] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[20] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[21] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[22] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[23] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[24] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[25] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[26] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore4[27] <= Weights4[(32'd508+32'd1)*32'd19-1:32'd508*32'd19];
			WeightsStore5[0] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[1] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[2] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[3] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[4] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[5] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[6] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[7] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[8] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[9] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[10] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[11] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[12] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[13] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[14] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[15] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[16] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[17] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[18] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[19] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[20] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[21] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[22] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[23] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[24] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[25] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[26] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore5[27] <= Weights5[(32'd509+32'd1)*32'd19-1:32'd509*32'd19];
			WeightsStore6[0] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[1] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[2] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[3] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[4] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[5] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[6] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[7] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[8] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[9] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[10] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[11] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[12] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[13] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[14] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[15] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[16] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[17] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[18] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[19] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[20] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[21] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[22] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[23] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[24] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[25] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[26] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore6[27] <= Weights6[(32'd510+32'd1)*32'd19-1:32'd510*32'd19];
			WeightsStore7[0] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[1] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[2] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[3] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[4] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[5] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[6] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[7] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[8] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[9] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[10] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[11] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[12] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[13] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[14] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[15] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[16] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[17] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[18] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[19] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[20] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[21] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[22] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[23] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[24] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[25] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[26] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore7[27] <= Weights7[(32'd511+32'd1)*32'd19-1:32'd511*32'd19];
			WeightsStore8[0] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[1] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[2] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[3] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[4] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[5] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[6] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[7] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[8] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[9] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[10] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[11] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[12] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[13] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[14] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[15] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[16] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[17] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[18] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[19] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[20] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[21] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[22] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[23] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[24] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[25] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[26] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore8[27] <= Weights8[(32'd512+32'd1)*32'd19-1:32'd512*32'd19];
			WeightsStore9[0] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[1] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[2] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[3] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[4] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[5] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[6] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[7] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[8] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[9] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[10] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[11] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[12] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[13] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[14] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[15] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[16] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[17] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[18] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[19] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[20] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[21] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[22] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[23] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[24] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[25] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[26] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
			WeightsStore9[27] <= Weights9[(32'd513+32'd1)*32'd19-1:32'd513*32'd19];
		end else if(switchCounter == 32'd19)begin
			PixelsStore[0] <= Pixels[(32'd532+32'd1)*32'd10-1:32'd532*32'd10];
			PixelsStore[1] <= Pixels[(32'd533+32'd1)*32'd10-1:32'd533*32'd10];
			PixelsStore[2] <= Pixels[(32'd534+32'd1)*32'd10-1:32'd534*32'd10];
			PixelsStore[3] <= Pixels[(32'd535+32'd1)*32'd10-1:32'd535*32'd10];
			PixelsStore[4] <= Pixels[(32'd536+32'd1)*32'd10-1:32'd536*32'd10];
			PixelsStore[5] <= Pixels[(32'd537+32'd1)*32'd10-1:32'd537*32'd10];
			PixelsStore[6] <= Pixels[(32'd538+32'd1)*32'd10-1:32'd538*32'd10];
			PixelsStore[7] <= Pixels[(32'd539+32'd1)*32'd10-1:32'd539*32'd10];
			PixelsStore[8] <= Pixels[(32'd540+32'd1)*32'd10-1:32'd540*32'd10];
			PixelsStore[9] <= Pixels[(32'd541+32'd1)*32'd10-1:32'd541*32'd10];
			PixelsStore[10] <= Pixels[(32'd542+32'd1)*32'd10-1:32'd542*32'd10];
			PixelsStore[11] <= Pixels[(32'd543+32'd1)*32'd10-1:32'd543*32'd10];
			PixelsStore[12] <= Pixels[(32'd544+32'd1)*32'd10-1:32'd544*32'd10];
			PixelsStore[13] <= Pixels[(32'd545+32'd1)*32'd10-1:32'd545*32'd10];
			PixelsStore[14] <= Pixels[(32'd546+32'd1)*32'd10-1:32'd546*32'd10];
			PixelsStore[15] <= Pixels[(32'd547+32'd1)*32'd10-1:32'd547*32'd10];
			PixelsStore[16] <= Pixels[(32'd548+32'd1)*32'd10-1:32'd548*32'd10];
			PixelsStore[17] <= Pixels[(32'd549+32'd1)*32'd10-1:32'd549*32'd10];
			PixelsStore[18] <= Pixels[(32'd550+32'd1)*32'd10-1:32'd550*32'd10];
			PixelsStore[19] <= Pixels[(32'd551+32'd1)*32'd10-1:32'd551*32'd10];
			PixelsStore[20] <= Pixels[(32'd552+32'd1)*32'd10-1:32'd552*32'd10];
			PixelsStore[21] <= Pixels[(32'd553+32'd1)*32'd10-1:32'd553*32'd10];
			PixelsStore[22] <= Pixels[(32'd554+32'd1)*32'd10-1:32'd554*32'd10];
			PixelsStore[23] <= Pixels[(32'd555+32'd1)*32'd10-1:32'd555*32'd10];
			PixelsStore[24] <= Pixels[(32'd556+32'd1)*32'd10-1:32'd556*32'd10];
			PixelsStore[25] <= Pixels[(32'd557+32'd1)*32'd10-1:32'd557*32'd10];
			PixelsStore[26] <= Pixels[(32'd558+32'd1)*32'd10-1:32'd558*32'd10];
			PixelsStore[27] <= Pixels[(32'd559+32'd1)*32'd10-1:32'd559*32'd10];
			WeightsStore0[0] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[1] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[2] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[3] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[4] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[5] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[6] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[7] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[8] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[9] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[10] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[11] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[12] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[13] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[14] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[15] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[16] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[17] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[18] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[19] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[20] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[21] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[22] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[23] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[24] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[25] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[26] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore0[27] <= Weights0[(32'd532+32'd1)*32'd19-1:32'd532*32'd19];
			WeightsStore1[0] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[1] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[2] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[3] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[4] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[5] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[6] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[7] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[8] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[9] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[10] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[11] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[12] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[13] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[14] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[15] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[16] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[17] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[18] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[19] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[20] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[21] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[22] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[23] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[24] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[25] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[26] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore1[27] <= Weights1[(32'd533+32'd1)*32'd19-1:32'd533*32'd19];
			WeightsStore2[0] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[1] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[2] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[3] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[4] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[5] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[6] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[7] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[8] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[9] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[10] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[11] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[12] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[13] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[14] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[15] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[16] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[17] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[18] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[19] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[20] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[21] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[22] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[23] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[24] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[25] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[26] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore2[27] <= Weights2[(32'd534+32'd1)*32'd19-1:32'd534*32'd19];
			WeightsStore3[0] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[1] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[2] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[3] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[4] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[5] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[6] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[7] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[8] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[9] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[10] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[11] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[12] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[13] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[14] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[15] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[16] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[17] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[18] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[19] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[20] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[21] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[22] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[23] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[24] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[25] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[26] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore3[27] <= Weights3[(32'd535+32'd1)*32'd19-1:32'd535*32'd19];
			WeightsStore4[0] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[1] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[2] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[3] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[4] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[5] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[6] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[7] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[8] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[9] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[10] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[11] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[12] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[13] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[14] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[15] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[16] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[17] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[18] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[19] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[20] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[21] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[22] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[23] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[24] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[25] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[26] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore4[27] <= Weights4[(32'd536+32'd1)*32'd19-1:32'd536*32'd19];
			WeightsStore5[0] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[1] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[2] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[3] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[4] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[5] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[6] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[7] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[8] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[9] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[10] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[11] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[12] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[13] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[14] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[15] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[16] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[17] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[18] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[19] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[20] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[21] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[22] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[23] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[24] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[25] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[26] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore5[27] <= Weights5[(32'd537+32'd1)*32'd19-1:32'd537*32'd19];
			WeightsStore6[0] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[1] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[2] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[3] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[4] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[5] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[6] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[7] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[8] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[9] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[10] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[11] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[12] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[13] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[14] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[15] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[16] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[17] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[18] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[19] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[20] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[21] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[22] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[23] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[24] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[25] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[26] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore6[27] <= Weights6[(32'd538+32'd1)*32'd19-1:32'd538*32'd19];
			WeightsStore7[0] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[1] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[2] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[3] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[4] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[5] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[6] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[7] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[8] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[9] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[10] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[11] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[12] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[13] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[14] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[15] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[16] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[17] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[18] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[19] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[20] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[21] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[22] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[23] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[24] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[25] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[26] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore7[27] <= Weights7[(32'd539+32'd1)*32'd19-1:32'd539*32'd19];
			WeightsStore8[0] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[1] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[2] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[3] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[4] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[5] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[6] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[7] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[8] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[9] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[10] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[11] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[12] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[13] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[14] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[15] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[16] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[17] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[18] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[19] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[20] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[21] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[22] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[23] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[24] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[25] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[26] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore8[27] <= Weights8[(32'd540+32'd1)*32'd19-1:32'd540*32'd19];
			WeightsStore9[0] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[1] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[2] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[3] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[4] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[5] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[6] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[7] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[8] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[9] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[10] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[11] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[12] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[13] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[14] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[15] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[16] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[17] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[18] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[19] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[20] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[21] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[22] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[23] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[24] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[25] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[26] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
			WeightsStore9[27] <= Weights9[(32'd541+32'd1)*32'd19-1:32'd541*32'd19];
		end else if(switchCounter == 32'd20)begin
			PixelsStore[0] <= Pixels[(32'd560+32'd1)*32'd10-1:32'd560*32'd10];
			PixelsStore[1] <= Pixels[(32'd561+32'd1)*32'd10-1:32'd561*32'd10];
			PixelsStore[2] <= Pixels[(32'd562+32'd1)*32'd10-1:32'd562*32'd10];
			PixelsStore[3] <= Pixels[(32'd563+32'd1)*32'd10-1:32'd563*32'd10];
			PixelsStore[4] <= Pixels[(32'd564+32'd1)*32'd10-1:32'd564*32'd10];
			PixelsStore[5] <= Pixels[(32'd565+32'd1)*32'd10-1:32'd565*32'd10];
			PixelsStore[6] <= Pixels[(32'd566+32'd1)*32'd10-1:32'd566*32'd10];
			PixelsStore[7] <= Pixels[(32'd567+32'd1)*32'd10-1:32'd567*32'd10];
			PixelsStore[8] <= Pixels[(32'd568+32'd1)*32'd10-1:32'd568*32'd10];
			PixelsStore[9] <= Pixels[(32'd569+32'd1)*32'd10-1:32'd569*32'd10];
			PixelsStore[10] <= Pixels[(32'd570+32'd1)*32'd10-1:32'd570*32'd10];
			PixelsStore[11] <= Pixels[(32'd571+32'd1)*32'd10-1:32'd571*32'd10];
			PixelsStore[12] <= Pixels[(32'd572+32'd1)*32'd10-1:32'd572*32'd10];
			PixelsStore[13] <= Pixels[(32'd573+32'd1)*32'd10-1:32'd573*32'd10];
			PixelsStore[14] <= Pixels[(32'd574+32'd1)*32'd10-1:32'd574*32'd10];
			PixelsStore[15] <= Pixels[(32'd575+32'd1)*32'd10-1:32'd575*32'd10];
			PixelsStore[16] <= Pixels[(32'd576+32'd1)*32'd10-1:32'd576*32'd10];
			PixelsStore[17] <= Pixels[(32'd577+32'd1)*32'd10-1:32'd577*32'd10];
			PixelsStore[18] <= Pixels[(32'd578+32'd1)*32'd10-1:32'd578*32'd10];
			PixelsStore[19] <= Pixels[(32'd579+32'd1)*32'd10-1:32'd579*32'd10];
			PixelsStore[20] <= Pixels[(32'd580+32'd1)*32'd10-1:32'd580*32'd10];
			PixelsStore[21] <= Pixels[(32'd581+32'd1)*32'd10-1:32'd581*32'd10];
			PixelsStore[22] <= Pixels[(32'd582+32'd1)*32'd10-1:32'd582*32'd10];
			PixelsStore[23] <= Pixels[(32'd583+32'd1)*32'd10-1:32'd583*32'd10];
			PixelsStore[24] <= Pixels[(32'd584+32'd1)*32'd10-1:32'd584*32'd10];
			PixelsStore[25] <= Pixels[(32'd585+32'd1)*32'd10-1:32'd585*32'd10];
			PixelsStore[26] <= Pixels[(32'd586+32'd1)*32'd10-1:32'd586*32'd10];
			PixelsStore[27] <= Pixels[(32'd587+32'd1)*32'd10-1:32'd587*32'd10];
			WeightsStore0[0] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[1] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[2] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[3] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[4] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[5] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[6] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[7] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[8] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[9] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[10] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[11] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[12] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[13] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[14] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[15] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[16] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[17] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[18] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[19] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[20] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[21] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[22] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[23] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[24] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[25] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[26] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore0[27] <= Weights0[(32'd560+32'd1)*32'd19-1:32'd560*32'd19];
			WeightsStore1[0] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[1] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[2] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[3] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[4] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[5] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[6] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[7] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[8] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[9] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[10] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[11] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[12] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[13] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[14] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[15] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[16] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[17] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[18] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[19] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[20] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[21] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[22] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[23] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[24] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[25] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[26] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore1[27] <= Weights1[(32'd561+32'd1)*32'd19-1:32'd561*32'd19];
			WeightsStore2[0] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[1] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[2] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[3] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[4] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[5] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[6] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[7] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[8] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[9] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[10] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[11] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[12] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[13] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[14] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[15] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[16] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[17] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[18] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[19] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[20] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[21] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[22] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[23] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[24] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[25] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[26] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore2[27] <= Weights2[(32'd562+32'd1)*32'd19-1:32'd562*32'd19];
			WeightsStore3[0] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[1] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[2] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[3] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[4] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[5] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[6] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[7] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[8] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[9] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[10] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[11] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[12] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[13] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[14] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[15] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[16] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[17] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[18] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[19] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[20] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[21] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[22] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[23] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[24] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[25] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[26] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore3[27] <= Weights3[(32'd563+32'd1)*32'd19-1:32'd563*32'd19];
			WeightsStore4[0] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[1] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[2] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[3] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[4] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[5] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[6] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[7] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[8] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[9] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[10] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[11] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[12] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[13] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[14] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[15] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[16] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[17] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[18] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[19] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[20] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[21] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[22] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[23] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[24] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[25] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[26] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore4[27] <= Weights4[(32'd564+32'd1)*32'd19-1:32'd564*32'd19];
			WeightsStore5[0] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[1] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[2] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[3] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[4] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[5] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[6] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[7] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[8] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[9] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[10] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[11] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[12] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[13] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[14] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[15] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[16] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[17] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[18] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[19] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[20] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[21] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[22] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[23] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[24] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[25] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[26] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore5[27] <= Weights5[(32'd565+32'd1)*32'd19-1:32'd565*32'd19];
			WeightsStore6[0] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[1] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[2] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[3] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[4] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[5] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[6] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[7] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[8] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[9] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[10] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[11] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[12] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[13] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[14] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[15] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[16] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[17] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[18] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[19] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[20] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[21] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[22] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[23] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[24] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[25] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[26] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore6[27] <= Weights6[(32'd566+32'd1)*32'd19-1:32'd566*32'd19];
			WeightsStore7[0] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[1] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[2] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[3] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[4] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[5] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[6] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[7] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[8] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[9] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[10] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[11] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[12] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[13] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[14] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[15] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[16] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[17] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[18] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[19] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[20] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[21] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[22] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[23] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[24] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[25] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[26] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore7[27] <= Weights7[(32'd567+32'd1)*32'd19-1:32'd567*32'd19];
			WeightsStore8[0] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[1] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[2] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[3] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[4] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[5] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[6] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[7] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[8] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[9] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[10] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[11] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[12] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[13] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[14] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[15] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[16] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[17] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[18] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[19] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[20] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[21] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[22] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[23] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[24] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[25] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[26] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore8[27] <= Weights8[(32'd568+32'd1)*32'd19-1:32'd568*32'd19];
			WeightsStore9[0] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[1] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[2] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[3] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[4] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[5] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[6] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[7] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[8] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[9] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[10] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[11] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[12] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[13] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[14] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[15] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[16] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[17] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[18] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[19] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[20] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[21] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[22] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[23] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[24] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[25] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[26] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
			WeightsStore9[27] <= Weights9[(32'd569+32'd1)*32'd19-1:32'd569*32'd19];
		end else if(switchCounter == 32'd21)begin
			PixelsStore[0] <= Pixels[(32'd588+32'd1)*32'd10-1:32'd588*32'd10];
			PixelsStore[1] <= Pixels[(32'd589+32'd1)*32'd10-1:32'd589*32'd10];
			PixelsStore[2] <= Pixels[(32'd590+32'd1)*32'd10-1:32'd590*32'd10];
			PixelsStore[3] <= Pixels[(32'd591+32'd1)*32'd10-1:32'd591*32'd10];
			PixelsStore[4] <= Pixels[(32'd592+32'd1)*32'd10-1:32'd592*32'd10];
			PixelsStore[5] <= Pixels[(32'd593+32'd1)*32'd10-1:32'd593*32'd10];
			PixelsStore[6] <= Pixels[(32'd594+32'd1)*32'd10-1:32'd594*32'd10];
			PixelsStore[7] <= Pixels[(32'd595+32'd1)*32'd10-1:32'd595*32'd10];
			PixelsStore[8] <= Pixels[(32'd596+32'd1)*32'd10-1:32'd596*32'd10];
			PixelsStore[9] <= Pixels[(32'd597+32'd1)*32'd10-1:32'd597*32'd10];
			PixelsStore[10] <= Pixels[(32'd598+32'd1)*32'd10-1:32'd598*32'd10];
			PixelsStore[11] <= Pixels[(32'd599+32'd1)*32'd10-1:32'd599*32'd10];
			PixelsStore[12] <= Pixels[(32'd600+32'd1)*32'd10-1:32'd600*32'd10];
			PixelsStore[13] <= Pixels[(32'd601+32'd1)*32'd10-1:32'd601*32'd10];
			PixelsStore[14] <= Pixels[(32'd602+32'd1)*32'd10-1:32'd602*32'd10];
			PixelsStore[15] <= Pixels[(32'd603+32'd1)*32'd10-1:32'd603*32'd10];
			PixelsStore[16] <= Pixels[(32'd604+32'd1)*32'd10-1:32'd604*32'd10];
			PixelsStore[17] <= Pixels[(32'd605+32'd1)*32'd10-1:32'd605*32'd10];
			PixelsStore[18] <= Pixels[(32'd606+32'd1)*32'd10-1:32'd606*32'd10];
			PixelsStore[19] <= Pixels[(32'd607+32'd1)*32'd10-1:32'd607*32'd10];
			PixelsStore[20] <= Pixels[(32'd608+32'd1)*32'd10-1:32'd608*32'd10];
			PixelsStore[21] <= Pixels[(32'd609+32'd1)*32'd10-1:32'd609*32'd10];
			PixelsStore[22] <= Pixels[(32'd610+32'd1)*32'd10-1:32'd610*32'd10];
			PixelsStore[23] <= Pixels[(32'd611+32'd1)*32'd10-1:32'd611*32'd10];
			PixelsStore[24] <= Pixels[(32'd612+32'd1)*32'd10-1:32'd612*32'd10];
			PixelsStore[25] <= Pixels[(32'd613+32'd1)*32'd10-1:32'd613*32'd10];
			PixelsStore[26] <= Pixels[(32'd614+32'd1)*32'd10-1:32'd614*32'd10];
			PixelsStore[27] <= Pixels[(32'd615+32'd1)*32'd10-1:32'd615*32'd10];
			WeightsStore0[0] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[1] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[2] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[3] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[4] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[5] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[6] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[7] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[8] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[9] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[10] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[11] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[12] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[13] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[14] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[15] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[16] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[17] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[18] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[19] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[20] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[21] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[22] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[23] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[24] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[25] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[26] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore0[27] <= Weights0[(32'd588+32'd1)*32'd19-1:32'd588*32'd19];
			WeightsStore1[0] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[1] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[2] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[3] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[4] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[5] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[6] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[7] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[8] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[9] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[10] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[11] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[12] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[13] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[14] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[15] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[16] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[17] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[18] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[19] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[20] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[21] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[22] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[23] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[24] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[25] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[26] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore1[27] <= Weights1[(32'd589+32'd1)*32'd19-1:32'd589*32'd19];
			WeightsStore2[0] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[1] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[2] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[3] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[4] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[5] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[6] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[7] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[8] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[9] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[10] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[11] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[12] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[13] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[14] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[15] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[16] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[17] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[18] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[19] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[20] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[21] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[22] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[23] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[24] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[25] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[26] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore2[27] <= Weights2[(32'd590+32'd1)*32'd19-1:32'd590*32'd19];
			WeightsStore3[0] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[1] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[2] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[3] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[4] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[5] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[6] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[7] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[8] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[9] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[10] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[11] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[12] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[13] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[14] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[15] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[16] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[17] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[18] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[19] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[20] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[21] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[22] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[23] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[24] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[25] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[26] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore3[27] <= Weights3[(32'd591+32'd1)*32'd19-1:32'd591*32'd19];
			WeightsStore4[0] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[1] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[2] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[3] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[4] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[5] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[6] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[7] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[8] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[9] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[10] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[11] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[12] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[13] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[14] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[15] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[16] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[17] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[18] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[19] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[20] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[21] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[22] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[23] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[24] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[25] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[26] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore4[27] <= Weights4[(32'd592+32'd1)*32'd19-1:32'd592*32'd19];
			WeightsStore5[0] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[1] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[2] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[3] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[4] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[5] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[6] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[7] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[8] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[9] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[10] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[11] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[12] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[13] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[14] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[15] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[16] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[17] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[18] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[19] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[20] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[21] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[22] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[23] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[24] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[25] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[26] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore5[27] <= Weights5[(32'd593+32'd1)*32'd19-1:32'd593*32'd19];
			WeightsStore6[0] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[1] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[2] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[3] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[4] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[5] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[6] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[7] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[8] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[9] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[10] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[11] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[12] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[13] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[14] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[15] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[16] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[17] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[18] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[19] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[20] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[21] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[22] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[23] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[24] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[25] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[26] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore6[27] <= Weights6[(32'd594+32'd1)*32'd19-1:32'd594*32'd19];
			WeightsStore7[0] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[1] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[2] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[3] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[4] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[5] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[6] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[7] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[8] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[9] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[10] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[11] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[12] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[13] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[14] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[15] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[16] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[17] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[18] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[19] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[20] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[21] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[22] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[23] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[24] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[25] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[26] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore7[27] <= Weights7[(32'd595+32'd1)*32'd19-1:32'd595*32'd19];
			WeightsStore8[0] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[1] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[2] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[3] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[4] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[5] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[6] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[7] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[8] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[9] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[10] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[11] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[12] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[13] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[14] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[15] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[16] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[17] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[18] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[19] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[20] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[21] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[22] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[23] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[24] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[25] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[26] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore8[27] <= Weights8[(32'd596+32'd1)*32'd19-1:32'd596*32'd19];
			WeightsStore9[0] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[1] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[2] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[3] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[4] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[5] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[6] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[7] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[8] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[9] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[10] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[11] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[12] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[13] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[14] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[15] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[16] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[17] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[18] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[19] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[20] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[21] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[22] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[23] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[24] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[25] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[26] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
			WeightsStore9[27] <= Weights9[(32'd597+32'd1)*32'd19-1:32'd597*32'd19];
		end else if(switchCounter == 32'd22)begin
			PixelsStore[0] <= Pixels[(32'd616+32'd1)*32'd10-1:32'd616*32'd10];
			PixelsStore[1] <= Pixels[(32'd617+32'd1)*32'd10-1:32'd617*32'd10];
			PixelsStore[2] <= Pixels[(32'd618+32'd1)*32'd10-1:32'd618*32'd10];
			PixelsStore[3] <= Pixels[(32'd619+32'd1)*32'd10-1:32'd619*32'd10];
			PixelsStore[4] <= Pixels[(32'd620+32'd1)*32'd10-1:32'd620*32'd10];
			PixelsStore[5] <= Pixels[(32'd621+32'd1)*32'd10-1:32'd621*32'd10];
			PixelsStore[6] <= Pixels[(32'd622+32'd1)*32'd10-1:32'd622*32'd10];
			PixelsStore[7] <= Pixels[(32'd623+32'd1)*32'd10-1:32'd623*32'd10];
			PixelsStore[8] <= Pixels[(32'd624+32'd1)*32'd10-1:32'd624*32'd10];
			PixelsStore[9] <= Pixels[(32'd625+32'd1)*32'd10-1:32'd625*32'd10];
			PixelsStore[10] <= Pixels[(32'd626+32'd1)*32'd10-1:32'd626*32'd10];
			PixelsStore[11] <= Pixels[(32'd627+32'd1)*32'd10-1:32'd627*32'd10];
			PixelsStore[12] <= Pixels[(32'd628+32'd1)*32'd10-1:32'd628*32'd10];
			PixelsStore[13] <= Pixels[(32'd629+32'd1)*32'd10-1:32'd629*32'd10];
			PixelsStore[14] <= Pixels[(32'd630+32'd1)*32'd10-1:32'd630*32'd10];
			PixelsStore[15] <= Pixels[(32'd631+32'd1)*32'd10-1:32'd631*32'd10];
			PixelsStore[16] <= Pixels[(32'd632+32'd1)*32'd10-1:32'd632*32'd10];
			PixelsStore[17] <= Pixels[(32'd633+32'd1)*32'd10-1:32'd633*32'd10];
			PixelsStore[18] <= Pixels[(32'd634+32'd1)*32'd10-1:32'd634*32'd10];
			PixelsStore[19] <= Pixels[(32'd635+32'd1)*32'd10-1:32'd635*32'd10];
			PixelsStore[20] <= Pixels[(32'd636+32'd1)*32'd10-1:32'd636*32'd10];
			PixelsStore[21] <= Pixels[(32'd637+32'd1)*32'd10-1:32'd637*32'd10];
			PixelsStore[22] <= Pixels[(32'd638+32'd1)*32'd10-1:32'd638*32'd10];
			PixelsStore[23] <= Pixels[(32'd639+32'd1)*32'd10-1:32'd639*32'd10];
			PixelsStore[24] <= Pixels[(32'd640+32'd1)*32'd10-1:32'd640*32'd10];
			PixelsStore[25] <= Pixels[(32'd641+32'd1)*32'd10-1:32'd641*32'd10];
			PixelsStore[26] <= Pixels[(32'd642+32'd1)*32'd10-1:32'd642*32'd10];
			PixelsStore[27] <= Pixels[(32'd643+32'd1)*32'd10-1:32'd643*32'd10];
			WeightsStore0[0] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[1] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[2] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[3] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[4] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[5] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[6] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[7] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[8] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[9] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[10] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[11] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[12] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[13] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[14] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[15] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[16] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[17] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[18] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[19] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[20] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[21] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[22] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[23] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[24] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[25] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[26] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore0[27] <= Weights0[(32'd616+32'd1)*32'd19-1:32'd616*32'd19];
			WeightsStore1[0] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[1] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[2] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[3] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[4] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[5] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[6] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[7] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[8] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[9] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[10] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[11] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[12] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[13] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[14] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[15] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[16] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[17] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[18] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[19] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[20] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[21] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[22] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[23] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[24] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[25] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[26] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore1[27] <= Weights1[(32'd617+32'd1)*32'd19-1:32'd617*32'd19];
			WeightsStore2[0] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[1] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[2] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[3] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[4] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[5] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[6] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[7] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[8] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[9] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[10] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[11] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[12] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[13] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[14] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[15] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[16] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[17] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[18] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[19] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[20] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[21] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[22] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[23] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[24] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[25] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[26] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore2[27] <= Weights2[(32'd618+32'd1)*32'd19-1:32'd618*32'd19];
			WeightsStore3[0] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[1] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[2] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[3] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[4] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[5] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[6] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[7] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[8] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[9] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[10] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[11] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[12] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[13] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[14] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[15] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[16] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[17] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[18] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[19] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[20] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[21] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[22] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[23] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[24] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[25] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[26] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore3[27] <= Weights3[(32'd619+32'd1)*32'd19-1:32'd619*32'd19];
			WeightsStore4[0] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[1] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[2] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[3] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[4] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[5] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[6] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[7] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[8] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[9] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[10] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[11] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[12] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[13] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[14] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[15] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[16] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[17] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[18] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[19] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[20] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[21] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[22] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[23] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[24] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[25] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[26] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore4[27] <= Weights4[(32'd620+32'd1)*32'd19-1:32'd620*32'd19];
			WeightsStore5[0] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[1] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[2] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[3] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[4] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[5] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[6] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[7] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[8] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[9] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[10] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[11] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[12] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[13] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[14] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[15] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[16] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[17] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[18] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[19] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[20] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[21] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[22] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[23] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[24] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[25] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[26] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore5[27] <= Weights5[(32'd621+32'd1)*32'd19-1:32'd621*32'd19];
			WeightsStore6[0] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[1] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[2] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[3] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[4] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[5] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[6] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[7] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[8] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[9] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[10] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[11] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[12] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[13] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[14] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[15] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[16] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[17] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[18] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[19] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[20] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[21] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[22] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[23] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[24] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[25] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[26] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore6[27] <= Weights6[(32'd622+32'd1)*32'd19-1:32'd622*32'd19];
			WeightsStore7[0] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[1] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[2] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[3] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[4] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[5] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[6] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[7] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[8] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[9] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[10] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[11] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[12] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[13] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[14] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[15] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[16] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[17] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[18] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[19] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[20] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[21] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[22] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[23] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[24] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[25] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[26] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore7[27] <= Weights7[(32'd623+32'd1)*32'd19-1:32'd623*32'd19];
			WeightsStore8[0] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[1] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[2] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[3] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[4] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[5] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[6] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[7] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[8] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[9] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[10] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[11] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[12] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[13] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[14] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[15] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[16] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[17] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[18] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[19] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[20] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[21] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[22] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[23] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[24] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[25] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[26] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore8[27] <= Weights8[(32'd624+32'd1)*32'd19-1:32'd624*32'd19];
			WeightsStore9[0] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[1] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[2] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[3] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[4] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[5] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[6] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[7] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[8] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[9] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[10] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[11] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[12] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[13] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[14] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[15] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[16] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[17] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[18] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[19] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[20] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[21] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[22] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[23] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[24] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[25] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[26] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
			WeightsStore9[27] <= Weights9[(32'd625+32'd1)*32'd19-1:32'd625*32'd19];
		end else if(switchCounter == 32'd23)begin
			PixelsStore[0] <= Pixels[(32'd644+32'd1)*32'd10-1:32'd644*32'd10];
			PixelsStore[1] <= Pixels[(32'd645+32'd1)*32'd10-1:32'd645*32'd10];
			PixelsStore[2] <= Pixels[(32'd646+32'd1)*32'd10-1:32'd646*32'd10];
			PixelsStore[3] <= Pixels[(32'd647+32'd1)*32'd10-1:32'd647*32'd10];
			PixelsStore[4] <= Pixels[(32'd648+32'd1)*32'd10-1:32'd648*32'd10];
			PixelsStore[5] <= Pixels[(32'd649+32'd1)*32'd10-1:32'd649*32'd10];
			PixelsStore[6] <= Pixels[(32'd650+32'd1)*32'd10-1:32'd650*32'd10];
			PixelsStore[7] <= Pixels[(32'd651+32'd1)*32'd10-1:32'd651*32'd10];
			PixelsStore[8] <= Pixels[(32'd652+32'd1)*32'd10-1:32'd652*32'd10];
			PixelsStore[9] <= Pixels[(32'd653+32'd1)*32'd10-1:32'd653*32'd10];
			PixelsStore[10] <= Pixels[(32'd654+32'd1)*32'd10-1:32'd654*32'd10];
			PixelsStore[11] <= Pixels[(32'd655+32'd1)*32'd10-1:32'd655*32'd10];
			PixelsStore[12] <= Pixels[(32'd656+32'd1)*32'd10-1:32'd656*32'd10];
			PixelsStore[13] <= Pixels[(32'd657+32'd1)*32'd10-1:32'd657*32'd10];
			PixelsStore[14] <= Pixels[(32'd658+32'd1)*32'd10-1:32'd658*32'd10];
			PixelsStore[15] <= Pixels[(32'd659+32'd1)*32'd10-1:32'd659*32'd10];
			PixelsStore[16] <= Pixels[(32'd660+32'd1)*32'd10-1:32'd660*32'd10];
			PixelsStore[17] <= Pixels[(32'd661+32'd1)*32'd10-1:32'd661*32'd10];
			PixelsStore[18] <= Pixels[(32'd662+32'd1)*32'd10-1:32'd662*32'd10];
			PixelsStore[19] <= Pixels[(32'd663+32'd1)*32'd10-1:32'd663*32'd10];
			PixelsStore[20] <= Pixels[(32'd664+32'd1)*32'd10-1:32'd664*32'd10];
			PixelsStore[21] <= Pixels[(32'd665+32'd1)*32'd10-1:32'd665*32'd10];
			PixelsStore[22] <= Pixels[(32'd666+32'd1)*32'd10-1:32'd666*32'd10];
			PixelsStore[23] <= Pixels[(32'd667+32'd1)*32'd10-1:32'd667*32'd10];
			PixelsStore[24] <= Pixels[(32'd668+32'd1)*32'd10-1:32'd668*32'd10];
			PixelsStore[25] <= Pixels[(32'd669+32'd1)*32'd10-1:32'd669*32'd10];
			PixelsStore[26] <= Pixels[(32'd670+32'd1)*32'd10-1:32'd670*32'd10];
			PixelsStore[27] <= Pixels[(32'd671+32'd1)*32'd10-1:32'd671*32'd10];
			WeightsStore0[0] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[1] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[2] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[3] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[4] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[5] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[6] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[7] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[8] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[9] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[10] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[11] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[12] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[13] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[14] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[15] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[16] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[17] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[18] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[19] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[20] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[21] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[22] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[23] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[24] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[25] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[26] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore0[27] <= Weights0[(32'd644+32'd1)*32'd19-1:32'd644*32'd19];
			WeightsStore1[0] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[1] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[2] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[3] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[4] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[5] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[6] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[7] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[8] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[9] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[10] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[11] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[12] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[13] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[14] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[15] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[16] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[17] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[18] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[19] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[20] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[21] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[22] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[23] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[24] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[25] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[26] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore1[27] <= Weights1[(32'd645+32'd1)*32'd19-1:32'd645*32'd19];
			WeightsStore2[0] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[1] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[2] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[3] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[4] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[5] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[6] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[7] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[8] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[9] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[10] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[11] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[12] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[13] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[14] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[15] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[16] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[17] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[18] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[19] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[20] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[21] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[22] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[23] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[24] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[25] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[26] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore2[27] <= Weights2[(32'd646+32'd1)*32'd19-1:32'd646*32'd19];
			WeightsStore3[0] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[1] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[2] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[3] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[4] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[5] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[6] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[7] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[8] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[9] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[10] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[11] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[12] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[13] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[14] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[15] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[16] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[17] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[18] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[19] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[20] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[21] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[22] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[23] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[24] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[25] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[26] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore3[27] <= Weights3[(32'd647+32'd1)*32'd19-1:32'd647*32'd19];
			WeightsStore4[0] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[1] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[2] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[3] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[4] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[5] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[6] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[7] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[8] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[9] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[10] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[11] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[12] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[13] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[14] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[15] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[16] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[17] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[18] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[19] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[20] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[21] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[22] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[23] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[24] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[25] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[26] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore4[27] <= Weights4[(32'd648+32'd1)*32'd19-1:32'd648*32'd19];
			WeightsStore5[0] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[1] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[2] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[3] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[4] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[5] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[6] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[7] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[8] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[9] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[10] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[11] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[12] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[13] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[14] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[15] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[16] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[17] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[18] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[19] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[20] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[21] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[22] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[23] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[24] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[25] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[26] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore5[27] <= Weights5[(32'd649+32'd1)*32'd19-1:32'd649*32'd19];
			WeightsStore6[0] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[1] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[2] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[3] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[4] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[5] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[6] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[7] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[8] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[9] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[10] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[11] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[12] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[13] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[14] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[15] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[16] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[17] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[18] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[19] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[20] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[21] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[22] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[23] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[24] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[25] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[26] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore6[27] <= Weights6[(32'd650+32'd1)*32'd19-1:32'd650*32'd19];
			WeightsStore7[0] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[1] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[2] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[3] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[4] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[5] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[6] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[7] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[8] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[9] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[10] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[11] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[12] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[13] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[14] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[15] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[16] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[17] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[18] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[19] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[20] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[21] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[22] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[23] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[24] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[25] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[26] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore7[27] <= Weights7[(32'd651+32'd1)*32'd19-1:32'd651*32'd19];
			WeightsStore8[0] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[1] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[2] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[3] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[4] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[5] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[6] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[7] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[8] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[9] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[10] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[11] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[12] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[13] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[14] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[15] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[16] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[17] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[18] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[19] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[20] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[21] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[22] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[23] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[24] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[25] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[26] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore8[27] <= Weights8[(32'd652+32'd1)*32'd19-1:32'd652*32'd19];
			WeightsStore9[0] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[1] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[2] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[3] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[4] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[5] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[6] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[7] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[8] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[9] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[10] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[11] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[12] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[13] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[14] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[15] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[16] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[17] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[18] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[19] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[20] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[21] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[22] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[23] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[24] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[25] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[26] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
			WeightsStore9[27] <= Weights9[(32'd653+32'd1)*32'd19-1:32'd653*32'd19];
		end else if(switchCounter == 32'd24)begin
			PixelsStore[0] <= Pixels[(32'd672+32'd1)*32'd10-1:32'd672*32'd10];
			PixelsStore[1] <= Pixels[(32'd673+32'd1)*32'd10-1:32'd673*32'd10];
			PixelsStore[2] <= Pixels[(32'd674+32'd1)*32'd10-1:32'd674*32'd10];
			PixelsStore[3] <= Pixels[(32'd675+32'd1)*32'd10-1:32'd675*32'd10];
			PixelsStore[4] <= Pixels[(32'd676+32'd1)*32'd10-1:32'd676*32'd10];
			PixelsStore[5] <= Pixels[(32'd677+32'd1)*32'd10-1:32'd677*32'd10];
			PixelsStore[6] <= Pixels[(32'd678+32'd1)*32'd10-1:32'd678*32'd10];
			PixelsStore[7] <= Pixels[(32'd679+32'd1)*32'd10-1:32'd679*32'd10];
			PixelsStore[8] <= Pixels[(32'd680+32'd1)*32'd10-1:32'd680*32'd10];
			PixelsStore[9] <= Pixels[(32'd681+32'd1)*32'd10-1:32'd681*32'd10];
			PixelsStore[10] <= Pixels[(32'd682+32'd1)*32'd10-1:32'd682*32'd10];
			PixelsStore[11] <= Pixels[(32'd683+32'd1)*32'd10-1:32'd683*32'd10];
			PixelsStore[12] <= Pixels[(32'd684+32'd1)*32'd10-1:32'd684*32'd10];
			PixelsStore[13] <= Pixels[(32'd685+32'd1)*32'd10-1:32'd685*32'd10];
			PixelsStore[14] <= Pixels[(32'd686+32'd1)*32'd10-1:32'd686*32'd10];
			PixelsStore[15] <= Pixels[(32'd687+32'd1)*32'd10-1:32'd687*32'd10];
			PixelsStore[16] <= Pixels[(32'd688+32'd1)*32'd10-1:32'd688*32'd10];
			PixelsStore[17] <= Pixels[(32'd689+32'd1)*32'd10-1:32'd689*32'd10];
			PixelsStore[18] <= Pixels[(32'd690+32'd1)*32'd10-1:32'd690*32'd10];
			PixelsStore[19] <= Pixels[(32'd691+32'd1)*32'd10-1:32'd691*32'd10];
			PixelsStore[20] <= Pixels[(32'd692+32'd1)*32'd10-1:32'd692*32'd10];
			PixelsStore[21] <= Pixels[(32'd693+32'd1)*32'd10-1:32'd693*32'd10];
			PixelsStore[22] <= Pixels[(32'd694+32'd1)*32'd10-1:32'd694*32'd10];
			PixelsStore[23] <= Pixels[(32'd695+32'd1)*32'd10-1:32'd695*32'd10];
			PixelsStore[24] <= Pixels[(32'd696+32'd1)*32'd10-1:32'd696*32'd10];
			PixelsStore[25] <= Pixels[(32'd697+32'd1)*32'd10-1:32'd697*32'd10];
			PixelsStore[26] <= Pixels[(32'd698+32'd1)*32'd10-1:32'd698*32'd10];
			PixelsStore[27] <= Pixels[(32'd699+32'd1)*32'd10-1:32'd699*32'd10];
			WeightsStore0[0] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[1] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[2] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[3] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[4] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[5] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[6] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[7] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[8] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[9] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[10] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[11] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[12] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[13] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[14] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[15] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[16] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[17] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[18] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[19] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[20] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[21] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[22] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[23] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[24] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[25] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[26] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore0[27] <= Weights0[(32'd672+32'd1)*32'd19-1:32'd672*32'd19];
			WeightsStore1[0] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[1] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[2] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[3] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[4] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[5] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[6] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[7] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[8] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[9] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[10] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[11] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[12] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[13] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[14] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[15] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[16] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[17] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[18] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[19] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[20] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[21] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[22] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[23] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[24] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[25] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[26] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore1[27] <= Weights1[(32'd673+32'd1)*32'd19-1:32'd673*32'd19];
			WeightsStore2[0] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[1] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[2] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[3] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[4] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[5] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[6] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[7] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[8] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[9] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[10] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[11] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[12] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[13] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[14] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[15] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[16] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[17] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[18] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[19] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[20] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[21] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[22] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[23] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[24] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[25] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[26] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore2[27] <= Weights2[(32'd674+32'd1)*32'd19-1:32'd674*32'd19];
			WeightsStore3[0] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[1] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[2] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[3] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[4] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[5] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[6] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[7] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[8] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[9] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[10] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[11] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[12] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[13] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[14] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[15] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[16] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[17] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[18] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[19] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[20] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[21] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[22] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[23] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[24] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[25] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[26] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore3[27] <= Weights3[(32'd675+32'd1)*32'd19-1:32'd675*32'd19];
			WeightsStore4[0] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[1] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[2] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[3] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[4] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[5] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[6] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[7] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[8] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[9] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[10] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[11] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[12] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[13] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[14] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[15] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[16] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[17] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[18] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[19] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[20] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[21] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[22] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[23] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[24] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[25] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[26] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore4[27] <= Weights4[(32'd676+32'd1)*32'd19-1:32'd676*32'd19];
			WeightsStore5[0] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[1] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[2] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[3] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[4] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[5] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[6] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[7] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[8] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[9] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[10] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[11] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[12] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[13] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[14] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[15] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[16] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[17] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[18] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[19] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[20] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[21] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[22] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[23] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[24] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[25] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[26] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore5[27] <= Weights5[(32'd677+32'd1)*32'd19-1:32'd677*32'd19];
			WeightsStore6[0] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[1] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[2] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[3] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[4] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[5] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[6] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[7] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[8] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[9] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[10] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[11] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[12] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[13] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[14] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[15] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[16] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[17] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[18] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[19] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[20] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[21] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[22] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[23] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[24] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[25] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[26] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore6[27] <= Weights6[(32'd678+32'd1)*32'd19-1:32'd678*32'd19];
			WeightsStore7[0] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[1] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[2] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[3] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[4] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[5] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[6] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[7] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[8] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[9] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[10] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[11] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[12] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[13] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[14] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[15] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[16] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[17] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[18] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[19] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[20] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[21] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[22] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[23] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[24] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[25] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[26] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore7[27] <= Weights7[(32'd679+32'd1)*32'd19-1:32'd679*32'd19];
			WeightsStore8[0] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[1] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[2] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[3] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[4] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[5] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[6] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[7] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[8] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[9] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[10] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[11] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[12] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[13] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[14] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[15] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[16] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[17] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[18] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[19] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[20] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[21] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[22] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[23] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[24] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[25] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[26] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore8[27] <= Weights8[(32'd680+32'd1)*32'd19-1:32'd680*32'd19];
			WeightsStore9[0] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[1] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[2] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[3] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[4] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[5] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[6] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[7] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[8] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[9] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[10] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[11] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[12] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[13] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[14] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[15] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[16] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[17] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[18] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[19] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[20] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[21] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[22] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[23] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[24] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[25] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[26] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
			WeightsStore9[27] <= Weights9[(32'd681+32'd1)*32'd19-1:32'd681*32'd19];
		end else if(switchCounter == 32'd25)begin
			PixelsStore[0] <= Pixels[(32'd700+32'd1)*32'd10-1:32'd700*32'd10];
			PixelsStore[1] <= Pixels[(32'd701+32'd1)*32'd10-1:32'd701*32'd10];
			PixelsStore[2] <= Pixels[(32'd702+32'd1)*32'd10-1:32'd702*32'd10];
			PixelsStore[3] <= Pixels[(32'd703+32'd1)*32'd10-1:32'd703*32'd10];
			PixelsStore[4] <= Pixels[(32'd704+32'd1)*32'd10-1:32'd704*32'd10];
			PixelsStore[5] <= Pixels[(32'd705+32'd1)*32'd10-1:32'd705*32'd10];
			PixelsStore[6] <= Pixels[(32'd706+32'd1)*32'd10-1:32'd706*32'd10];
			PixelsStore[7] <= Pixels[(32'd707+32'd1)*32'd10-1:32'd707*32'd10];
			PixelsStore[8] <= Pixels[(32'd708+32'd1)*32'd10-1:32'd708*32'd10];
			PixelsStore[9] <= Pixels[(32'd709+32'd1)*32'd10-1:32'd709*32'd10];
			PixelsStore[10] <= Pixels[(32'd710+32'd1)*32'd10-1:32'd710*32'd10];
			PixelsStore[11] <= Pixels[(32'd711+32'd1)*32'd10-1:32'd711*32'd10];
			PixelsStore[12] <= Pixels[(32'd712+32'd1)*32'd10-1:32'd712*32'd10];
			PixelsStore[13] <= Pixels[(32'd713+32'd1)*32'd10-1:32'd713*32'd10];
			PixelsStore[14] <= Pixels[(32'd714+32'd1)*32'd10-1:32'd714*32'd10];
			PixelsStore[15] <= Pixels[(32'd715+32'd1)*32'd10-1:32'd715*32'd10];
			PixelsStore[16] <= Pixels[(32'd716+32'd1)*32'd10-1:32'd716*32'd10];
			PixelsStore[17] <= Pixels[(32'd717+32'd1)*32'd10-1:32'd717*32'd10];
			PixelsStore[18] <= Pixels[(32'd718+32'd1)*32'd10-1:32'd718*32'd10];
			PixelsStore[19] <= Pixels[(32'd719+32'd1)*32'd10-1:32'd719*32'd10];
			PixelsStore[20] <= Pixels[(32'd720+32'd1)*32'd10-1:32'd720*32'd10];
			PixelsStore[21] <= Pixels[(32'd721+32'd1)*32'd10-1:32'd721*32'd10];
			PixelsStore[22] <= Pixels[(32'd722+32'd1)*32'd10-1:32'd722*32'd10];
			PixelsStore[23] <= Pixels[(32'd723+32'd1)*32'd10-1:32'd723*32'd10];
			PixelsStore[24] <= Pixels[(32'd724+32'd1)*32'd10-1:32'd724*32'd10];
			PixelsStore[25] <= Pixels[(32'd725+32'd1)*32'd10-1:32'd725*32'd10];
			PixelsStore[26] <= Pixels[(32'd726+32'd1)*32'd10-1:32'd726*32'd10];
			PixelsStore[27] <= Pixels[(32'd727+32'd1)*32'd10-1:32'd727*32'd10];
			WeightsStore0[0] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[1] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[2] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[3] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[4] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[5] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[6] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[7] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[8] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[9] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[10] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[11] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[12] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[13] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[14] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[15] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[16] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[17] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[18] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[19] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[20] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[21] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[22] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[23] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[24] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[25] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[26] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore0[27] <= Weights0[(32'd700+32'd1)*32'd19-1:32'd700*32'd19];
			WeightsStore1[0] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[1] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[2] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[3] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[4] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[5] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[6] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[7] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[8] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[9] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[10] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[11] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[12] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[13] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[14] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[15] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[16] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[17] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[18] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[19] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[20] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[21] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[22] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[23] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[24] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[25] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[26] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore1[27] <= Weights1[(32'd701+32'd1)*32'd19-1:32'd701*32'd19];
			WeightsStore2[0] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[1] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[2] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[3] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[4] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[5] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[6] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[7] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[8] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[9] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[10] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[11] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[12] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[13] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[14] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[15] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[16] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[17] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[18] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[19] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[20] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[21] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[22] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[23] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[24] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[25] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[26] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore2[27] <= Weights2[(32'd702+32'd1)*32'd19-1:32'd702*32'd19];
			WeightsStore3[0] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[1] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[2] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[3] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[4] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[5] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[6] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[7] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[8] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[9] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[10] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[11] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[12] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[13] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[14] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[15] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[16] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[17] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[18] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[19] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[20] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[21] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[22] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[23] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[24] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[25] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[26] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore3[27] <= Weights3[(32'd703+32'd1)*32'd19-1:32'd703*32'd19];
			WeightsStore4[0] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[1] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[2] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[3] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[4] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[5] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[6] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[7] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[8] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[9] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[10] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[11] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[12] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[13] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[14] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[15] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[16] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[17] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[18] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[19] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[20] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[21] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[22] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[23] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[24] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[25] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[26] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore4[27] <= Weights4[(32'd704+32'd1)*32'd19-1:32'd704*32'd19];
			WeightsStore5[0] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[1] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[2] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[3] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[4] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[5] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[6] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[7] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[8] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[9] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[10] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[11] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[12] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[13] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[14] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[15] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[16] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[17] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[18] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[19] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[20] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[21] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[22] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[23] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[24] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[25] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[26] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore5[27] <= Weights5[(32'd705+32'd1)*32'd19-1:32'd705*32'd19];
			WeightsStore6[0] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[1] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[2] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[3] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[4] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[5] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[6] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[7] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[8] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[9] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[10] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[11] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[12] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[13] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[14] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[15] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[16] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[17] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[18] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[19] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[20] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[21] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[22] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[23] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[24] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[25] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[26] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore6[27] <= Weights6[(32'd706+32'd1)*32'd19-1:32'd706*32'd19];
			WeightsStore7[0] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[1] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[2] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[3] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[4] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[5] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[6] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[7] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[8] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[9] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[10] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[11] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[12] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[13] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[14] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[15] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[16] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[17] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[18] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[19] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[20] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[21] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[22] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[23] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[24] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[25] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[26] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore7[27] <= Weights7[(32'd707+32'd1)*32'd19-1:32'd707*32'd19];
			WeightsStore8[0] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[1] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[2] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[3] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[4] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[5] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[6] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[7] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[8] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[9] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[10] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[11] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[12] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[13] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[14] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[15] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[16] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[17] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[18] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[19] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[20] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[21] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[22] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[23] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[24] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[25] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[26] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore8[27] <= Weights8[(32'd708+32'd1)*32'd19-1:32'd708*32'd19];
			WeightsStore9[0] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[1] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[2] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[3] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[4] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[5] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[6] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[7] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[8] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[9] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[10] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[11] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[12] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[13] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[14] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[15] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[16] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[17] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[18] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[19] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[20] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[21] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[22] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[23] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[24] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[25] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[26] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
			WeightsStore9[27] <= Weights9[(32'd709+32'd1)*32'd19-1:32'd709*32'd19];
		end else if(switchCounter == 32'd26)begin
			PixelsStore[0] <= Pixels[(32'd728+32'd1)*32'd10-1:32'd728*32'd10];
			PixelsStore[1] <= Pixels[(32'd729+32'd1)*32'd10-1:32'd729*32'd10];
			PixelsStore[2] <= Pixels[(32'd730+32'd1)*32'd10-1:32'd730*32'd10];
			PixelsStore[3] <= Pixels[(32'd731+32'd1)*32'd10-1:32'd731*32'd10];
			PixelsStore[4] <= Pixels[(32'd732+32'd1)*32'd10-1:32'd732*32'd10];
			PixelsStore[5] <= Pixels[(32'd733+32'd1)*32'd10-1:32'd733*32'd10];
			PixelsStore[6] <= Pixels[(32'd734+32'd1)*32'd10-1:32'd734*32'd10];
			PixelsStore[7] <= Pixels[(32'd735+32'd1)*32'd10-1:32'd735*32'd10];
			PixelsStore[8] <= Pixels[(32'd736+32'd1)*32'd10-1:32'd736*32'd10];
			PixelsStore[9] <= Pixels[(32'd737+32'd1)*32'd10-1:32'd737*32'd10];
			PixelsStore[10] <= Pixels[(32'd738+32'd1)*32'd10-1:32'd738*32'd10];
			PixelsStore[11] <= Pixels[(32'd739+32'd1)*32'd10-1:32'd739*32'd10];
			PixelsStore[12] <= Pixels[(32'd740+32'd1)*32'd10-1:32'd740*32'd10];
			PixelsStore[13] <= Pixels[(32'd741+32'd1)*32'd10-1:32'd741*32'd10];
			PixelsStore[14] <= Pixels[(32'd742+32'd1)*32'd10-1:32'd742*32'd10];
			PixelsStore[15] <= Pixels[(32'd743+32'd1)*32'd10-1:32'd743*32'd10];
			PixelsStore[16] <= Pixels[(32'd744+32'd1)*32'd10-1:32'd744*32'd10];
			PixelsStore[17] <= Pixels[(32'd745+32'd1)*32'd10-1:32'd745*32'd10];
			PixelsStore[18] <= Pixels[(32'd746+32'd1)*32'd10-1:32'd746*32'd10];
			PixelsStore[19] <= Pixels[(32'd747+32'd1)*32'd10-1:32'd747*32'd10];
			PixelsStore[20] <= Pixels[(32'd748+32'd1)*32'd10-1:32'd748*32'd10];
			PixelsStore[21] <= Pixels[(32'd749+32'd1)*32'd10-1:32'd749*32'd10];
			PixelsStore[22] <= Pixels[(32'd750+32'd1)*32'd10-1:32'd750*32'd10];
			PixelsStore[23] <= Pixels[(32'd751+32'd1)*32'd10-1:32'd751*32'd10];
			PixelsStore[24] <= Pixels[(32'd752+32'd1)*32'd10-1:32'd752*32'd10];
			PixelsStore[25] <= Pixels[(32'd753+32'd1)*32'd10-1:32'd753*32'd10];
			PixelsStore[26] <= Pixels[(32'd754+32'd1)*32'd10-1:32'd754*32'd10];
			PixelsStore[27] <= Pixels[(32'd755+32'd1)*32'd10-1:32'd755*32'd10];
			WeightsStore0[0] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[1] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[2] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[3] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[4] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[5] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[6] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[7] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[8] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[9] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[10] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[11] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[12] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[13] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[14] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[15] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[16] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[17] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[18] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[19] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[20] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[21] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[22] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[23] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[24] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[25] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[26] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore0[27] <= Weights0[(32'd728+32'd1)*32'd19-1:32'd728*32'd19];
			WeightsStore1[0] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[1] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[2] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[3] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[4] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[5] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[6] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[7] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[8] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[9] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[10] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[11] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[12] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[13] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[14] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[15] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[16] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[17] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[18] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[19] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[20] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[21] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[22] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[23] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[24] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[25] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[26] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore1[27] <= Weights1[(32'd729+32'd1)*32'd19-1:32'd729*32'd19];
			WeightsStore2[0] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[1] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[2] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[3] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[4] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[5] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[6] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[7] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[8] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[9] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[10] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[11] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[12] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[13] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[14] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[15] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[16] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[17] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[18] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[19] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[20] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[21] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[22] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[23] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[24] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[25] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[26] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore2[27] <= Weights2[(32'd730+32'd1)*32'd19-1:32'd730*32'd19];
			WeightsStore3[0] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[1] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[2] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[3] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[4] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[5] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[6] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[7] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[8] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[9] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[10] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[11] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[12] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[13] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[14] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[15] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[16] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[17] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[18] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[19] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[20] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[21] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[22] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[23] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[24] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[25] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[26] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore3[27] <= Weights3[(32'd731+32'd1)*32'd19-1:32'd731*32'd19];
			WeightsStore4[0] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[1] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[2] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[3] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[4] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[5] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[6] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[7] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[8] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[9] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[10] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[11] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[12] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[13] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[14] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[15] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[16] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[17] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[18] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[19] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[20] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[21] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[22] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[23] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[24] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[25] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[26] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore4[27] <= Weights4[(32'd732+32'd1)*32'd19-1:32'd732*32'd19];
			WeightsStore5[0] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[1] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[2] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[3] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[4] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[5] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[6] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[7] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[8] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[9] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[10] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[11] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[12] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[13] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[14] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[15] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[16] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[17] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[18] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[19] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[20] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[21] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[22] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[23] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[24] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[25] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[26] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore5[27] <= Weights5[(32'd733+32'd1)*32'd19-1:32'd733*32'd19];
			WeightsStore6[0] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[1] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[2] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[3] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[4] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[5] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[6] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[7] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[8] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[9] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[10] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[11] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[12] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[13] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[14] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[15] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[16] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[17] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[18] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[19] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[20] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[21] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[22] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[23] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[24] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[25] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[26] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore6[27] <= Weights6[(32'd734+32'd1)*32'd19-1:32'd734*32'd19];
			WeightsStore7[0] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[1] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[2] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[3] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[4] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[5] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[6] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[7] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[8] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[9] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[10] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[11] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[12] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[13] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[14] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[15] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[16] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[17] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[18] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[19] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[20] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[21] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[22] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[23] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[24] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[25] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[26] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore7[27] <= Weights7[(32'd735+32'd1)*32'd19-1:32'd735*32'd19];
			WeightsStore8[0] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[1] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[2] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[3] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[4] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[5] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[6] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[7] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[8] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[9] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[10] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[11] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[12] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[13] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[14] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[15] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[16] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[17] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[18] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[19] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[20] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[21] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[22] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[23] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[24] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[25] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[26] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore8[27] <= Weights8[(32'd736+32'd1)*32'd19-1:32'd736*32'd19];
			WeightsStore9[0] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[1] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[2] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[3] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[4] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[5] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[6] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[7] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[8] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[9] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[10] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[11] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[12] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[13] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[14] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[15] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[16] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[17] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[18] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[19] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[20] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[21] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[22] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[23] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[24] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[25] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[26] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
			WeightsStore9[27] <= Weights9[(32'd737+32'd1)*32'd19-1:32'd737*32'd19];
		end else if(switchCounter == 32'd27)begin
			PixelsStore[0] <= Pixels[(32'd756+32'd1)*32'd10-1:32'd756*32'd10];
			PixelsStore[1] <= Pixels[(32'd757+32'd1)*32'd10-1:32'd757*32'd10];
			PixelsStore[2] <= Pixels[(32'd758+32'd1)*32'd10-1:32'd758*32'd10];
			PixelsStore[3] <= Pixels[(32'd759+32'd1)*32'd10-1:32'd759*32'd10];
			PixelsStore[4] <= Pixels[(32'd760+32'd1)*32'd10-1:32'd760*32'd10];
			PixelsStore[5] <= Pixels[(32'd761+32'd1)*32'd10-1:32'd761*32'd10];
			PixelsStore[6] <= Pixels[(32'd762+32'd1)*32'd10-1:32'd762*32'd10];
			PixelsStore[7] <= Pixels[(32'd763+32'd1)*32'd10-1:32'd763*32'd10];
			PixelsStore[8] <= Pixels[(32'd764+32'd1)*32'd10-1:32'd764*32'd10];
			PixelsStore[9] <= Pixels[(32'd765+32'd1)*32'd10-1:32'd765*32'd10];
			PixelsStore[10] <= Pixels[(32'd766+32'd1)*32'd10-1:32'd766*32'd10];
			PixelsStore[11] <= Pixels[(32'd767+32'd1)*32'd10-1:32'd767*32'd10];
			PixelsStore[12] <= Pixels[(32'd768+32'd1)*32'd10-1:32'd768*32'd10];
			PixelsStore[13] <= Pixels[(32'd769+32'd1)*32'd10-1:32'd769*32'd10];
			PixelsStore[14] <= Pixels[(32'd770+32'd1)*32'd10-1:32'd770*32'd10];
			PixelsStore[15] <= Pixels[(32'd771+32'd1)*32'd10-1:32'd771*32'd10];
			PixelsStore[16] <= Pixels[(32'd772+32'd1)*32'd10-1:32'd772*32'd10];
			PixelsStore[17] <= Pixels[(32'd773+32'd1)*32'd10-1:32'd773*32'd10];
			PixelsStore[18] <= Pixels[(32'd774+32'd1)*32'd10-1:32'd774*32'd10];
			PixelsStore[19] <= Pixels[(32'd775+32'd1)*32'd10-1:32'd775*32'd10];
			PixelsStore[20] <= Pixels[(32'd776+32'd1)*32'd10-1:32'd776*32'd10];
			PixelsStore[21] <= Pixels[(32'd777+32'd1)*32'd10-1:32'd777*32'd10];
			PixelsStore[22] <= Pixels[(32'd778+32'd1)*32'd10-1:32'd778*32'd10];
			PixelsStore[23] <= Pixels[(32'd779+32'd1)*32'd10-1:32'd779*32'd10];
			PixelsStore[24] <= Pixels[(32'd780+32'd1)*32'd10-1:32'd780*32'd10];
			PixelsStore[25] <= Pixels[(32'd781+32'd1)*32'd10-1:32'd781*32'd10];
			PixelsStore[26] <= Pixels[(32'd782+32'd1)*32'd10-1:32'd782*32'd10];
			PixelsStore[27] <= Pixels[(32'd783+32'd1)*32'd10-1:32'd783*32'd10];
			WeightsStore0[0] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[1] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[2] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[3] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[4] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[5] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[6] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[7] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[8] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[9] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[10] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[11] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[12] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[13] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[14] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[15] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[16] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[17] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[18] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[19] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[20] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[21] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[22] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[23] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[24] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[25] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[26] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore0[27] <= Weights0[(32'd756+32'd1)*32'd19-1:32'd756*32'd19];
			WeightsStore1[0] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[1] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[2] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[3] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[4] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[5] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[6] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[7] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[8] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[9] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[10] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[11] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[12] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[13] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[14] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[15] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[16] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[17] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[18] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[19] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[20] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[21] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[22] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[23] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[24] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[25] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[26] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore1[27] <= Weights1[(32'd757+32'd1)*32'd19-1:32'd757*32'd19];
			WeightsStore2[0] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[1] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[2] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[3] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[4] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[5] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[6] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[7] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[8] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[9] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[10] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[11] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[12] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[13] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[14] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[15] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[16] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[17] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[18] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[19] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[20] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[21] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[22] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[23] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[24] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[25] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[26] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore2[27] <= Weights2[(32'd758+32'd1)*32'd19-1:32'd758*32'd19];
			WeightsStore3[0] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[1] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[2] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[3] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[4] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[5] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[6] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[7] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[8] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[9] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[10] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[11] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[12] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[13] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[14] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[15] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[16] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[17] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[18] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[19] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[20] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[21] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[22] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[23] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[24] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[25] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[26] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore3[27] <= Weights3[(32'd759+32'd1)*32'd19-1:32'd759*32'd19];
			WeightsStore4[0] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[1] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[2] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[3] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[4] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[5] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[6] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[7] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[8] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[9] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[10] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[11] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[12] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[13] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[14] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[15] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[16] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[17] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[18] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[19] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[20] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[21] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[22] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[23] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[24] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[25] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[26] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore4[27] <= Weights4[(32'd760+32'd1)*32'd19-1:32'd760*32'd19];
			WeightsStore5[0] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[1] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[2] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[3] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[4] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[5] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[6] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[7] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[8] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[9] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[10] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[11] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[12] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[13] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[14] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[15] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[16] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[17] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[18] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[19] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[20] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[21] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[22] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[23] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[24] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[25] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[26] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore5[27] <= Weights5[(32'd761+32'd1)*32'd19-1:32'd761*32'd19];
			WeightsStore6[0] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[1] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[2] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[3] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[4] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[5] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[6] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[7] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[8] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[9] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[10] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[11] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[12] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[13] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[14] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[15] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[16] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[17] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[18] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[19] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[20] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[21] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[22] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[23] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[24] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[25] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[26] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore6[27] <= Weights6[(32'd762+32'd1)*32'd19-1:32'd762*32'd19];
			WeightsStore7[0] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[1] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[2] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[3] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[4] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[5] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[6] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[7] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[8] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[9] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[10] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[11] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[12] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[13] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[14] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[15] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[16] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[17] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[18] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[19] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[20] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[21] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[22] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[23] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[24] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[25] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[26] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore7[27] <= Weights7[(32'd763+32'd1)*32'd19-1:32'd763*32'd19];
			WeightsStore8[0] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[1] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[2] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[3] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[4] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[5] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[6] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[7] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[8] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[9] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[10] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[11] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[12] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[13] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[14] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[15] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[16] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[17] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[18] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[19] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[20] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[21] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[22] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[23] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[24] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[25] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[26] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore8[27] <= Weights8[(32'd764+32'd1)*32'd19-1:32'd764*32'd19];
			WeightsStore9[0] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[1] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[2] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[3] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[4] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[5] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[6] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[7] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[8] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[9] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[10] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[11] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[12] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[13] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[14] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[15] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[16] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[17] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[18] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[19] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[20] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[21] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[22] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[23] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[24] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[25] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[26] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
			WeightsStore9[27] <= Weights9[(32'd765+32'd1)*32'd19-1:32'd765*32'd19];
		end
		switchCounter <= switchCounter + 32'd1;
	end
end

endmodule
