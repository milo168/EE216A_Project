module Image_Classifier
#(parameter NEURONS = 10,
  parameter PIXEL_N = 785,
  parameter WEIGHT_SIZE = 19,
  parameter PIXEL_SIZE = 10,
  parameter FPM_DELAY = 6,
  parameter FPA_DELAY = 2,
  parameter PARALLEL = 2,
  parameter BUS_WIDTH = 1,
  parameter VAL_SIZE = 26)
(
input clk,
input GlobalReset,
input Input_Valid,
input [WEIGHT_SIZE-1:0] Wgt_0_0,input [WEIGHT_SIZE-1:0] Wgt_0_1,input [WEIGHT_SIZE-1:0] Wgt_0_2,input [WEIGHT_SIZE-1:0] Wgt_0_3,input [WEIGHT_SIZE-1:0] Wgt_0_4,input [WEIGHT_SIZE-1:0] Wgt_0_5,input [WEIGHT_SIZE-1:0] Wgt_0_6,input [WEIGHT_SIZE-1:0] Wgt_0_7,input [WEIGHT_SIZE-1:0] Wgt_0_8,input [WEIGHT_SIZE-1:0] Wgt_0_9,input [WEIGHT_SIZE-1:0] Wgt_0_10,input [WEIGHT_SIZE-1:0] Wgt_0_11,input [WEIGHT_SIZE-1:0] Wgt_0_12,input [WEIGHT_SIZE-1:0] Wgt_0_13,input [WEIGHT_SIZE-1:0] Wgt_0_14,input [WEIGHT_SIZE-1:0] Wgt_0_15,input [WEIGHT_SIZE-1:0] Wgt_0_16,input [WEIGHT_SIZE-1:0] Wgt_0_17,input [WEIGHT_SIZE-1:0] Wgt_0_18,input [WEIGHT_SIZE-1:0] Wgt_0_19,input [WEIGHT_SIZE-1:0] Wgt_0_20,input [WEIGHT_SIZE-1:0] Wgt_0_21,input [WEIGHT_SIZE-1:0] Wgt_0_22,input [WEIGHT_SIZE-1:0] Wgt_0_23,input [WEIGHT_SIZE-1:0] Wgt_0_24,input [WEIGHT_SIZE-1:0] Wgt_0_25,input [WEIGHT_SIZE-1:0] Wgt_0_26,input [WEIGHT_SIZE-1:0] Wgt_0_27,input [WEIGHT_SIZE-1:0] Wgt_0_28,input [WEIGHT_SIZE-1:0] Wgt_0_29,input [WEIGHT_SIZE-1:0] Wgt_0_30,input [WEIGHT_SIZE-1:0] Wgt_0_31,input [WEIGHT_SIZE-1:0] Wgt_0_32,input [WEIGHT_SIZE-1:0] Wgt_0_33,input [WEIGHT_SIZE-1:0] Wgt_0_34,input [WEIGHT_SIZE-1:0] Wgt_0_35,input [WEIGHT_SIZE-1:0] Wgt_0_36,input [WEIGHT_SIZE-1:0] Wgt_0_37,input [WEIGHT_SIZE-1:0] Wgt_0_38,input [WEIGHT_SIZE-1:0] Wgt_0_39,input [WEIGHT_SIZE-1:0] Wgt_0_40,input [WEIGHT_SIZE-1:0] Wgt_0_41,input [WEIGHT_SIZE-1:0] Wgt_0_42,input [WEIGHT_SIZE-1:0] Wgt_0_43,input [WEIGHT_SIZE-1:0] Wgt_0_44,input [WEIGHT_SIZE-1:0] Wgt_0_45,input [WEIGHT_SIZE-1:0] Wgt_0_46,input [WEIGHT_SIZE-1:0] Wgt_0_47,input [WEIGHT_SIZE-1:0] Wgt_0_48,input [WEIGHT_SIZE-1:0] Wgt_0_49,input [WEIGHT_SIZE-1:0] Wgt_0_50,input [WEIGHT_SIZE-1:0] Wgt_0_51,input [WEIGHT_SIZE-1:0] Wgt_0_52,input [WEIGHT_SIZE-1:0] Wgt_0_53,input [WEIGHT_SIZE-1:0] Wgt_0_54,input [WEIGHT_SIZE-1:0] Wgt_0_55,input [WEIGHT_SIZE-1:0] Wgt_0_56,input [WEIGHT_SIZE-1:0] Wgt_0_57,input [WEIGHT_SIZE-1:0] Wgt_0_58,input [WEIGHT_SIZE-1:0] Wgt_0_59,input [WEIGHT_SIZE-1:0] Wgt_0_60,input [WEIGHT_SIZE-1:0] Wgt_0_61,input [WEIGHT_SIZE-1:0] Wgt_0_62,input [WEIGHT_SIZE-1:0] Wgt_0_63,input [WEIGHT_SIZE-1:0] Wgt_0_64,input [WEIGHT_SIZE-1:0] Wgt_0_65,input [WEIGHT_SIZE-1:0] Wgt_0_66,input [WEIGHT_SIZE-1:0] Wgt_0_67,input [WEIGHT_SIZE-1:0] Wgt_0_68,input [WEIGHT_SIZE-1:0] Wgt_0_69,input [WEIGHT_SIZE-1:0] Wgt_0_70,input [WEIGHT_SIZE-1:0] Wgt_0_71,input [WEIGHT_SIZE-1:0] Wgt_0_72,input [WEIGHT_SIZE-1:0] Wgt_0_73,input [WEIGHT_SIZE-1:0] Wgt_0_74,input [WEIGHT_SIZE-1:0] Wgt_0_75,input [WEIGHT_SIZE-1:0] Wgt_0_76,input [WEIGHT_SIZE-1:0] Wgt_0_77,input [WEIGHT_SIZE-1:0] Wgt_0_78,input [WEIGHT_SIZE-1:0] Wgt_0_79,input [WEIGHT_SIZE-1:0] Wgt_0_80,input [WEIGHT_SIZE-1:0] Wgt_0_81,input [WEIGHT_SIZE-1:0] Wgt_0_82,input [WEIGHT_SIZE-1:0] Wgt_0_83,input [WEIGHT_SIZE-1:0] Wgt_0_84,input [WEIGHT_SIZE-1:0] Wgt_0_85,input [WEIGHT_SIZE-1:0] Wgt_0_86,input [WEIGHT_SIZE-1:0] Wgt_0_87,input [WEIGHT_SIZE-1:0] Wgt_0_88,input [WEIGHT_SIZE-1:0] Wgt_0_89,input [WEIGHT_SIZE-1:0] Wgt_0_90,input [WEIGHT_SIZE-1:0] Wgt_0_91,input [WEIGHT_SIZE-1:0] Wgt_0_92,input [WEIGHT_SIZE-1:0] Wgt_0_93,input [WEIGHT_SIZE-1:0] Wgt_0_94,input [WEIGHT_SIZE-1:0] Wgt_0_95,input [WEIGHT_SIZE-1:0] Wgt_0_96,input [WEIGHT_SIZE-1:0] Wgt_0_97,input [WEIGHT_SIZE-1:0] Wgt_0_98,input [WEIGHT_SIZE-1:0] Wgt_0_99,input [WEIGHT_SIZE-1:0] Wgt_0_100,input [WEIGHT_SIZE-1:0] Wgt_0_101,input [WEIGHT_SIZE-1:0] Wgt_0_102,input [WEIGHT_SIZE-1:0] Wgt_0_103,input [WEIGHT_SIZE-1:0] Wgt_0_104,input [WEIGHT_SIZE-1:0] Wgt_0_105,input [WEIGHT_SIZE-1:0] Wgt_0_106,input [WEIGHT_SIZE-1:0] Wgt_0_107,input [WEIGHT_SIZE-1:0] Wgt_0_108,input [WEIGHT_SIZE-1:0] Wgt_0_109,input [WEIGHT_SIZE-1:0] Wgt_0_110,input [WEIGHT_SIZE-1:0] Wgt_0_111,input [WEIGHT_SIZE-1:0] Wgt_0_112,input [WEIGHT_SIZE-1:0] Wgt_0_113,input [WEIGHT_SIZE-1:0] Wgt_0_114,input [WEIGHT_SIZE-1:0] Wgt_0_115,input [WEIGHT_SIZE-1:0] Wgt_0_116,input [WEIGHT_SIZE-1:0] Wgt_0_117,input [WEIGHT_SIZE-1:0] Wgt_0_118,input [WEIGHT_SIZE-1:0] Wgt_0_119,input [WEIGHT_SIZE-1:0] Wgt_0_120,input [WEIGHT_SIZE-1:0] Wgt_0_121,input [WEIGHT_SIZE-1:0] Wgt_0_122,input [WEIGHT_SIZE-1:0] Wgt_0_123,input [WEIGHT_SIZE-1:0] Wgt_0_124,input [WEIGHT_SIZE-1:0] Wgt_0_125,input [WEIGHT_SIZE-1:0] Wgt_0_126,input [WEIGHT_SIZE-1:0] Wgt_0_127,input [WEIGHT_SIZE-1:0] Wgt_0_128,input [WEIGHT_SIZE-1:0] Wgt_0_129,input [WEIGHT_SIZE-1:0] Wgt_0_130,input [WEIGHT_SIZE-1:0] Wgt_0_131,input [WEIGHT_SIZE-1:0] Wgt_0_132,input [WEIGHT_SIZE-1:0] Wgt_0_133,input [WEIGHT_SIZE-1:0] Wgt_0_134,input [WEIGHT_SIZE-1:0] Wgt_0_135,input [WEIGHT_SIZE-1:0] Wgt_0_136,input [WEIGHT_SIZE-1:0] Wgt_0_137,input [WEIGHT_SIZE-1:0] Wgt_0_138,input [WEIGHT_SIZE-1:0] Wgt_0_139,input [WEIGHT_SIZE-1:0] Wgt_0_140,input [WEIGHT_SIZE-1:0] Wgt_0_141,input [WEIGHT_SIZE-1:0] Wgt_0_142,input [WEIGHT_SIZE-1:0] Wgt_0_143,input [WEIGHT_SIZE-1:0] Wgt_0_144,input [WEIGHT_SIZE-1:0] Wgt_0_145,input [WEIGHT_SIZE-1:0] Wgt_0_146,input [WEIGHT_SIZE-1:0] Wgt_0_147,input [WEIGHT_SIZE-1:0] Wgt_0_148,input [WEIGHT_SIZE-1:0] Wgt_0_149,input [WEIGHT_SIZE-1:0] Wgt_0_150,input [WEIGHT_SIZE-1:0] Wgt_0_151,input [WEIGHT_SIZE-1:0] Wgt_0_152,input [WEIGHT_SIZE-1:0] Wgt_0_153,input [WEIGHT_SIZE-1:0] Wgt_0_154,input [WEIGHT_SIZE-1:0] Wgt_0_155,input [WEIGHT_SIZE-1:0] Wgt_0_156,input [WEIGHT_SIZE-1:0] Wgt_0_157,input [WEIGHT_SIZE-1:0] Wgt_0_158,input [WEIGHT_SIZE-1:0] Wgt_0_159,input [WEIGHT_SIZE-1:0] Wgt_0_160,input [WEIGHT_SIZE-1:0] Wgt_0_161,input [WEIGHT_SIZE-1:0] Wgt_0_162,input [WEIGHT_SIZE-1:0] Wgt_0_163,input [WEIGHT_SIZE-1:0] Wgt_0_164,input [WEIGHT_SIZE-1:0] Wgt_0_165,input [WEIGHT_SIZE-1:0] Wgt_0_166,input [WEIGHT_SIZE-1:0] Wgt_0_167,input [WEIGHT_SIZE-1:0] Wgt_0_168,input [WEIGHT_SIZE-1:0] Wgt_0_169,input [WEIGHT_SIZE-1:0] Wgt_0_170,input [WEIGHT_SIZE-1:0] Wgt_0_171,input [WEIGHT_SIZE-1:0] Wgt_0_172,input [WEIGHT_SIZE-1:0] Wgt_0_173,input [WEIGHT_SIZE-1:0] Wgt_0_174,input [WEIGHT_SIZE-1:0] Wgt_0_175,input [WEIGHT_SIZE-1:0] Wgt_0_176,input [WEIGHT_SIZE-1:0] Wgt_0_177,input [WEIGHT_SIZE-1:0] Wgt_0_178,input [WEIGHT_SIZE-1:0] Wgt_0_179,input [WEIGHT_SIZE-1:0] Wgt_0_180,input [WEIGHT_SIZE-1:0] Wgt_0_181,input [WEIGHT_SIZE-1:0] Wgt_0_182,input [WEIGHT_SIZE-1:0] Wgt_0_183,input [WEIGHT_SIZE-1:0] Wgt_0_184,input [WEIGHT_SIZE-1:0] Wgt_0_185,input [WEIGHT_SIZE-1:0] Wgt_0_186,input [WEIGHT_SIZE-1:0] Wgt_0_187,input [WEIGHT_SIZE-1:0] Wgt_0_188,input [WEIGHT_SIZE-1:0] Wgt_0_189,input [WEIGHT_SIZE-1:0] Wgt_0_190,input [WEIGHT_SIZE-1:0] Wgt_0_191,input [WEIGHT_SIZE-1:0] Wgt_0_192,input [WEIGHT_SIZE-1:0] Wgt_0_193,input [WEIGHT_SIZE-1:0] Wgt_0_194,input [WEIGHT_SIZE-1:0] Wgt_0_195,input [WEIGHT_SIZE-1:0] Wgt_0_196,input [WEIGHT_SIZE-1:0] Wgt_0_197,input [WEIGHT_SIZE-1:0] Wgt_0_198,input [WEIGHT_SIZE-1:0] Wgt_0_199,input [WEIGHT_SIZE-1:0] Wgt_0_200,input [WEIGHT_SIZE-1:0] Wgt_0_201,input [WEIGHT_SIZE-1:0] Wgt_0_202,input [WEIGHT_SIZE-1:0] Wgt_0_203,input [WEIGHT_SIZE-1:0] Wgt_0_204,input [WEIGHT_SIZE-1:0] Wgt_0_205,input [WEIGHT_SIZE-1:0] Wgt_0_206,input [WEIGHT_SIZE-1:0] Wgt_0_207,input [WEIGHT_SIZE-1:0] Wgt_0_208,input [WEIGHT_SIZE-1:0] Wgt_0_209,input [WEIGHT_SIZE-1:0] Wgt_0_210,input [WEIGHT_SIZE-1:0] Wgt_0_211,input [WEIGHT_SIZE-1:0] Wgt_0_212,input [WEIGHT_SIZE-1:0] Wgt_0_213,input [WEIGHT_SIZE-1:0] Wgt_0_214,input [WEIGHT_SIZE-1:0] Wgt_0_215,input [WEIGHT_SIZE-1:0] Wgt_0_216,input [WEIGHT_SIZE-1:0] Wgt_0_217,input [WEIGHT_SIZE-1:0] Wgt_0_218,input [WEIGHT_SIZE-1:0] Wgt_0_219,input [WEIGHT_SIZE-1:0] Wgt_0_220,input [WEIGHT_SIZE-1:0] Wgt_0_221,input [WEIGHT_SIZE-1:0] Wgt_0_222,input [WEIGHT_SIZE-1:0] Wgt_0_223,input [WEIGHT_SIZE-1:0] Wgt_0_224,input [WEIGHT_SIZE-1:0] Wgt_0_225,input [WEIGHT_SIZE-1:0] Wgt_0_226,input [WEIGHT_SIZE-1:0] Wgt_0_227,input [WEIGHT_SIZE-1:0] Wgt_0_228,input [WEIGHT_SIZE-1:0] Wgt_0_229,input [WEIGHT_SIZE-1:0] Wgt_0_230,input [WEIGHT_SIZE-1:0] Wgt_0_231,input [WEIGHT_SIZE-1:0] Wgt_0_232,input [WEIGHT_SIZE-1:0] Wgt_0_233,input [WEIGHT_SIZE-1:0] Wgt_0_234,input [WEIGHT_SIZE-1:0] Wgt_0_235,input [WEIGHT_SIZE-1:0] Wgt_0_236,input [WEIGHT_SIZE-1:0] Wgt_0_237,input [WEIGHT_SIZE-1:0] Wgt_0_238,input [WEIGHT_SIZE-1:0] Wgt_0_239,input [WEIGHT_SIZE-1:0] Wgt_0_240,input [WEIGHT_SIZE-1:0] Wgt_0_241,input [WEIGHT_SIZE-1:0] Wgt_0_242,input [WEIGHT_SIZE-1:0] Wgt_0_243,input [WEIGHT_SIZE-1:0] Wgt_0_244,input [WEIGHT_SIZE-1:0] Wgt_0_245,input [WEIGHT_SIZE-1:0] Wgt_0_246,input [WEIGHT_SIZE-1:0] Wgt_0_247,input [WEIGHT_SIZE-1:0] Wgt_0_248,input [WEIGHT_SIZE-1:0] Wgt_0_249,input [WEIGHT_SIZE-1:0] Wgt_0_250,input [WEIGHT_SIZE-1:0] Wgt_0_251,input [WEIGHT_SIZE-1:0] Wgt_0_252,input [WEIGHT_SIZE-1:0] Wgt_0_253,input [WEIGHT_SIZE-1:0] Wgt_0_254,input [WEIGHT_SIZE-1:0] Wgt_0_255,input [WEIGHT_SIZE-1:0] Wgt_0_256,input [WEIGHT_SIZE-1:0] Wgt_0_257,input [WEIGHT_SIZE-1:0] Wgt_0_258,input [WEIGHT_SIZE-1:0] Wgt_0_259,input [WEIGHT_SIZE-1:0] Wgt_0_260,input [WEIGHT_SIZE-1:0] Wgt_0_261,input [WEIGHT_SIZE-1:0] Wgt_0_262,input [WEIGHT_SIZE-1:0] Wgt_0_263,input [WEIGHT_SIZE-1:0] Wgt_0_264,input [WEIGHT_SIZE-1:0] Wgt_0_265,input [WEIGHT_SIZE-1:0] Wgt_0_266,input [WEIGHT_SIZE-1:0] Wgt_0_267,input [WEIGHT_SIZE-1:0] Wgt_0_268,input [WEIGHT_SIZE-1:0] Wgt_0_269,input [WEIGHT_SIZE-1:0] Wgt_0_270,input [WEIGHT_SIZE-1:0] Wgt_0_271,input [WEIGHT_SIZE-1:0] Wgt_0_272,input [WEIGHT_SIZE-1:0] Wgt_0_273,input [WEIGHT_SIZE-1:0] Wgt_0_274,input [WEIGHT_SIZE-1:0] Wgt_0_275,input [WEIGHT_SIZE-1:0] Wgt_0_276,input [WEIGHT_SIZE-1:0] Wgt_0_277,input [WEIGHT_SIZE-1:0] Wgt_0_278,input [WEIGHT_SIZE-1:0] Wgt_0_279,input [WEIGHT_SIZE-1:0] Wgt_0_280,input [WEIGHT_SIZE-1:0] Wgt_0_281,input [WEIGHT_SIZE-1:0] Wgt_0_282,input [WEIGHT_SIZE-1:0] Wgt_0_283,input [WEIGHT_SIZE-1:0] Wgt_0_284,input [WEIGHT_SIZE-1:0] Wgt_0_285,input [WEIGHT_SIZE-1:0] Wgt_0_286,input [WEIGHT_SIZE-1:0] Wgt_0_287,input [WEIGHT_SIZE-1:0] Wgt_0_288,input [WEIGHT_SIZE-1:0] Wgt_0_289,input [WEIGHT_SIZE-1:0] Wgt_0_290,input [WEIGHT_SIZE-1:0] Wgt_0_291,input [WEIGHT_SIZE-1:0] Wgt_0_292,input [WEIGHT_SIZE-1:0] Wgt_0_293,input [WEIGHT_SIZE-1:0] Wgt_0_294,input [WEIGHT_SIZE-1:0] Wgt_0_295,input [WEIGHT_SIZE-1:0] Wgt_0_296,input [WEIGHT_SIZE-1:0] Wgt_0_297,input [WEIGHT_SIZE-1:0] Wgt_0_298,input [WEIGHT_SIZE-1:0] Wgt_0_299,input [WEIGHT_SIZE-1:0] Wgt_0_300,input [WEIGHT_SIZE-1:0] Wgt_0_301,input [WEIGHT_SIZE-1:0] Wgt_0_302,input [WEIGHT_SIZE-1:0] Wgt_0_303,input [WEIGHT_SIZE-1:0] Wgt_0_304,input [WEIGHT_SIZE-1:0] Wgt_0_305,input [WEIGHT_SIZE-1:0] Wgt_0_306,input [WEIGHT_SIZE-1:0] Wgt_0_307,input [WEIGHT_SIZE-1:0] Wgt_0_308,input [WEIGHT_SIZE-1:0] Wgt_0_309,input [WEIGHT_SIZE-1:0] Wgt_0_310,input [WEIGHT_SIZE-1:0] Wgt_0_311,input [WEIGHT_SIZE-1:0] Wgt_0_312,input [WEIGHT_SIZE-1:0] Wgt_0_313,input [WEIGHT_SIZE-1:0] Wgt_0_314,input [WEIGHT_SIZE-1:0] Wgt_0_315,input [WEIGHT_SIZE-1:0] Wgt_0_316,input [WEIGHT_SIZE-1:0] Wgt_0_317,input [WEIGHT_SIZE-1:0] Wgt_0_318,input [WEIGHT_SIZE-1:0] Wgt_0_319,input [WEIGHT_SIZE-1:0] Wgt_0_320,input [WEIGHT_SIZE-1:0] Wgt_0_321,input [WEIGHT_SIZE-1:0] Wgt_0_322,input [WEIGHT_SIZE-1:0] Wgt_0_323,input [WEIGHT_SIZE-1:0] Wgt_0_324,input [WEIGHT_SIZE-1:0] Wgt_0_325,input [WEIGHT_SIZE-1:0] Wgt_0_326,input [WEIGHT_SIZE-1:0] Wgt_0_327,input [WEIGHT_SIZE-1:0] Wgt_0_328,input [WEIGHT_SIZE-1:0] Wgt_0_329,input [WEIGHT_SIZE-1:0] Wgt_0_330,input [WEIGHT_SIZE-1:0] Wgt_0_331,input [WEIGHT_SIZE-1:0] Wgt_0_332,input [WEIGHT_SIZE-1:0] Wgt_0_333,input [WEIGHT_SIZE-1:0] Wgt_0_334,input [WEIGHT_SIZE-1:0] Wgt_0_335,input [WEIGHT_SIZE-1:0] Wgt_0_336,input [WEIGHT_SIZE-1:0] Wgt_0_337,input [WEIGHT_SIZE-1:0] Wgt_0_338,input [WEIGHT_SIZE-1:0] Wgt_0_339,input [WEIGHT_SIZE-1:0] Wgt_0_340,input [WEIGHT_SIZE-1:0] Wgt_0_341,input [WEIGHT_SIZE-1:0] Wgt_0_342,input [WEIGHT_SIZE-1:0] Wgt_0_343,input [WEIGHT_SIZE-1:0] Wgt_0_344,input [WEIGHT_SIZE-1:0] Wgt_0_345,input [WEIGHT_SIZE-1:0] Wgt_0_346,input [WEIGHT_SIZE-1:0] Wgt_0_347,input [WEIGHT_SIZE-1:0] Wgt_0_348,input [WEIGHT_SIZE-1:0] Wgt_0_349,input [WEIGHT_SIZE-1:0] Wgt_0_350,input [WEIGHT_SIZE-1:0] Wgt_0_351,input [WEIGHT_SIZE-1:0] Wgt_0_352,input [WEIGHT_SIZE-1:0] Wgt_0_353,input [WEIGHT_SIZE-1:0] Wgt_0_354,input [WEIGHT_SIZE-1:0] Wgt_0_355,input [WEIGHT_SIZE-1:0] Wgt_0_356,input [WEIGHT_SIZE-1:0] Wgt_0_357,input [WEIGHT_SIZE-1:0] Wgt_0_358,input [WEIGHT_SIZE-1:0] Wgt_0_359,input [WEIGHT_SIZE-1:0] Wgt_0_360,input [WEIGHT_SIZE-1:0] Wgt_0_361,input [WEIGHT_SIZE-1:0] Wgt_0_362,input [WEIGHT_SIZE-1:0] Wgt_0_363,input [WEIGHT_SIZE-1:0] Wgt_0_364,input [WEIGHT_SIZE-1:0] Wgt_0_365,input [WEIGHT_SIZE-1:0] Wgt_0_366,input [WEIGHT_SIZE-1:0] Wgt_0_367,input [WEIGHT_SIZE-1:0] Wgt_0_368,input [WEIGHT_SIZE-1:0] Wgt_0_369,input [WEIGHT_SIZE-1:0] Wgt_0_370,input [WEIGHT_SIZE-1:0] Wgt_0_371,input [WEIGHT_SIZE-1:0] Wgt_0_372,input [WEIGHT_SIZE-1:0] Wgt_0_373,input [WEIGHT_SIZE-1:0] Wgt_0_374,input [WEIGHT_SIZE-1:0] Wgt_0_375,input [WEIGHT_SIZE-1:0] Wgt_0_376,input [WEIGHT_SIZE-1:0] Wgt_0_377,input [WEIGHT_SIZE-1:0] Wgt_0_378,input [WEIGHT_SIZE-1:0] Wgt_0_379,input [WEIGHT_SIZE-1:0] Wgt_0_380,input [WEIGHT_SIZE-1:0] Wgt_0_381,input [WEIGHT_SIZE-1:0] Wgt_0_382,input [WEIGHT_SIZE-1:0] Wgt_0_383,input [WEIGHT_SIZE-1:0] Wgt_0_384,input [WEIGHT_SIZE-1:0] Wgt_0_385,input [WEIGHT_SIZE-1:0] Wgt_0_386,input [WEIGHT_SIZE-1:0] Wgt_0_387,input [WEIGHT_SIZE-1:0] Wgt_0_388,input [WEIGHT_SIZE-1:0] Wgt_0_389,input [WEIGHT_SIZE-1:0] Wgt_0_390,input [WEIGHT_SIZE-1:0] Wgt_0_391,input [WEIGHT_SIZE-1:0] Wgt_0_392,input [WEIGHT_SIZE-1:0] Wgt_0_393,input [WEIGHT_SIZE-1:0] Wgt_0_394,input [WEIGHT_SIZE-1:0] Wgt_0_395,input [WEIGHT_SIZE-1:0] Wgt_0_396,input [WEIGHT_SIZE-1:0] Wgt_0_397,input [WEIGHT_SIZE-1:0] Wgt_0_398,input [WEIGHT_SIZE-1:0] Wgt_0_399,input [WEIGHT_SIZE-1:0] Wgt_0_400,input [WEIGHT_SIZE-1:0] Wgt_0_401,input [WEIGHT_SIZE-1:0] Wgt_0_402,input [WEIGHT_SIZE-1:0] Wgt_0_403,input [WEIGHT_SIZE-1:0] Wgt_0_404,input [WEIGHT_SIZE-1:0] Wgt_0_405,input [WEIGHT_SIZE-1:0] Wgt_0_406,input [WEIGHT_SIZE-1:0] Wgt_0_407,input [WEIGHT_SIZE-1:0] Wgt_0_408,input [WEIGHT_SIZE-1:0] Wgt_0_409,input [WEIGHT_SIZE-1:0] Wgt_0_410,input [WEIGHT_SIZE-1:0] Wgt_0_411,input [WEIGHT_SIZE-1:0] Wgt_0_412,input [WEIGHT_SIZE-1:0] Wgt_0_413,input [WEIGHT_SIZE-1:0] Wgt_0_414,input [WEIGHT_SIZE-1:0] Wgt_0_415,input [WEIGHT_SIZE-1:0] Wgt_0_416,input [WEIGHT_SIZE-1:0] Wgt_0_417,input [WEIGHT_SIZE-1:0] Wgt_0_418,input [WEIGHT_SIZE-1:0] Wgt_0_419,input [WEIGHT_SIZE-1:0] Wgt_0_420,input [WEIGHT_SIZE-1:0] Wgt_0_421,input [WEIGHT_SIZE-1:0] Wgt_0_422,input [WEIGHT_SIZE-1:0] Wgt_0_423,input [WEIGHT_SIZE-1:0] Wgt_0_424,input [WEIGHT_SIZE-1:0] Wgt_0_425,input [WEIGHT_SIZE-1:0] Wgt_0_426,input [WEIGHT_SIZE-1:0] Wgt_0_427,input [WEIGHT_SIZE-1:0] Wgt_0_428,input [WEIGHT_SIZE-1:0] Wgt_0_429,input [WEIGHT_SIZE-1:0] Wgt_0_430,input [WEIGHT_SIZE-1:0] Wgt_0_431,input [WEIGHT_SIZE-1:0] Wgt_0_432,input [WEIGHT_SIZE-1:0] Wgt_0_433,input [WEIGHT_SIZE-1:0] Wgt_0_434,input [WEIGHT_SIZE-1:0] Wgt_0_435,input [WEIGHT_SIZE-1:0] Wgt_0_436,input [WEIGHT_SIZE-1:0] Wgt_0_437,input [WEIGHT_SIZE-1:0] Wgt_0_438,input [WEIGHT_SIZE-1:0] Wgt_0_439,input [WEIGHT_SIZE-1:0] Wgt_0_440,input [WEIGHT_SIZE-1:0] Wgt_0_441,input [WEIGHT_SIZE-1:0] Wgt_0_442,input [WEIGHT_SIZE-1:0] Wgt_0_443,input [WEIGHT_SIZE-1:0] Wgt_0_444,input [WEIGHT_SIZE-1:0] Wgt_0_445,input [WEIGHT_SIZE-1:0] Wgt_0_446,input [WEIGHT_SIZE-1:0] Wgt_0_447,input [WEIGHT_SIZE-1:0] Wgt_0_448,input [WEIGHT_SIZE-1:0] Wgt_0_449,input [WEIGHT_SIZE-1:0] Wgt_0_450,input [WEIGHT_SIZE-1:0] Wgt_0_451,input [WEIGHT_SIZE-1:0] Wgt_0_452,input [WEIGHT_SIZE-1:0] Wgt_0_453,input [WEIGHT_SIZE-1:0] Wgt_0_454,input [WEIGHT_SIZE-1:0] Wgt_0_455,input [WEIGHT_SIZE-1:0] Wgt_0_456,input [WEIGHT_SIZE-1:0] Wgt_0_457,input [WEIGHT_SIZE-1:0] Wgt_0_458,input [WEIGHT_SIZE-1:0] Wgt_0_459,input [WEIGHT_SIZE-1:0] Wgt_0_460,input [WEIGHT_SIZE-1:0] Wgt_0_461,input [WEIGHT_SIZE-1:0] Wgt_0_462,input [WEIGHT_SIZE-1:0] Wgt_0_463,input [WEIGHT_SIZE-1:0] Wgt_0_464,input [WEIGHT_SIZE-1:0] Wgt_0_465,input [WEIGHT_SIZE-1:0] Wgt_0_466,input [WEIGHT_SIZE-1:0] Wgt_0_467,input [WEIGHT_SIZE-1:0] Wgt_0_468,input [WEIGHT_SIZE-1:0] Wgt_0_469,input [WEIGHT_SIZE-1:0] Wgt_0_470,input [WEIGHT_SIZE-1:0] Wgt_0_471,input [WEIGHT_SIZE-1:0] Wgt_0_472,input [WEIGHT_SIZE-1:0] Wgt_0_473,input [WEIGHT_SIZE-1:0] Wgt_0_474,input [WEIGHT_SIZE-1:0] Wgt_0_475,input [WEIGHT_SIZE-1:0] Wgt_0_476,input [WEIGHT_SIZE-1:0] Wgt_0_477,input [WEIGHT_SIZE-1:0] Wgt_0_478,input [WEIGHT_SIZE-1:0] Wgt_0_479,input [WEIGHT_SIZE-1:0] Wgt_0_480,input [WEIGHT_SIZE-1:0] Wgt_0_481,input [WEIGHT_SIZE-1:0] Wgt_0_482,input [WEIGHT_SIZE-1:0] Wgt_0_483,input [WEIGHT_SIZE-1:0] Wgt_0_484,input [WEIGHT_SIZE-1:0] Wgt_0_485,input [WEIGHT_SIZE-1:0] Wgt_0_486,input [WEIGHT_SIZE-1:0] Wgt_0_487,input [WEIGHT_SIZE-1:0] Wgt_0_488,input [WEIGHT_SIZE-1:0] Wgt_0_489,input [WEIGHT_SIZE-1:0] Wgt_0_490,input [WEIGHT_SIZE-1:0] Wgt_0_491,input [WEIGHT_SIZE-1:0] Wgt_0_492,input [WEIGHT_SIZE-1:0] Wgt_0_493,input [WEIGHT_SIZE-1:0] Wgt_0_494,input [WEIGHT_SIZE-1:0] Wgt_0_495,input [WEIGHT_SIZE-1:0] Wgt_0_496,input [WEIGHT_SIZE-1:0] Wgt_0_497,input [WEIGHT_SIZE-1:0] Wgt_0_498,input [WEIGHT_SIZE-1:0] Wgt_0_499,input [WEIGHT_SIZE-1:0] Wgt_0_500,input [WEIGHT_SIZE-1:0] Wgt_0_501,input [WEIGHT_SIZE-1:0] Wgt_0_502,input [WEIGHT_SIZE-1:0] Wgt_0_503,input [WEIGHT_SIZE-1:0] Wgt_0_504,input [WEIGHT_SIZE-1:0] Wgt_0_505,input [WEIGHT_SIZE-1:0] Wgt_0_506,input [WEIGHT_SIZE-1:0] Wgt_0_507,input [WEIGHT_SIZE-1:0] Wgt_0_508,input [WEIGHT_SIZE-1:0] Wgt_0_509,input [WEIGHT_SIZE-1:0] Wgt_0_510,input [WEIGHT_SIZE-1:0] Wgt_0_511,input [WEIGHT_SIZE-1:0] Wgt_0_512,input [WEIGHT_SIZE-1:0] Wgt_0_513,input [WEIGHT_SIZE-1:0] Wgt_0_514,input [WEIGHT_SIZE-1:0] Wgt_0_515,input [WEIGHT_SIZE-1:0] Wgt_0_516,input [WEIGHT_SIZE-1:0] Wgt_0_517,input [WEIGHT_SIZE-1:0] Wgt_0_518,input [WEIGHT_SIZE-1:0] Wgt_0_519,input [WEIGHT_SIZE-1:0] Wgt_0_520,input [WEIGHT_SIZE-1:0] Wgt_0_521,input [WEIGHT_SIZE-1:0] Wgt_0_522,input [WEIGHT_SIZE-1:0] Wgt_0_523,input [WEIGHT_SIZE-1:0] Wgt_0_524,input [WEIGHT_SIZE-1:0] Wgt_0_525,input [WEIGHT_SIZE-1:0] Wgt_0_526,input [WEIGHT_SIZE-1:0] Wgt_0_527,input [WEIGHT_SIZE-1:0] Wgt_0_528,input [WEIGHT_SIZE-1:0] Wgt_0_529,input [WEIGHT_SIZE-1:0] Wgt_0_530,input [WEIGHT_SIZE-1:0] Wgt_0_531,input [WEIGHT_SIZE-1:0] Wgt_0_532,input [WEIGHT_SIZE-1:0] Wgt_0_533,input [WEIGHT_SIZE-1:0] Wgt_0_534,input [WEIGHT_SIZE-1:0] Wgt_0_535,input [WEIGHT_SIZE-1:0] Wgt_0_536,input [WEIGHT_SIZE-1:0] Wgt_0_537,input [WEIGHT_SIZE-1:0] Wgt_0_538,input [WEIGHT_SIZE-1:0] Wgt_0_539,input [WEIGHT_SIZE-1:0] Wgt_0_540,input [WEIGHT_SIZE-1:0] Wgt_0_541,input [WEIGHT_SIZE-1:0] Wgt_0_542,input [WEIGHT_SIZE-1:0] Wgt_0_543,input [WEIGHT_SIZE-1:0] Wgt_0_544,input [WEIGHT_SIZE-1:0] Wgt_0_545,input [WEIGHT_SIZE-1:0] Wgt_0_546,input [WEIGHT_SIZE-1:0] Wgt_0_547,input [WEIGHT_SIZE-1:0] Wgt_0_548,input [WEIGHT_SIZE-1:0] Wgt_0_549,input [WEIGHT_SIZE-1:0] Wgt_0_550,input [WEIGHT_SIZE-1:0] Wgt_0_551,input [WEIGHT_SIZE-1:0] Wgt_0_552,input [WEIGHT_SIZE-1:0] Wgt_0_553,input [WEIGHT_SIZE-1:0] Wgt_0_554,input [WEIGHT_SIZE-1:0] Wgt_0_555,input [WEIGHT_SIZE-1:0] Wgt_0_556,input [WEIGHT_SIZE-1:0] Wgt_0_557,input [WEIGHT_SIZE-1:0] Wgt_0_558,input [WEIGHT_SIZE-1:0] Wgt_0_559,input [WEIGHT_SIZE-1:0] Wgt_0_560,input [WEIGHT_SIZE-1:0] Wgt_0_561,input [WEIGHT_SIZE-1:0] Wgt_0_562,input [WEIGHT_SIZE-1:0] Wgt_0_563,input [WEIGHT_SIZE-1:0] Wgt_0_564,input [WEIGHT_SIZE-1:0] Wgt_0_565,input [WEIGHT_SIZE-1:0] Wgt_0_566,input [WEIGHT_SIZE-1:0] Wgt_0_567,input [WEIGHT_SIZE-1:0] Wgt_0_568,input [WEIGHT_SIZE-1:0] Wgt_0_569,input [WEIGHT_SIZE-1:0] Wgt_0_570,input [WEIGHT_SIZE-1:0] Wgt_0_571,input [WEIGHT_SIZE-1:0] Wgt_0_572,input [WEIGHT_SIZE-1:0] Wgt_0_573,input [WEIGHT_SIZE-1:0] Wgt_0_574,input [WEIGHT_SIZE-1:0] Wgt_0_575,input [WEIGHT_SIZE-1:0] Wgt_0_576,input [WEIGHT_SIZE-1:0] Wgt_0_577,input [WEIGHT_SIZE-1:0] Wgt_0_578,input [WEIGHT_SIZE-1:0] Wgt_0_579,input [WEIGHT_SIZE-1:0] Wgt_0_580,input [WEIGHT_SIZE-1:0] Wgt_0_581,input [WEIGHT_SIZE-1:0] Wgt_0_582,input [WEIGHT_SIZE-1:0] Wgt_0_583,input [WEIGHT_SIZE-1:0] Wgt_0_584,input [WEIGHT_SIZE-1:0] Wgt_0_585,input [WEIGHT_SIZE-1:0] Wgt_0_586,input [WEIGHT_SIZE-1:0] Wgt_0_587,input [WEIGHT_SIZE-1:0] Wgt_0_588,input [WEIGHT_SIZE-1:0] Wgt_0_589,input [WEIGHT_SIZE-1:0] Wgt_0_590,input [WEIGHT_SIZE-1:0] Wgt_0_591,input [WEIGHT_SIZE-1:0] Wgt_0_592,input [WEIGHT_SIZE-1:0] Wgt_0_593,input [WEIGHT_SIZE-1:0] Wgt_0_594,input [WEIGHT_SIZE-1:0] Wgt_0_595,input [WEIGHT_SIZE-1:0] Wgt_0_596,input [WEIGHT_SIZE-1:0] Wgt_0_597,input [WEIGHT_SIZE-1:0] Wgt_0_598,input [WEIGHT_SIZE-1:0] Wgt_0_599,input [WEIGHT_SIZE-1:0] Wgt_0_600,input [WEIGHT_SIZE-1:0] Wgt_0_601,input [WEIGHT_SIZE-1:0] Wgt_0_602,input [WEIGHT_SIZE-1:0] Wgt_0_603,input [WEIGHT_SIZE-1:0] Wgt_0_604,input [WEIGHT_SIZE-1:0] Wgt_0_605,input [WEIGHT_SIZE-1:0] Wgt_0_606,input [WEIGHT_SIZE-1:0] Wgt_0_607,input [WEIGHT_SIZE-1:0] Wgt_0_608,input [WEIGHT_SIZE-1:0] Wgt_0_609,input [WEIGHT_SIZE-1:0] Wgt_0_610,input [WEIGHT_SIZE-1:0] Wgt_0_611,input [WEIGHT_SIZE-1:0] Wgt_0_612,input [WEIGHT_SIZE-1:0] Wgt_0_613,input [WEIGHT_SIZE-1:0] Wgt_0_614,input [WEIGHT_SIZE-1:0] Wgt_0_615,input [WEIGHT_SIZE-1:0] Wgt_0_616,input [WEIGHT_SIZE-1:0] Wgt_0_617,input [WEIGHT_SIZE-1:0] Wgt_0_618,input [WEIGHT_SIZE-1:0] Wgt_0_619,input [WEIGHT_SIZE-1:0] Wgt_0_620,input [WEIGHT_SIZE-1:0] Wgt_0_621,input [WEIGHT_SIZE-1:0] Wgt_0_622,input [WEIGHT_SIZE-1:0] Wgt_0_623,input [WEIGHT_SIZE-1:0] Wgt_0_624,input [WEIGHT_SIZE-1:0] Wgt_0_625,input [WEIGHT_SIZE-1:0] Wgt_0_626,input [WEIGHT_SIZE-1:0] Wgt_0_627,input [WEIGHT_SIZE-1:0] Wgt_0_628,input [WEIGHT_SIZE-1:0] Wgt_0_629,input [WEIGHT_SIZE-1:0] Wgt_0_630,input [WEIGHT_SIZE-1:0] Wgt_0_631,input [WEIGHT_SIZE-1:0] Wgt_0_632,input [WEIGHT_SIZE-1:0] Wgt_0_633,input [WEIGHT_SIZE-1:0] Wgt_0_634,input [WEIGHT_SIZE-1:0] Wgt_0_635,input [WEIGHT_SIZE-1:0] Wgt_0_636,input [WEIGHT_SIZE-1:0] Wgt_0_637,input [WEIGHT_SIZE-1:0] Wgt_0_638,input [WEIGHT_SIZE-1:0] Wgt_0_639,input [WEIGHT_SIZE-1:0] Wgt_0_640,input [WEIGHT_SIZE-1:0] Wgt_0_641,input [WEIGHT_SIZE-1:0] Wgt_0_642,input [WEIGHT_SIZE-1:0] Wgt_0_643,input [WEIGHT_SIZE-1:0] Wgt_0_644,input [WEIGHT_SIZE-1:0] Wgt_0_645,input [WEIGHT_SIZE-1:0] Wgt_0_646,input [WEIGHT_SIZE-1:0] Wgt_0_647,input [WEIGHT_SIZE-1:0] Wgt_0_648,input [WEIGHT_SIZE-1:0] Wgt_0_649,input [WEIGHT_SIZE-1:0] Wgt_0_650,input [WEIGHT_SIZE-1:0] Wgt_0_651,input [WEIGHT_SIZE-1:0] Wgt_0_652,input [WEIGHT_SIZE-1:0] Wgt_0_653,input [WEIGHT_SIZE-1:0] Wgt_0_654,input [WEIGHT_SIZE-1:0] Wgt_0_655,input [WEIGHT_SIZE-1:0] Wgt_0_656,input [WEIGHT_SIZE-1:0] Wgt_0_657,input [WEIGHT_SIZE-1:0] Wgt_0_658,input [WEIGHT_SIZE-1:0] Wgt_0_659,input [WEIGHT_SIZE-1:0] Wgt_0_660,input [WEIGHT_SIZE-1:0] Wgt_0_661,input [WEIGHT_SIZE-1:0] Wgt_0_662,input [WEIGHT_SIZE-1:0] Wgt_0_663,input [WEIGHT_SIZE-1:0] Wgt_0_664,input [WEIGHT_SIZE-1:0] Wgt_0_665,input [WEIGHT_SIZE-1:0] Wgt_0_666,input [WEIGHT_SIZE-1:0] Wgt_0_667,input [WEIGHT_SIZE-1:0] Wgt_0_668,input [WEIGHT_SIZE-1:0] Wgt_0_669,input [WEIGHT_SIZE-1:0] Wgt_0_670,input [WEIGHT_SIZE-1:0] Wgt_0_671,input [WEIGHT_SIZE-1:0] Wgt_0_672,input [WEIGHT_SIZE-1:0] Wgt_0_673,input [WEIGHT_SIZE-1:0] Wgt_0_674,input [WEIGHT_SIZE-1:0] Wgt_0_675,input [WEIGHT_SIZE-1:0] Wgt_0_676,input [WEIGHT_SIZE-1:0] Wgt_0_677,input [WEIGHT_SIZE-1:0] Wgt_0_678,input [WEIGHT_SIZE-1:0] Wgt_0_679,input [WEIGHT_SIZE-1:0] Wgt_0_680,input [WEIGHT_SIZE-1:0] Wgt_0_681,input [WEIGHT_SIZE-1:0] Wgt_0_682,input [WEIGHT_SIZE-1:0] Wgt_0_683,input [WEIGHT_SIZE-1:0] Wgt_0_684,input [WEIGHT_SIZE-1:0] Wgt_0_685,input [WEIGHT_SIZE-1:0] Wgt_0_686,input [WEIGHT_SIZE-1:0] Wgt_0_687,input [WEIGHT_SIZE-1:0] Wgt_0_688,input [WEIGHT_SIZE-1:0] Wgt_0_689,input [WEIGHT_SIZE-1:0] Wgt_0_690,input [WEIGHT_SIZE-1:0] Wgt_0_691,input [WEIGHT_SIZE-1:0] Wgt_0_692,input [WEIGHT_SIZE-1:0] Wgt_0_693,input [WEIGHT_SIZE-1:0] Wgt_0_694,input [WEIGHT_SIZE-1:0] Wgt_0_695,input [WEIGHT_SIZE-1:0] Wgt_0_696,input [WEIGHT_SIZE-1:0] Wgt_0_697,input [WEIGHT_SIZE-1:0] Wgt_0_698,input [WEIGHT_SIZE-1:0] Wgt_0_699,input [WEIGHT_SIZE-1:0] Wgt_0_700,input [WEIGHT_SIZE-1:0] Wgt_0_701,input [WEIGHT_SIZE-1:0] Wgt_0_702,input [WEIGHT_SIZE-1:0] Wgt_0_703,input [WEIGHT_SIZE-1:0] Wgt_0_704,input [WEIGHT_SIZE-1:0] Wgt_0_705,input [WEIGHT_SIZE-1:0] Wgt_0_706,input [WEIGHT_SIZE-1:0] Wgt_0_707,input [WEIGHT_SIZE-1:0] Wgt_0_708,input [WEIGHT_SIZE-1:0] Wgt_0_709,input [WEIGHT_SIZE-1:0] Wgt_0_710,input [WEIGHT_SIZE-1:0] Wgt_0_711,input [WEIGHT_SIZE-1:0] Wgt_0_712,input [WEIGHT_SIZE-1:0] Wgt_0_713,input [WEIGHT_SIZE-1:0] Wgt_0_714,input [WEIGHT_SIZE-1:0] Wgt_0_715,input [WEIGHT_SIZE-1:0] Wgt_0_716,input [WEIGHT_SIZE-1:0] Wgt_0_717,input [WEIGHT_SIZE-1:0] Wgt_0_718,input [WEIGHT_SIZE-1:0] Wgt_0_719,input [WEIGHT_SIZE-1:0] Wgt_0_720,input [WEIGHT_SIZE-1:0] Wgt_0_721,input [WEIGHT_SIZE-1:0] Wgt_0_722,input [WEIGHT_SIZE-1:0] Wgt_0_723,input [WEIGHT_SIZE-1:0] Wgt_0_724,input [WEIGHT_SIZE-1:0] Wgt_0_725,input [WEIGHT_SIZE-1:0] Wgt_0_726,input [WEIGHT_SIZE-1:0] Wgt_0_727,input [WEIGHT_SIZE-1:0] Wgt_0_728,input [WEIGHT_SIZE-1:0] Wgt_0_729,input [WEIGHT_SIZE-1:0] Wgt_0_730,input [WEIGHT_SIZE-1:0] Wgt_0_731,input [WEIGHT_SIZE-1:0] Wgt_0_732,input [WEIGHT_SIZE-1:0] Wgt_0_733,input [WEIGHT_SIZE-1:0] Wgt_0_734,input [WEIGHT_SIZE-1:0] Wgt_0_735,input [WEIGHT_SIZE-1:0] Wgt_0_736,input [WEIGHT_SIZE-1:0] Wgt_0_737,input [WEIGHT_SIZE-1:0] Wgt_0_738,input [WEIGHT_SIZE-1:0] Wgt_0_739,input [WEIGHT_SIZE-1:0] Wgt_0_740,input [WEIGHT_SIZE-1:0] Wgt_0_741,input [WEIGHT_SIZE-1:0] Wgt_0_742,input [WEIGHT_SIZE-1:0] Wgt_0_743,input [WEIGHT_SIZE-1:0] Wgt_0_744,input [WEIGHT_SIZE-1:0] Wgt_0_745,input [WEIGHT_SIZE-1:0] Wgt_0_746,input [WEIGHT_SIZE-1:0] Wgt_0_747,input [WEIGHT_SIZE-1:0] Wgt_0_748,input [WEIGHT_SIZE-1:0] Wgt_0_749,input [WEIGHT_SIZE-1:0] Wgt_0_750,input [WEIGHT_SIZE-1:0] Wgt_0_751,input [WEIGHT_SIZE-1:0] Wgt_0_752,input [WEIGHT_SIZE-1:0] Wgt_0_753,input [WEIGHT_SIZE-1:0] Wgt_0_754,input [WEIGHT_SIZE-1:0] Wgt_0_755,input [WEIGHT_SIZE-1:0] Wgt_0_756,input [WEIGHT_SIZE-1:0] Wgt_0_757,input [WEIGHT_SIZE-1:0] Wgt_0_758,input [WEIGHT_SIZE-1:0] Wgt_0_759,input [WEIGHT_SIZE-1:0] Wgt_0_760,input [WEIGHT_SIZE-1:0] Wgt_0_761,input [WEIGHT_SIZE-1:0] Wgt_0_762,input [WEIGHT_SIZE-1:0] Wgt_0_763,input [WEIGHT_SIZE-1:0] Wgt_0_764,input [WEIGHT_SIZE-1:0] Wgt_0_765,input [WEIGHT_SIZE-1:0] Wgt_0_766,input [WEIGHT_SIZE-1:0] Wgt_0_767,input [WEIGHT_SIZE-1:0] Wgt_0_768,input [WEIGHT_SIZE-1:0] Wgt_0_769,input [WEIGHT_SIZE-1:0] Wgt_0_770,input [WEIGHT_SIZE-1:0] Wgt_0_771,input [WEIGHT_SIZE-1:0] Wgt_0_772,input [WEIGHT_SIZE-1:0] Wgt_0_773,input [WEIGHT_SIZE-1:0] Wgt_0_774,input [WEIGHT_SIZE-1:0] Wgt_0_775,input [WEIGHT_SIZE-1:0] Wgt_0_776,input [WEIGHT_SIZE-1:0] Wgt_0_777,input [WEIGHT_SIZE-1:0] Wgt_0_778,input [WEIGHT_SIZE-1:0] Wgt_0_779,input [WEIGHT_SIZE-1:0] Wgt_0_780,input [WEIGHT_SIZE-1:0] Wgt_0_781,input [WEIGHT_SIZE-1:0] Wgt_0_782,input [WEIGHT_SIZE-1:0] Wgt_0_783,input [WEIGHT_SIZE-1:0] Wgt_0_784,input [WEIGHT_SIZE-1:0] Wgt_1_0,input [WEIGHT_SIZE-1:0] Wgt_1_1,input [WEIGHT_SIZE-1:0] Wgt_1_2,input [WEIGHT_SIZE-1:0] Wgt_1_3,input [WEIGHT_SIZE-1:0] Wgt_1_4,input [WEIGHT_SIZE-1:0] Wgt_1_5,input [WEIGHT_SIZE-1:0] Wgt_1_6,input [WEIGHT_SIZE-1:0] Wgt_1_7,input [WEIGHT_SIZE-1:0] Wgt_1_8,input [WEIGHT_SIZE-1:0] Wgt_1_9,input [WEIGHT_SIZE-1:0] Wgt_1_10,input [WEIGHT_SIZE-1:0] Wgt_1_11,input [WEIGHT_SIZE-1:0] Wgt_1_12,input [WEIGHT_SIZE-1:0] Wgt_1_13,input [WEIGHT_SIZE-1:0] Wgt_1_14,input [WEIGHT_SIZE-1:0] Wgt_1_15,input [WEIGHT_SIZE-1:0] Wgt_1_16,input [WEIGHT_SIZE-1:0] Wgt_1_17,input [WEIGHT_SIZE-1:0] Wgt_1_18,input [WEIGHT_SIZE-1:0] Wgt_1_19,input [WEIGHT_SIZE-1:0] Wgt_1_20,input [WEIGHT_SIZE-1:0] Wgt_1_21,input [WEIGHT_SIZE-1:0] Wgt_1_22,input [WEIGHT_SIZE-1:0] Wgt_1_23,input [WEIGHT_SIZE-1:0] Wgt_1_24,input [WEIGHT_SIZE-1:0] Wgt_1_25,input [WEIGHT_SIZE-1:0] Wgt_1_26,input [WEIGHT_SIZE-1:0] Wgt_1_27,input [WEIGHT_SIZE-1:0] Wgt_1_28,input [WEIGHT_SIZE-1:0] Wgt_1_29,input [WEIGHT_SIZE-1:0] Wgt_1_30,input [WEIGHT_SIZE-1:0] Wgt_1_31,input [WEIGHT_SIZE-1:0] Wgt_1_32,input [WEIGHT_SIZE-1:0] Wgt_1_33,input [WEIGHT_SIZE-1:0] Wgt_1_34,input [WEIGHT_SIZE-1:0] Wgt_1_35,input [WEIGHT_SIZE-1:0] Wgt_1_36,input [WEIGHT_SIZE-1:0] Wgt_1_37,input [WEIGHT_SIZE-1:0] Wgt_1_38,input [WEIGHT_SIZE-1:0] Wgt_1_39,input [WEIGHT_SIZE-1:0] Wgt_1_40,input [WEIGHT_SIZE-1:0] Wgt_1_41,input [WEIGHT_SIZE-1:0] Wgt_1_42,input [WEIGHT_SIZE-1:0] Wgt_1_43,input [WEIGHT_SIZE-1:0] Wgt_1_44,input [WEIGHT_SIZE-1:0] Wgt_1_45,input [WEIGHT_SIZE-1:0] Wgt_1_46,input [WEIGHT_SIZE-1:0] Wgt_1_47,input [WEIGHT_SIZE-1:0] Wgt_1_48,input [WEIGHT_SIZE-1:0] Wgt_1_49,input [WEIGHT_SIZE-1:0] Wgt_1_50,input [WEIGHT_SIZE-1:0] Wgt_1_51,input [WEIGHT_SIZE-1:0] Wgt_1_52,input [WEIGHT_SIZE-1:0] Wgt_1_53,input [WEIGHT_SIZE-1:0] Wgt_1_54,input [WEIGHT_SIZE-1:0] Wgt_1_55,input [WEIGHT_SIZE-1:0] Wgt_1_56,input [WEIGHT_SIZE-1:0] Wgt_1_57,input [WEIGHT_SIZE-1:0] Wgt_1_58,input [WEIGHT_SIZE-1:0] Wgt_1_59,input [WEIGHT_SIZE-1:0] Wgt_1_60,input [WEIGHT_SIZE-1:0] Wgt_1_61,input [WEIGHT_SIZE-1:0] Wgt_1_62,input [WEIGHT_SIZE-1:0] Wgt_1_63,input [WEIGHT_SIZE-1:0] Wgt_1_64,input [WEIGHT_SIZE-1:0] Wgt_1_65,input [WEIGHT_SIZE-1:0] Wgt_1_66,input [WEIGHT_SIZE-1:0] Wgt_1_67,input [WEIGHT_SIZE-1:0] Wgt_1_68,input [WEIGHT_SIZE-1:0] Wgt_1_69,input [WEIGHT_SIZE-1:0] Wgt_1_70,input [WEIGHT_SIZE-1:0] Wgt_1_71,input [WEIGHT_SIZE-1:0] Wgt_1_72,input [WEIGHT_SIZE-1:0] Wgt_1_73,input [WEIGHT_SIZE-1:0] Wgt_1_74,input [WEIGHT_SIZE-1:0] Wgt_1_75,input [WEIGHT_SIZE-1:0] Wgt_1_76,input [WEIGHT_SIZE-1:0] Wgt_1_77,input [WEIGHT_SIZE-1:0] Wgt_1_78,input [WEIGHT_SIZE-1:0] Wgt_1_79,input [WEIGHT_SIZE-1:0] Wgt_1_80,input [WEIGHT_SIZE-1:0] Wgt_1_81,input [WEIGHT_SIZE-1:0] Wgt_1_82,input [WEIGHT_SIZE-1:0] Wgt_1_83,input [WEIGHT_SIZE-1:0] Wgt_1_84,input [WEIGHT_SIZE-1:0] Wgt_1_85,input [WEIGHT_SIZE-1:0] Wgt_1_86,input [WEIGHT_SIZE-1:0] Wgt_1_87,input [WEIGHT_SIZE-1:0] Wgt_1_88,input [WEIGHT_SIZE-1:0] Wgt_1_89,input [WEIGHT_SIZE-1:0] Wgt_1_90,input [WEIGHT_SIZE-1:0] Wgt_1_91,input [WEIGHT_SIZE-1:0] Wgt_1_92,input [WEIGHT_SIZE-1:0] Wgt_1_93,input [WEIGHT_SIZE-1:0] Wgt_1_94,input [WEIGHT_SIZE-1:0] Wgt_1_95,input [WEIGHT_SIZE-1:0] Wgt_1_96,input [WEIGHT_SIZE-1:0] Wgt_1_97,input [WEIGHT_SIZE-1:0] Wgt_1_98,input [WEIGHT_SIZE-1:0] Wgt_1_99,input [WEIGHT_SIZE-1:0] Wgt_1_100,input [WEIGHT_SIZE-1:0] Wgt_1_101,input [WEIGHT_SIZE-1:0] Wgt_1_102,input [WEIGHT_SIZE-1:0] Wgt_1_103,input [WEIGHT_SIZE-1:0] Wgt_1_104,input [WEIGHT_SIZE-1:0] Wgt_1_105,input [WEIGHT_SIZE-1:0] Wgt_1_106,input [WEIGHT_SIZE-1:0] Wgt_1_107,input [WEIGHT_SIZE-1:0] Wgt_1_108,input [WEIGHT_SIZE-1:0] Wgt_1_109,input [WEIGHT_SIZE-1:0] Wgt_1_110,input [WEIGHT_SIZE-1:0] Wgt_1_111,input [WEIGHT_SIZE-1:0] Wgt_1_112,input [WEIGHT_SIZE-1:0] Wgt_1_113,input [WEIGHT_SIZE-1:0] Wgt_1_114,input [WEIGHT_SIZE-1:0] Wgt_1_115,input [WEIGHT_SIZE-1:0] Wgt_1_116,input [WEIGHT_SIZE-1:0] Wgt_1_117,input [WEIGHT_SIZE-1:0] Wgt_1_118,input [WEIGHT_SIZE-1:0] Wgt_1_119,input [WEIGHT_SIZE-1:0] Wgt_1_120,input [WEIGHT_SIZE-1:0] Wgt_1_121,input [WEIGHT_SIZE-1:0] Wgt_1_122,input [WEIGHT_SIZE-1:0] Wgt_1_123,input [WEIGHT_SIZE-1:0] Wgt_1_124,input [WEIGHT_SIZE-1:0] Wgt_1_125,input [WEIGHT_SIZE-1:0] Wgt_1_126,input [WEIGHT_SIZE-1:0] Wgt_1_127,input [WEIGHT_SIZE-1:0] Wgt_1_128,input [WEIGHT_SIZE-1:0] Wgt_1_129,input [WEIGHT_SIZE-1:0] Wgt_1_130,input [WEIGHT_SIZE-1:0] Wgt_1_131,input [WEIGHT_SIZE-1:0] Wgt_1_132,input [WEIGHT_SIZE-1:0] Wgt_1_133,input [WEIGHT_SIZE-1:0] Wgt_1_134,input [WEIGHT_SIZE-1:0] Wgt_1_135,input [WEIGHT_SIZE-1:0] Wgt_1_136,input [WEIGHT_SIZE-1:0] Wgt_1_137,input [WEIGHT_SIZE-1:0] Wgt_1_138,input [WEIGHT_SIZE-1:0] Wgt_1_139,input [WEIGHT_SIZE-1:0] Wgt_1_140,input [WEIGHT_SIZE-1:0] Wgt_1_141,input [WEIGHT_SIZE-1:0] Wgt_1_142,input [WEIGHT_SIZE-1:0] Wgt_1_143,input [WEIGHT_SIZE-1:0] Wgt_1_144,input [WEIGHT_SIZE-1:0] Wgt_1_145,input [WEIGHT_SIZE-1:0] Wgt_1_146,input [WEIGHT_SIZE-1:0] Wgt_1_147,input [WEIGHT_SIZE-1:0] Wgt_1_148,input [WEIGHT_SIZE-1:0] Wgt_1_149,input [WEIGHT_SIZE-1:0] Wgt_1_150,input [WEIGHT_SIZE-1:0] Wgt_1_151,input [WEIGHT_SIZE-1:0] Wgt_1_152,input [WEIGHT_SIZE-1:0] Wgt_1_153,input [WEIGHT_SIZE-1:0] Wgt_1_154,input [WEIGHT_SIZE-1:0] Wgt_1_155,input [WEIGHT_SIZE-1:0] Wgt_1_156,input [WEIGHT_SIZE-1:0] Wgt_1_157,input [WEIGHT_SIZE-1:0] Wgt_1_158,input [WEIGHT_SIZE-1:0] Wgt_1_159,input [WEIGHT_SIZE-1:0] Wgt_1_160,input [WEIGHT_SIZE-1:0] Wgt_1_161,input [WEIGHT_SIZE-1:0] Wgt_1_162,input [WEIGHT_SIZE-1:0] Wgt_1_163,input [WEIGHT_SIZE-1:0] Wgt_1_164,input [WEIGHT_SIZE-1:0] Wgt_1_165,input [WEIGHT_SIZE-1:0] Wgt_1_166,input [WEIGHT_SIZE-1:0] Wgt_1_167,input [WEIGHT_SIZE-1:0] Wgt_1_168,input [WEIGHT_SIZE-1:0] Wgt_1_169,input [WEIGHT_SIZE-1:0] Wgt_1_170,input [WEIGHT_SIZE-1:0] Wgt_1_171,input [WEIGHT_SIZE-1:0] Wgt_1_172,input [WEIGHT_SIZE-1:0] Wgt_1_173,input [WEIGHT_SIZE-1:0] Wgt_1_174,input [WEIGHT_SIZE-1:0] Wgt_1_175,input [WEIGHT_SIZE-1:0] Wgt_1_176,input [WEIGHT_SIZE-1:0] Wgt_1_177,input [WEIGHT_SIZE-1:0] Wgt_1_178,input [WEIGHT_SIZE-1:0] Wgt_1_179,input [WEIGHT_SIZE-1:0] Wgt_1_180,input [WEIGHT_SIZE-1:0] Wgt_1_181,input [WEIGHT_SIZE-1:0] Wgt_1_182,input [WEIGHT_SIZE-1:0] Wgt_1_183,input [WEIGHT_SIZE-1:0] Wgt_1_184,input [WEIGHT_SIZE-1:0] Wgt_1_185,input [WEIGHT_SIZE-1:0] Wgt_1_186,input [WEIGHT_SIZE-1:0] Wgt_1_187,input [WEIGHT_SIZE-1:0] Wgt_1_188,input [WEIGHT_SIZE-1:0] Wgt_1_189,input [WEIGHT_SIZE-1:0] Wgt_1_190,input [WEIGHT_SIZE-1:0] Wgt_1_191,input [WEIGHT_SIZE-1:0] Wgt_1_192,input [WEIGHT_SIZE-1:0] Wgt_1_193,input [WEIGHT_SIZE-1:0] Wgt_1_194,input [WEIGHT_SIZE-1:0] Wgt_1_195,input [WEIGHT_SIZE-1:0] Wgt_1_196,input [WEIGHT_SIZE-1:0] Wgt_1_197,input [WEIGHT_SIZE-1:0] Wgt_1_198,input [WEIGHT_SIZE-1:0] Wgt_1_199,input [WEIGHT_SIZE-1:0] Wgt_1_200,input [WEIGHT_SIZE-1:0] Wgt_1_201,input [WEIGHT_SIZE-1:0] Wgt_1_202,input [WEIGHT_SIZE-1:0] Wgt_1_203,input [WEIGHT_SIZE-1:0] Wgt_1_204,input [WEIGHT_SIZE-1:0] Wgt_1_205,input [WEIGHT_SIZE-1:0] Wgt_1_206,input [WEIGHT_SIZE-1:0] Wgt_1_207,input [WEIGHT_SIZE-1:0] Wgt_1_208,input [WEIGHT_SIZE-1:0] Wgt_1_209,input [WEIGHT_SIZE-1:0] Wgt_1_210,input [WEIGHT_SIZE-1:0] Wgt_1_211,input [WEIGHT_SIZE-1:0] Wgt_1_212,input [WEIGHT_SIZE-1:0] Wgt_1_213,input [WEIGHT_SIZE-1:0] Wgt_1_214,input [WEIGHT_SIZE-1:0] Wgt_1_215,input [WEIGHT_SIZE-1:0] Wgt_1_216,input [WEIGHT_SIZE-1:0] Wgt_1_217,input [WEIGHT_SIZE-1:0] Wgt_1_218,input [WEIGHT_SIZE-1:0] Wgt_1_219,input [WEIGHT_SIZE-1:0] Wgt_1_220,input [WEIGHT_SIZE-1:0] Wgt_1_221,input [WEIGHT_SIZE-1:0] Wgt_1_222,input [WEIGHT_SIZE-1:0] Wgt_1_223,input [WEIGHT_SIZE-1:0] Wgt_1_224,input [WEIGHT_SIZE-1:0] Wgt_1_225,input [WEIGHT_SIZE-1:0] Wgt_1_226,input [WEIGHT_SIZE-1:0] Wgt_1_227,input [WEIGHT_SIZE-1:0] Wgt_1_228,input [WEIGHT_SIZE-1:0] Wgt_1_229,input [WEIGHT_SIZE-1:0] Wgt_1_230,input [WEIGHT_SIZE-1:0] Wgt_1_231,input [WEIGHT_SIZE-1:0] Wgt_1_232,input [WEIGHT_SIZE-1:0] Wgt_1_233,input [WEIGHT_SIZE-1:0] Wgt_1_234,input [WEIGHT_SIZE-1:0] Wgt_1_235,input [WEIGHT_SIZE-1:0] Wgt_1_236,input [WEIGHT_SIZE-1:0] Wgt_1_237,input [WEIGHT_SIZE-1:0] Wgt_1_238,input [WEIGHT_SIZE-1:0] Wgt_1_239,input [WEIGHT_SIZE-1:0] Wgt_1_240,input [WEIGHT_SIZE-1:0] Wgt_1_241,input [WEIGHT_SIZE-1:0] Wgt_1_242,input [WEIGHT_SIZE-1:0] Wgt_1_243,input [WEIGHT_SIZE-1:0] Wgt_1_244,input [WEIGHT_SIZE-1:0] Wgt_1_245,input [WEIGHT_SIZE-1:0] Wgt_1_246,input [WEIGHT_SIZE-1:0] Wgt_1_247,input [WEIGHT_SIZE-1:0] Wgt_1_248,input [WEIGHT_SIZE-1:0] Wgt_1_249,input [WEIGHT_SIZE-1:0] Wgt_1_250,input [WEIGHT_SIZE-1:0] Wgt_1_251,input [WEIGHT_SIZE-1:0] Wgt_1_252,input [WEIGHT_SIZE-1:0] Wgt_1_253,input [WEIGHT_SIZE-1:0] Wgt_1_254,input [WEIGHT_SIZE-1:0] Wgt_1_255,input [WEIGHT_SIZE-1:0] Wgt_1_256,input [WEIGHT_SIZE-1:0] Wgt_1_257,input [WEIGHT_SIZE-1:0] Wgt_1_258,input [WEIGHT_SIZE-1:0] Wgt_1_259,input [WEIGHT_SIZE-1:0] Wgt_1_260,input [WEIGHT_SIZE-1:0] Wgt_1_261,input [WEIGHT_SIZE-1:0] Wgt_1_262,input [WEIGHT_SIZE-1:0] Wgt_1_263,input [WEIGHT_SIZE-1:0] Wgt_1_264,input [WEIGHT_SIZE-1:0] Wgt_1_265,input [WEIGHT_SIZE-1:0] Wgt_1_266,input [WEIGHT_SIZE-1:0] Wgt_1_267,input [WEIGHT_SIZE-1:0] Wgt_1_268,input [WEIGHT_SIZE-1:0] Wgt_1_269,input [WEIGHT_SIZE-1:0] Wgt_1_270,input [WEIGHT_SIZE-1:0] Wgt_1_271,input [WEIGHT_SIZE-1:0] Wgt_1_272,input [WEIGHT_SIZE-1:0] Wgt_1_273,input [WEIGHT_SIZE-1:0] Wgt_1_274,input [WEIGHT_SIZE-1:0] Wgt_1_275,input [WEIGHT_SIZE-1:0] Wgt_1_276,input [WEIGHT_SIZE-1:0] Wgt_1_277,input [WEIGHT_SIZE-1:0] Wgt_1_278,input [WEIGHT_SIZE-1:0] Wgt_1_279,input [WEIGHT_SIZE-1:0] Wgt_1_280,input [WEIGHT_SIZE-1:0] Wgt_1_281,input [WEIGHT_SIZE-1:0] Wgt_1_282,input [WEIGHT_SIZE-1:0] Wgt_1_283,input [WEIGHT_SIZE-1:0] Wgt_1_284,input [WEIGHT_SIZE-1:0] Wgt_1_285,input [WEIGHT_SIZE-1:0] Wgt_1_286,input [WEIGHT_SIZE-1:0] Wgt_1_287,input [WEIGHT_SIZE-1:0] Wgt_1_288,input [WEIGHT_SIZE-1:0] Wgt_1_289,input [WEIGHT_SIZE-1:0] Wgt_1_290,input [WEIGHT_SIZE-1:0] Wgt_1_291,input [WEIGHT_SIZE-1:0] Wgt_1_292,input [WEIGHT_SIZE-1:0] Wgt_1_293,input [WEIGHT_SIZE-1:0] Wgt_1_294,input [WEIGHT_SIZE-1:0] Wgt_1_295,input [WEIGHT_SIZE-1:0] Wgt_1_296,input [WEIGHT_SIZE-1:0] Wgt_1_297,input [WEIGHT_SIZE-1:0] Wgt_1_298,input [WEIGHT_SIZE-1:0] Wgt_1_299,input [WEIGHT_SIZE-1:0] Wgt_1_300,input [WEIGHT_SIZE-1:0] Wgt_1_301,input [WEIGHT_SIZE-1:0] Wgt_1_302,input [WEIGHT_SIZE-1:0] Wgt_1_303,input [WEIGHT_SIZE-1:0] Wgt_1_304,input [WEIGHT_SIZE-1:0] Wgt_1_305,input [WEIGHT_SIZE-1:0] Wgt_1_306,input [WEIGHT_SIZE-1:0] Wgt_1_307,input [WEIGHT_SIZE-1:0] Wgt_1_308,input [WEIGHT_SIZE-1:0] Wgt_1_309,input [WEIGHT_SIZE-1:0] Wgt_1_310,input [WEIGHT_SIZE-1:0] Wgt_1_311,input [WEIGHT_SIZE-1:0] Wgt_1_312,input [WEIGHT_SIZE-1:0] Wgt_1_313,input [WEIGHT_SIZE-1:0] Wgt_1_314,input [WEIGHT_SIZE-1:0] Wgt_1_315,input [WEIGHT_SIZE-1:0] Wgt_1_316,input [WEIGHT_SIZE-1:0] Wgt_1_317,input [WEIGHT_SIZE-1:0] Wgt_1_318,input [WEIGHT_SIZE-1:0] Wgt_1_319,input [WEIGHT_SIZE-1:0] Wgt_1_320,input [WEIGHT_SIZE-1:0] Wgt_1_321,input [WEIGHT_SIZE-1:0] Wgt_1_322,input [WEIGHT_SIZE-1:0] Wgt_1_323,input [WEIGHT_SIZE-1:0] Wgt_1_324,input [WEIGHT_SIZE-1:0] Wgt_1_325,input [WEIGHT_SIZE-1:0] Wgt_1_326,input [WEIGHT_SIZE-1:0] Wgt_1_327,input [WEIGHT_SIZE-1:0] Wgt_1_328,input [WEIGHT_SIZE-1:0] Wgt_1_329,input [WEIGHT_SIZE-1:0] Wgt_1_330,input [WEIGHT_SIZE-1:0] Wgt_1_331,input [WEIGHT_SIZE-1:0] Wgt_1_332,input [WEIGHT_SIZE-1:0] Wgt_1_333,input [WEIGHT_SIZE-1:0] Wgt_1_334,input [WEIGHT_SIZE-1:0] Wgt_1_335,input [WEIGHT_SIZE-1:0] Wgt_1_336,input [WEIGHT_SIZE-1:0] Wgt_1_337,input [WEIGHT_SIZE-1:0] Wgt_1_338,input [WEIGHT_SIZE-1:0] Wgt_1_339,input [WEIGHT_SIZE-1:0] Wgt_1_340,input [WEIGHT_SIZE-1:0] Wgt_1_341,input [WEIGHT_SIZE-1:0] Wgt_1_342,input [WEIGHT_SIZE-1:0] Wgt_1_343,input [WEIGHT_SIZE-1:0] Wgt_1_344,input [WEIGHT_SIZE-1:0] Wgt_1_345,input [WEIGHT_SIZE-1:0] Wgt_1_346,input [WEIGHT_SIZE-1:0] Wgt_1_347,input [WEIGHT_SIZE-1:0] Wgt_1_348,input [WEIGHT_SIZE-1:0] Wgt_1_349,input [WEIGHT_SIZE-1:0] Wgt_1_350,input [WEIGHT_SIZE-1:0] Wgt_1_351,input [WEIGHT_SIZE-1:0] Wgt_1_352,input [WEIGHT_SIZE-1:0] Wgt_1_353,input [WEIGHT_SIZE-1:0] Wgt_1_354,input [WEIGHT_SIZE-1:0] Wgt_1_355,input [WEIGHT_SIZE-1:0] Wgt_1_356,input [WEIGHT_SIZE-1:0] Wgt_1_357,input [WEIGHT_SIZE-1:0] Wgt_1_358,input [WEIGHT_SIZE-1:0] Wgt_1_359,input [WEIGHT_SIZE-1:0] Wgt_1_360,input [WEIGHT_SIZE-1:0] Wgt_1_361,input [WEIGHT_SIZE-1:0] Wgt_1_362,input [WEIGHT_SIZE-1:0] Wgt_1_363,input [WEIGHT_SIZE-1:0] Wgt_1_364,input [WEIGHT_SIZE-1:0] Wgt_1_365,input [WEIGHT_SIZE-1:0] Wgt_1_366,input [WEIGHT_SIZE-1:0] Wgt_1_367,input [WEIGHT_SIZE-1:0] Wgt_1_368,input [WEIGHT_SIZE-1:0] Wgt_1_369,input [WEIGHT_SIZE-1:0] Wgt_1_370,input [WEIGHT_SIZE-1:0] Wgt_1_371,input [WEIGHT_SIZE-1:0] Wgt_1_372,input [WEIGHT_SIZE-1:0] Wgt_1_373,input [WEIGHT_SIZE-1:0] Wgt_1_374,input [WEIGHT_SIZE-1:0] Wgt_1_375,input [WEIGHT_SIZE-1:0] Wgt_1_376,input [WEIGHT_SIZE-1:0] Wgt_1_377,input [WEIGHT_SIZE-1:0] Wgt_1_378,input [WEIGHT_SIZE-1:0] Wgt_1_379,input [WEIGHT_SIZE-1:0] Wgt_1_380,input [WEIGHT_SIZE-1:0] Wgt_1_381,input [WEIGHT_SIZE-1:0] Wgt_1_382,input [WEIGHT_SIZE-1:0] Wgt_1_383,input [WEIGHT_SIZE-1:0] Wgt_1_384,input [WEIGHT_SIZE-1:0] Wgt_1_385,input [WEIGHT_SIZE-1:0] Wgt_1_386,input [WEIGHT_SIZE-1:0] Wgt_1_387,input [WEIGHT_SIZE-1:0] Wgt_1_388,input [WEIGHT_SIZE-1:0] Wgt_1_389,input [WEIGHT_SIZE-1:0] Wgt_1_390,input [WEIGHT_SIZE-1:0] Wgt_1_391,input [WEIGHT_SIZE-1:0] Wgt_1_392,input [WEIGHT_SIZE-1:0] Wgt_1_393,input [WEIGHT_SIZE-1:0] Wgt_1_394,input [WEIGHT_SIZE-1:0] Wgt_1_395,input [WEIGHT_SIZE-1:0] Wgt_1_396,input [WEIGHT_SIZE-1:0] Wgt_1_397,input [WEIGHT_SIZE-1:0] Wgt_1_398,input [WEIGHT_SIZE-1:0] Wgt_1_399,input [WEIGHT_SIZE-1:0] Wgt_1_400,input [WEIGHT_SIZE-1:0] Wgt_1_401,input [WEIGHT_SIZE-1:0] Wgt_1_402,input [WEIGHT_SIZE-1:0] Wgt_1_403,input [WEIGHT_SIZE-1:0] Wgt_1_404,input [WEIGHT_SIZE-1:0] Wgt_1_405,input [WEIGHT_SIZE-1:0] Wgt_1_406,input [WEIGHT_SIZE-1:0] Wgt_1_407,input [WEIGHT_SIZE-1:0] Wgt_1_408,input [WEIGHT_SIZE-1:0] Wgt_1_409,input [WEIGHT_SIZE-1:0] Wgt_1_410,input [WEIGHT_SIZE-1:0] Wgt_1_411,input [WEIGHT_SIZE-1:0] Wgt_1_412,input [WEIGHT_SIZE-1:0] Wgt_1_413,input [WEIGHT_SIZE-1:0] Wgt_1_414,input [WEIGHT_SIZE-1:0] Wgt_1_415,input [WEIGHT_SIZE-1:0] Wgt_1_416,input [WEIGHT_SIZE-1:0] Wgt_1_417,input [WEIGHT_SIZE-1:0] Wgt_1_418,input [WEIGHT_SIZE-1:0] Wgt_1_419,input [WEIGHT_SIZE-1:0] Wgt_1_420,input [WEIGHT_SIZE-1:0] Wgt_1_421,input [WEIGHT_SIZE-1:0] Wgt_1_422,input [WEIGHT_SIZE-1:0] Wgt_1_423,input [WEIGHT_SIZE-1:0] Wgt_1_424,input [WEIGHT_SIZE-1:0] Wgt_1_425,input [WEIGHT_SIZE-1:0] Wgt_1_426,input [WEIGHT_SIZE-1:0] Wgt_1_427,input [WEIGHT_SIZE-1:0] Wgt_1_428,input [WEIGHT_SIZE-1:0] Wgt_1_429,input [WEIGHT_SIZE-1:0] Wgt_1_430,input [WEIGHT_SIZE-1:0] Wgt_1_431,input [WEIGHT_SIZE-1:0] Wgt_1_432,input [WEIGHT_SIZE-1:0] Wgt_1_433,input [WEIGHT_SIZE-1:0] Wgt_1_434,input [WEIGHT_SIZE-1:0] Wgt_1_435,input [WEIGHT_SIZE-1:0] Wgt_1_436,input [WEIGHT_SIZE-1:0] Wgt_1_437,input [WEIGHT_SIZE-1:0] Wgt_1_438,input [WEIGHT_SIZE-1:0] Wgt_1_439,input [WEIGHT_SIZE-1:0] Wgt_1_440,input [WEIGHT_SIZE-1:0] Wgt_1_441,input [WEIGHT_SIZE-1:0] Wgt_1_442,input [WEIGHT_SIZE-1:0] Wgt_1_443,input [WEIGHT_SIZE-1:0] Wgt_1_444,input [WEIGHT_SIZE-1:0] Wgt_1_445,input [WEIGHT_SIZE-1:0] Wgt_1_446,input [WEIGHT_SIZE-1:0] Wgt_1_447,input [WEIGHT_SIZE-1:0] Wgt_1_448,input [WEIGHT_SIZE-1:0] Wgt_1_449,input [WEIGHT_SIZE-1:0] Wgt_1_450,input [WEIGHT_SIZE-1:0] Wgt_1_451,input [WEIGHT_SIZE-1:0] Wgt_1_452,input [WEIGHT_SIZE-1:0] Wgt_1_453,input [WEIGHT_SIZE-1:0] Wgt_1_454,input [WEIGHT_SIZE-1:0] Wgt_1_455,input [WEIGHT_SIZE-1:0] Wgt_1_456,input [WEIGHT_SIZE-1:0] Wgt_1_457,input [WEIGHT_SIZE-1:0] Wgt_1_458,input [WEIGHT_SIZE-1:0] Wgt_1_459,input [WEIGHT_SIZE-1:0] Wgt_1_460,input [WEIGHT_SIZE-1:0] Wgt_1_461,input [WEIGHT_SIZE-1:0] Wgt_1_462,input [WEIGHT_SIZE-1:0] Wgt_1_463,input [WEIGHT_SIZE-1:0] Wgt_1_464,input [WEIGHT_SIZE-1:0] Wgt_1_465,input [WEIGHT_SIZE-1:0] Wgt_1_466,input [WEIGHT_SIZE-1:0] Wgt_1_467,input [WEIGHT_SIZE-1:0] Wgt_1_468,input [WEIGHT_SIZE-1:0] Wgt_1_469,input [WEIGHT_SIZE-1:0] Wgt_1_470,input [WEIGHT_SIZE-1:0] Wgt_1_471,input [WEIGHT_SIZE-1:0] Wgt_1_472,input [WEIGHT_SIZE-1:0] Wgt_1_473,input [WEIGHT_SIZE-1:0] Wgt_1_474,input [WEIGHT_SIZE-1:0] Wgt_1_475,input [WEIGHT_SIZE-1:0] Wgt_1_476,input [WEIGHT_SIZE-1:0] Wgt_1_477,input [WEIGHT_SIZE-1:0] Wgt_1_478,input [WEIGHT_SIZE-1:0] Wgt_1_479,input [WEIGHT_SIZE-1:0] Wgt_1_480,input [WEIGHT_SIZE-1:0] Wgt_1_481,input [WEIGHT_SIZE-1:0] Wgt_1_482,input [WEIGHT_SIZE-1:0] Wgt_1_483,input [WEIGHT_SIZE-1:0] Wgt_1_484,input [WEIGHT_SIZE-1:0] Wgt_1_485,input [WEIGHT_SIZE-1:0] Wgt_1_486,input [WEIGHT_SIZE-1:0] Wgt_1_487,input [WEIGHT_SIZE-1:0] Wgt_1_488,input [WEIGHT_SIZE-1:0] Wgt_1_489,input [WEIGHT_SIZE-1:0] Wgt_1_490,input [WEIGHT_SIZE-1:0] Wgt_1_491,input [WEIGHT_SIZE-1:0] Wgt_1_492,input [WEIGHT_SIZE-1:0] Wgt_1_493,input [WEIGHT_SIZE-1:0] Wgt_1_494,input [WEIGHT_SIZE-1:0] Wgt_1_495,input [WEIGHT_SIZE-1:0] Wgt_1_496,input [WEIGHT_SIZE-1:0] Wgt_1_497,input [WEIGHT_SIZE-1:0] Wgt_1_498,input [WEIGHT_SIZE-1:0] Wgt_1_499,input [WEIGHT_SIZE-1:0] Wgt_1_500,input [WEIGHT_SIZE-1:0] Wgt_1_501,input [WEIGHT_SIZE-1:0] Wgt_1_502,input [WEIGHT_SIZE-1:0] Wgt_1_503,input [WEIGHT_SIZE-1:0] Wgt_1_504,input [WEIGHT_SIZE-1:0] Wgt_1_505,input [WEIGHT_SIZE-1:0] Wgt_1_506,input [WEIGHT_SIZE-1:0] Wgt_1_507,input [WEIGHT_SIZE-1:0] Wgt_1_508,input [WEIGHT_SIZE-1:0] Wgt_1_509,input [WEIGHT_SIZE-1:0] Wgt_1_510,input [WEIGHT_SIZE-1:0] Wgt_1_511,input [WEIGHT_SIZE-1:0] Wgt_1_512,input [WEIGHT_SIZE-1:0] Wgt_1_513,input [WEIGHT_SIZE-1:0] Wgt_1_514,input [WEIGHT_SIZE-1:0] Wgt_1_515,input [WEIGHT_SIZE-1:0] Wgt_1_516,input [WEIGHT_SIZE-1:0] Wgt_1_517,input [WEIGHT_SIZE-1:0] Wgt_1_518,input [WEIGHT_SIZE-1:0] Wgt_1_519,input [WEIGHT_SIZE-1:0] Wgt_1_520,input [WEIGHT_SIZE-1:0] Wgt_1_521,input [WEIGHT_SIZE-1:0] Wgt_1_522,input [WEIGHT_SIZE-1:0] Wgt_1_523,input [WEIGHT_SIZE-1:0] Wgt_1_524,input [WEIGHT_SIZE-1:0] Wgt_1_525,input [WEIGHT_SIZE-1:0] Wgt_1_526,input [WEIGHT_SIZE-1:0] Wgt_1_527,input [WEIGHT_SIZE-1:0] Wgt_1_528,input [WEIGHT_SIZE-1:0] Wgt_1_529,input [WEIGHT_SIZE-1:0] Wgt_1_530,input [WEIGHT_SIZE-1:0] Wgt_1_531,input [WEIGHT_SIZE-1:0] Wgt_1_532,input [WEIGHT_SIZE-1:0] Wgt_1_533,input [WEIGHT_SIZE-1:0] Wgt_1_534,input [WEIGHT_SIZE-1:0] Wgt_1_535,input [WEIGHT_SIZE-1:0] Wgt_1_536,input [WEIGHT_SIZE-1:0] Wgt_1_537,input [WEIGHT_SIZE-1:0] Wgt_1_538,input [WEIGHT_SIZE-1:0] Wgt_1_539,input [WEIGHT_SIZE-1:0] Wgt_1_540,input [WEIGHT_SIZE-1:0] Wgt_1_541,input [WEIGHT_SIZE-1:0] Wgt_1_542,input [WEIGHT_SIZE-1:0] Wgt_1_543,input [WEIGHT_SIZE-1:0] Wgt_1_544,input [WEIGHT_SIZE-1:0] Wgt_1_545,input [WEIGHT_SIZE-1:0] Wgt_1_546,input [WEIGHT_SIZE-1:0] Wgt_1_547,input [WEIGHT_SIZE-1:0] Wgt_1_548,input [WEIGHT_SIZE-1:0] Wgt_1_549,input [WEIGHT_SIZE-1:0] Wgt_1_550,input [WEIGHT_SIZE-1:0] Wgt_1_551,input [WEIGHT_SIZE-1:0] Wgt_1_552,input [WEIGHT_SIZE-1:0] Wgt_1_553,input [WEIGHT_SIZE-1:0] Wgt_1_554,input [WEIGHT_SIZE-1:0] Wgt_1_555,input [WEIGHT_SIZE-1:0] Wgt_1_556,input [WEIGHT_SIZE-1:0] Wgt_1_557,input [WEIGHT_SIZE-1:0] Wgt_1_558,input [WEIGHT_SIZE-1:0] Wgt_1_559,input [WEIGHT_SIZE-1:0] Wgt_1_560,input [WEIGHT_SIZE-1:0] Wgt_1_561,input [WEIGHT_SIZE-1:0] Wgt_1_562,input [WEIGHT_SIZE-1:0] Wgt_1_563,input [WEIGHT_SIZE-1:0] Wgt_1_564,input [WEIGHT_SIZE-1:0] Wgt_1_565,input [WEIGHT_SIZE-1:0] Wgt_1_566,input [WEIGHT_SIZE-1:0] Wgt_1_567,input [WEIGHT_SIZE-1:0] Wgt_1_568,input [WEIGHT_SIZE-1:0] Wgt_1_569,input [WEIGHT_SIZE-1:0] Wgt_1_570,input [WEIGHT_SIZE-1:0] Wgt_1_571,input [WEIGHT_SIZE-1:0] Wgt_1_572,input [WEIGHT_SIZE-1:0] Wgt_1_573,input [WEIGHT_SIZE-1:0] Wgt_1_574,input [WEIGHT_SIZE-1:0] Wgt_1_575,input [WEIGHT_SIZE-1:0] Wgt_1_576,input [WEIGHT_SIZE-1:0] Wgt_1_577,input [WEIGHT_SIZE-1:0] Wgt_1_578,input [WEIGHT_SIZE-1:0] Wgt_1_579,input [WEIGHT_SIZE-1:0] Wgt_1_580,input [WEIGHT_SIZE-1:0] Wgt_1_581,input [WEIGHT_SIZE-1:0] Wgt_1_582,input [WEIGHT_SIZE-1:0] Wgt_1_583,input [WEIGHT_SIZE-1:0] Wgt_1_584,input [WEIGHT_SIZE-1:0] Wgt_1_585,input [WEIGHT_SIZE-1:0] Wgt_1_586,input [WEIGHT_SIZE-1:0] Wgt_1_587,input [WEIGHT_SIZE-1:0] Wgt_1_588,input [WEIGHT_SIZE-1:0] Wgt_1_589,input [WEIGHT_SIZE-1:0] Wgt_1_590,input [WEIGHT_SIZE-1:0] Wgt_1_591,input [WEIGHT_SIZE-1:0] Wgt_1_592,input [WEIGHT_SIZE-1:0] Wgt_1_593,input [WEIGHT_SIZE-1:0] Wgt_1_594,input [WEIGHT_SIZE-1:0] Wgt_1_595,input [WEIGHT_SIZE-1:0] Wgt_1_596,input [WEIGHT_SIZE-1:0] Wgt_1_597,input [WEIGHT_SIZE-1:0] Wgt_1_598,input [WEIGHT_SIZE-1:0] Wgt_1_599,input [WEIGHT_SIZE-1:0] Wgt_1_600,input [WEIGHT_SIZE-1:0] Wgt_1_601,input [WEIGHT_SIZE-1:0] Wgt_1_602,input [WEIGHT_SIZE-1:0] Wgt_1_603,input [WEIGHT_SIZE-1:0] Wgt_1_604,input [WEIGHT_SIZE-1:0] Wgt_1_605,input [WEIGHT_SIZE-1:0] Wgt_1_606,input [WEIGHT_SIZE-1:0] Wgt_1_607,input [WEIGHT_SIZE-1:0] Wgt_1_608,input [WEIGHT_SIZE-1:0] Wgt_1_609,input [WEIGHT_SIZE-1:0] Wgt_1_610,input [WEIGHT_SIZE-1:0] Wgt_1_611,input [WEIGHT_SIZE-1:0] Wgt_1_612,input [WEIGHT_SIZE-1:0] Wgt_1_613,input [WEIGHT_SIZE-1:0] Wgt_1_614,input [WEIGHT_SIZE-1:0] Wgt_1_615,input [WEIGHT_SIZE-1:0] Wgt_1_616,input [WEIGHT_SIZE-1:0] Wgt_1_617,input [WEIGHT_SIZE-1:0] Wgt_1_618,input [WEIGHT_SIZE-1:0] Wgt_1_619,input [WEIGHT_SIZE-1:0] Wgt_1_620,input [WEIGHT_SIZE-1:0] Wgt_1_621,input [WEIGHT_SIZE-1:0] Wgt_1_622,input [WEIGHT_SIZE-1:0] Wgt_1_623,input [WEIGHT_SIZE-1:0] Wgt_1_624,input [WEIGHT_SIZE-1:0] Wgt_1_625,input [WEIGHT_SIZE-1:0] Wgt_1_626,input [WEIGHT_SIZE-1:0] Wgt_1_627,input [WEIGHT_SIZE-1:0] Wgt_1_628,input [WEIGHT_SIZE-1:0] Wgt_1_629,input [WEIGHT_SIZE-1:0] Wgt_1_630,input [WEIGHT_SIZE-1:0] Wgt_1_631,input [WEIGHT_SIZE-1:0] Wgt_1_632,input [WEIGHT_SIZE-1:0] Wgt_1_633,input [WEIGHT_SIZE-1:0] Wgt_1_634,input [WEIGHT_SIZE-1:0] Wgt_1_635,input [WEIGHT_SIZE-1:0] Wgt_1_636,input [WEIGHT_SIZE-1:0] Wgt_1_637,input [WEIGHT_SIZE-1:0] Wgt_1_638,input [WEIGHT_SIZE-1:0] Wgt_1_639,input [WEIGHT_SIZE-1:0] Wgt_1_640,input [WEIGHT_SIZE-1:0] Wgt_1_641,input [WEIGHT_SIZE-1:0] Wgt_1_642,input [WEIGHT_SIZE-1:0] Wgt_1_643,input [WEIGHT_SIZE-1:0] Wgt_1_644,input [WEIGHT_SIZE-1:0] Wgt_1_645,input [WEIGHT_SIZE-1:0] Wgt_1_646,input [WEIGHT_SIZE-1:0] Wgt_1_647,input [WEIGHT_SIZE-1:0] Wgt_1_648,input [WEIGHT_SIZE-1:0] Wgt_1_649,input [WEIGHT_SIZE-1:0] Wgt_1_650,input [WEIGHT_SIZE-1:0] Wgt_1_651,input [WEIGHT_SIZE-1:0] Wgt_1_652,input [WEIGHT_SIZE-1:0] Wgt_1_653,input [WEIGHT_SIZE-1:0] Wgt_1_654,input [WEIGHT_SIZE-1:0] Wgt_1_655,input [WEIGHT_SIZE-1:0] Wgt_1_656,input [WEIGHT_SIZE-1:0] Wgt_1_657,input [WEIGHT_SIZE-1:0] Wgt_1_658,input [WEIGHT_SIZE-1:0] Wgt_1_659,input [WEIGHT_SIZE-1:0] Wgt_1_660,input [WEIGHT_SIZE-1:0] Wgt_1_661,input [WEIGHT_SIZE-1:0] Wgt_1_662,input [WEIGHT_SIZE-1:0] Wgt_1_663,input [WEIGHT_SIZE-1:0] Wgt_1_664,input [WEIGHT_SIZE-1:0] Wgt_1_665,input [WEIGHT_SIZE-1:0] Wgt_1_666,input [WEIGHT_SIZE-1:0] Wgt_1_667,input [WEIGHT_SIZE-1:0] Wgt_1_668,input [WEIGHT_SIZE-1:0] Wgt_1_669,input [WEIGHT_SIZE-1:0] Wgt_1_670,input [WEIGHT_SIZE-1:0] Wgt_1_671,input [WEIGHT_SIZE-1:0] Wgt_1_672,input [WEIGHT_SIZE-1:0] Wgt_1_673,input [WEIGHT_SIZE-1:0] Wgt_1_674,input [WEIGHT_SIZE-1:0] Wgt_1_675,input [WEIGHT_SIZE-1:0] Wgt_1_676,input [WEIGHT_SIZE-1:0] Wgt_1_677,input [WEIGHT_SIZE-1:0] Wgt_1_678,input [WEIGHT_SIZE-1:0] Wgt_1_679,input [WEIGHT_SIZE-1:0] Wgt_1_680,input [WEIGHT_SIZE-1:0] Wgt_1_681,input [WEIGHT_SIZE-1:0] Wgt_1_682,input [WEIGHT_SIZE-1:0] Wgt_1_683,input [WEIGHT_SIZE-1:0] Wgt_1_684,input [WEIGHT_SIZE-1:0] Wgt_1_685,input [WEIGHT_SIZE-1:0] Wgt_1_686,input [WEIGHT_SIZE-1:0] Wgt_1_687,input [WEIGHT_SIZE-1:0] Wgt_1_688,input [WEIGHT_SIZE-1:0] Wgt_1_689,input [WEIGHT_SIZE-1:0] Wgt_1_690,input [WEIGHT_SIZE-1:0] Wgt_1_691,input [WEIGHT_SIZE-1:0] Wgt_1_692,input [WEIGHT_SIZE-1:0] Wgt_1_693,input [WEIGHT_SIZE-1:0] Wgt_1_694,input [WEIGHT_SIZE-1:0] Wgt_1_695,input [WEIGHT_SIZE-1:0] Wgt_1_696,input [WEIGHT_SIZE-1:0] Wgt_1_697,input [WEIGHT_SIZE-1:0] Wgt_1_698,input [WEIGHT_SIZE-1:0] Wgt_1_699,input [WEIGHT_SIZE-1:0] Wgt_1_700,input [WEIGHT_SIZE-1:0] Wgt_1_701,input [WEIGHT_SIZE-1:0] Wgt_1_702,input [WEIGHT_SIZE-1:0] Wgt_1_703,input [WEIGHT_SIZE-1:0] Wgt_1_704,input [WEIGHT_SIZE-1:0] Wgt_1_705,input [WEIGHT_SIZE-1:0] Wgt_1_706,input [WEIGHT_SIZE-1:0] Wgt_1_707,input [WEIGHT_SIZE-1:0] Wgt_1_708,input [WEIGHT_SIZE-1:0] Wgt_1_709,input [WEIGHT_SIZE-1:0] Wgt_1_710,input [WEIGHT_SIZE-1:0] Wgt_1_711,input [WEIGHT_SIZE-1:0] Wgt_1_712,input [WEIGHT_SIZE-1:0] Wgt_1_713,input [WEIGHT_SIZE-1:0] Wgt_1_714,input [WEIGHT_SIZE-1:0] Wgt_1_715,input [WEIGHT_SIZE-1:0] Wgt_1_716,input [WEIGHT_SIZE-1:0] Wgt_1_717,input [WEIGHT_SIZE-1:0] Wgt_1_718,input [WEIGHT_SIZE-1:0] Wgt_1_719,input [WEIGHT_SIZE-1:0] Wgt_1_720,input [WEIGHT_SIZE-1:0] Wgt_1_721,input [WEIGHT_SIZE-1:0] Wgt_1_722,input [WEIGHT_SIZE-1:0] Wgt_1_723,input [WEIGHT_SIZE-1:0] Wgt_1_724,input [WEIGHT_SIZE-1:0] Wgt_1_725,input [WEIGHT_SIZE-1:0] Wgt_1_726,input [WEIGHT_SIZE-1:0] Wgt_1_727,input [WEIGHT_SIZE-1:0] Wgt_1_728,input [WEIGHT_SIZE-1:0] Wgt_1_729,input [WEIGHT_SIZE-1:0] Wgt_1_730,input [WEIGHT_SIZE-1:0] Wgt_1_731,input [WEIGHT_SIZE-1:0] Wgt_1_732,input [WEIGHT_SIZE-1:0] Wgt_1_733,input [WEIGHT_SIZE-1:0] Wgt_1_734,input [WEIGHT_SIZE-1:0] Wgt_1_735,input [WEIGHT_SIZE-1:0] Wgt_1_736,input [WEIGHT_SIZE-1:0] Wgt_1_737,input [WEIGHT_SIZE-1:0] Wgt_1_738,input [WEIGHT_SIZE-1:0] Wgt_1_739,input [WEIGHT_SIZE-1:0] Wgt_1_740,input [WEIGHT_SIZE-1:0] Wgt_1_741,input [WEIGHT_SIZE-1:0] Wgt_1_742,input [WEIGHT_SIZE-1:0] Wgt_1_743,input [WEIGHT_SIZE-1:0] Wgt_1_744,input [WEIGHT_SIZE-1:0] Wgt_1_745,input [WEIGHT_SIZE-1:0] Wgt_1_746,input [WEIGHT_SIZE-1:0] Wgt_1_747,input [WEIGHT_SIZE-1:0] Wgt_1_748,input [WEIGHT_SIZE-1:0] Wgt_1_749,input [WEIGHT_SIZE-1:0] Wgt_1_750,input [WEIGHT_SIZE-1:0] Wgt_1_751,input [WEIGHT_SIZE-1:0] Wgt_1_752,input [WEIGHT_SIZE-1:0] Wgt_1_753,input [WEIGHT_SIZE-1:0] Wgt_1_754,input [WEIGHT_SIZE-1:0] Wgt_1_755,input [WEIGHT_SIZE-1:0] Wgt_1_756,input [WEIGHT_SIZE-1:0] Wgt_1_757,input [WEIGHT_SIZE-1:0] Wgt_1_758,input [WEIGHT_SIZE-1:0] Wgt_1_759,input [WEIGHT_SIZE-1:0] Wgt_1_760,input [WEIGHT_SIZE-1:0] Wgt_1_761,input [WEIGHT_SIZE-1:0] Wgt_1_762,input [WEIGHT_SIZE-1:0] Wgt_1_763,input [WEIGHT_SIZE-1:0] Wgt_1_764,input [WEIGHT_SIZE-1:0] Wgt_1_765,input [WEIGHT_SIZE-1:0] Wgt_1_766,input [WEIGHT_SIZE-1:0] Wgt_1_767,input [WEIGHT_SIZE-1:0] Wgt_1_768,input [WEIGHT_SIZE-1:0] Wgt_1_769,input [WEIGHT_SIZE-1:0] Wgt_1_770,input [WEIGHT_SIZE-1:0] Wgt_1_771,input [WEIGHT_SIZE-1:0] Wgt_1_772,input [WEIGHT_SIZE-1:0] Wgt_1_773,input [WEIGHT_SIZE-1:0] Wgt_1_774,input [WEIGHT_SIZE-1:0] Wgt_1_775,input [WEIGHT_SIZE-1:0] Wgt_1_776,input [WEIGHT_SIZE-1:0] Wgt_1_777,input [WEIGHT_SIZE-1:0] Wgt_1_778,input [WEIGHT_SIZE-1:0] Wgt_1_779,input [WEIGHT_SIZE-1:0] Wgt_1_780,input [WEIGHT_SIZE-1:0] Wgt_1_781,input [WEIGHT_SIZE-1:0] Wgt_1_782,input [WEIGHT_SIZE-1:0] Wgt_1_783,input [WEIGHT_SIZE-1:0] Wgt_1_784,input [WEIGHT_SIZE-1:0] Wgt_2_0,input [WEIGHT_SIZE-1:0] Wgt_2_1,input [WEIGHT_SIZE-1:0] Wgt_2_2,input [WEIGHT_SIZE-1:0] Wgt_2_3,input [WEIGHT_SIZE-1:0] Wgt_2_4,input [WEIGHT_SIZE-1:0] Wgt_2_5,input [WEIGHT_SIZE-1:0] Wgt_2_6,input [WEIGHT_SIZE-1:0] Wgt_2_7,input [WEIGHT_SIZE-1:0] Wgt_2_8,input [WEIGHT_SIZE-1:0] Wgt_2_9,input [WEIGHT_SIZE-1:0] Wgt_2_10,input [WEIGHT_SIZE-1:0] Wgt_2_11,input [WEIGHT_SIZE-1:0] Wgt_2_12,input [WEIGHT_SIZE-1:0] Wgt_2_13,input [WEIGHT_SIZE-1:0] Wgt_2_14,input [WEIGHT_SIZE-1:0] Wgt_2_15,input [WEIGHT_SIZE-1:0] Wgt_2_16,input [WEIGHT_SIZE-1:0] Wgt_2_17,input [WEIGHT_SIZE-1:0] Wgt_2_18,input [WEIGHT_SIZE-1:0] Wgt_2_19,input [WEIGHT_SIZE-1:0] Wgt_2_20,input [WEIGHT_SIZE-1:0] Wgt_2_21,input [WEIGHT_SIZE-1:0] Wgt_2_22,input [WEIGHT_SIZE-1:0] Wgt_2_23,input [WEIGHT_SIZE-1:0] Wgt_2_24,input [WEIGHT_SIZE-1:0] Wgt_2_25,input [WEIGHT_SIZE-1:0] Wgt_2_26,input [WEIGHT_SIZE-1:0] Wgt_2_27,input [WEIGHT_SIZE-1:0] Wgt_2_28,input [WEIGHT_SIZE-1:0] Wgt_2_29,input [WEIGHT_SIZE-1:0] Wgt_2_30,input [WEIGHT_SIZE-1:0] Wgt_2_31,input [WEIGHT_SIZE-1:0] Wgt_2_32,input [WEIGHT_SIZE-1:0] Wgt_2_33,input [WEIGHT_SIZE-1:0] Wgt_2_34,input [WEIGHT_SIZE-1:0] Wgt_2_35,input [WEIGHT_SIZE-1:0] Wgt_2_36,input [WEIGHT_SIZE-1:0] Wgt_2_37,input [WEIGHT_SIZE-1:0] Wgt_2_38,input [WEIGHT_SIZE-1:0] Wgt_2_39,input [WEIGHT_SIZE-1:0] Wgt_2_40,input [WEIGHT_SIZE-1:0] Wgt_2_41,input [WEIGHT_SIZE-1:0] Wgt_2_42,input [WEIGHT_SIZE-1:0] Wgt_2_43,input [WEIGHT_SIZE-1:0] Wgt_2_44,input [WEIGHT_SIZE-1:0] Wgt_2_45,input [WEIGHT_SIZE-1:0] Wgt_2_46,input [WEIGHT_SIZE-1:0] Wgt_2_47,input [WEIGHT_SIZE-1:0] Wgt_2_48,input [WEIGHT_SIZE-1:0] Wgt_2_49,input [WEIGHT_SIZE-1:0] Wgt_2_50,input [WEIGHT_SIZE-1:0] Wgt_2_51,input [WEIGHT_SIZE-1:0] Wgt_2_52,input [WEIGHT_SIZE-1:0] Wgt_2_53,input [WEIGHT_SIZE-1:0] Wgt_2_54,input [WEIGHT_SIZE-1:0] Wgt_2_55,input [WEIGHT_SIZE-1:0] Wgt_2_56,input [WEIGHT_SIZE-1:0] Wgt_2_57,input [WEIGHT_SIZE-1:0] Wgt_2_58,input [WEIGHT_SIZE-1:0] Wgt_2_59,input [WEIGHT_SIZE-1:0] Wgt_2_60,input [WEIGHT_SIZE-1:0] Wgt_2_61,input [WEIGHT_SIZE-1:0] Wgt_2_62,input [WEIGHT_SIZE-1:0] Wgt_2_63,input [WEIGHT_SIZE-1:0] Wgt_2_64,input [WEIGHT_SIZE-1:0] Wgt_2_65,input [WEIGHT_SIZE-1:0] Wgt_2_66,input [WEIGHT_SIZE-1:0] Wgt_2_67,input [WEIGHT_SIZE-1:0] Wgt_2_68,input [WEIGHT_SIZE-1:0] Wgt_2_69,input [WEIGHT_SIZE-1:0] Wgt_2_70,input [WEIGHT_SIZE-1:0] Wgt_2_71,input [WEIGHT_SIZE-1:0] Wgt_2_72,input [WEIGHT_SIZE-1:0] Wgt_2_73,input [WEIGHT_SIZE-1:0] Wgt_2_74,input [WEIGHT_SIZE-1:0] Wgt_2_75,input [WEIGHT_SIZE-1:0] Wgt_2_76,input [WEIGHT_SIZE-1:0] Wgt_2_77,input [WEIGHT_SIZE-1:0] Wgt_2_78,input [WEIGHT_SIZE-1:0] Wgt_2_79,input [WEIGHT_SIZE-1:0] Wgt_2_80,input [WEIGHT_SIZE-1:0] Wgt_2_81,input [WEIGHT_SIZE-1:0] Wgt_2_82,input [WEIGHT_SIZE-1:0] Wgt_2_83,input [WEIGHT_SIZE-1:0] Wgt_2_84,input [WEIGHT_SIZE-1:0] Wgt_2_85,input [WEIGHT_SIZE-1:0] Wgt_2_86,input [WEIGHT_SIZE-1:0] Wgt_2_87,input [WEIGHT_SIZE-1:0] Wgt_2_88,input [WEIGHT_SIZE-1:0] Wgt_2_89,input [WEIGHT_SIZE-1:0] Wgt_2_90,input [WEIGHT_SIZE-1:0] Wgt_2_91,input [WEIGHT_SIZE-1:0] Wgt_2_92,input [WEIGHT_SIZE-1:0] Wgt_2_93,input [WEIGHT_SIZE-1:0] Wgt_2_94,input [WEIGHT_SIZE-1:0] Wgt_2_95,input [WEIGHT_SIZE-1:0] Wgt_2_96,input [WEIGHT_SIZE-1:0] Wgt_2_97,input [WEIGHT_SIZE-1:0] Wgt_2_98,input [WEIGHT_SIZE-1:0] Wgt_2_99,input [WEIGHT_SIZE-1:0] Wgt_2_100,input [WEIGHT_SIZE-1:0] Wgt_2_101,input [WEIGHT_SIZE-1:0] Wgt_2_102,input [WEIGHT_SIZE-1:0] Wgt_2_103,input [WEIGHT_SIZE-1:0] Wgt_2_104,input [WEIGHT_SIZE-1:0] Wgt_2_105,input [WEIGHT_SIZE-1:0] Wgt_2_106,input [WEIGHT_SIZE-1:0] Wgt_2_107,input [WEIGHT_SIZE-1:0] Wgt_2_108,input [WEIGHT_SIZE-1:0] Wgt_2_109,input [WEIGHT_SIZE-1:0] Wgt_2_110,input [WEIGHT_SIZE-1:0] Wgt_2_111,input [WEIGHT_SIZE-1:0] Wgt_2_112,input [WEIGHT_SIZE-1:0] Wgt_2_113,input [WEIGHT_SIZE-1:0] Wgt_2_114,input [WEIGHT_SIZE-1:0] Wgt_2_115,input [WEIGHT_SIZE-1:0] Wgt_2_116,input [WEIGHT_SIZE-1:0] Wgt_2_117,input [WEIGHT_SIZE-1:0] Wgt_2_118,input [WEIGHT_SIZE-1:0] Wgt_2_119,input [WEIGHT_SIZE-1:0] Wgt_2_120,input [WEIGHT_SIZE-1:0] Wgt_2_121,input [WEIGHT_SIZE-1:0] Wgt_2_122,input [WEIGHT_SIZE-1:0] Wgt_2_123,input [WEIGHT_SIZE-1:0] Wgt_2_124,input [WEIGHT_SIZE-1:0] Wgt_2_125,input [WEIGHT_SIZE-1:0] Wgt_2_126,input [WEIGHT_SIZE-1:0] Wgt_2_127,input [WEIGHT_SIZE-1:0] Wgt_2_128,input [WEIGHT_SIZE-1:0] Wgt_2_129,input [WEIGHT_SIZE-1:0] Wgt_2_130,input [WEIGHT_SIZE-1:0] Wgt_2_131,input [WEIGHT_SIZE-1:0] Wgt_2_132,input [WEIGHT_SIZE-1:0] Wgt_2_133,input [WEIGHT_SIZE-1:0] Wgt_2_134,input [WEIGHT_SIZE-1:0] Wgt_2_135,input [WEIGHT_SIZE-1:0] Wgt_2_136,input [WEIGHT_SIZE-1:0] Wgt_2_137,input [WEIGHT_SIZE-1:0] Wgt_2_138,input [WEIGHT_SIZE-1:0] Wgt_2_139,input [WEIGHT_SIZE-1:0] Wgt_2_140,input [WEIGHT_SIZE-1:0] Wgt_2_141,input [WEIGHT_SIZE-1:0] Wgt_2_142,input [WEIGHT_SIZE-1:0] Wgt_2_143,input [WEIGHT_SIZE-1:0] Wgt_2_144,input [WEIGHT_SIZE-1:0] Wgt_2_145,input [WEIGHT_SIZE-1:0] Wgt_2_146,input [WEIGHT_SIZE-1:0] Wgt_2_147,input [WEIGHT_SIZE-1:0] Wgt_2_148,input [WEIGHT_SIZE-1:0] Wgt_2_149,input [WEIGHT_SIZE-1:0] Wgt_2_150,input [WEIGHT_SIZE-1:0] Wgt_2_151,input [WEIGHT_SIZE-1:0] Wgt_2_152,input [WEIGHT_SIZE-1:0] Wgt_2_153,input [WEIGHT_SIZE-1:0] Wgt_2_154,input [WEIGHT_SIZE-1:0] Wgt_2_155,input [WEIGHT_SIZE-1:0] Wgt_2_156,input [WEIGHT_SIZE-1:0] Wgt_2_157,input [WEIGHT_SIZE-1:0] Wgt_2_158,input [WEIGHT_SIZE-1:0] Wgt_2_159,input [WEIGHT_SIZE-1:0] Wgt_2_160,input [WEIGHT_SIZE-1:0] Wgt_2_161,input [WEIGHT_SIZE-1:0] Wgt_2_162,input [WEIGHT_SIZE-1:0] Wgt_2_163,input [WEIGHT_SIZE-1:0] Wgt_2_164,input [WEIGHT_SIZE-1:0] Wgt_2_165,input [WEIGHT_SIZE-1:0] Wgt_2_166,input [WEIGHT_SIZE-1:0] Wgt_2_167,input [WEIGHT_SIZE-1:0] Wgt_2_168,input [WEIGHT_SIZE-1:0] Wgt_2_169,input [WEIGHT_SIZE-1:0] Wgt_2_170,input [WEIGHT_SIZE-1:0] Wgt_2_171,input [WEIGHT_SIZE-1:0] Wgt_2_172,input [WEIGHT_SIZE-1:0] Wgt_2_173,input [WEIGHT_SIZE-1:0] Wgt_2_174,input [WEIGHT_SIZE-1:0] Wgt_2_175,input [WEIGHT_SIZE-1:0] Wgt_2_176,input [WEIGHT_SIZE-1:0] Wgt_2_177,input [WEIGHT_SIZE-1:0] Wgt_2_178,input [WEIGHT_SIZE-1:0] Wgt_2_179,input [WEIGHT_SIZE-1:0] Wgt_2_180,input [WEIGHT_SIZE-1:0] Wgt_2_181,input [WEIGHT_SIZE-1:0] Wgt_2_182,input [WEIGHT_SIZE-1:0] Wgt_2_183,input [WEIGHT_SIZE-1:0] Wgt_2_184,input [WEIGHT_SIZE-1:0] Wgt_2_185,input [WEIGHT_SIZE-1:0] Wgt_2_186,input [WEIGHT_SIZE-1:0] Wgt_2_187,input [WEIGHT_SIZE-1:0] Wgt_2_188,input [WEIGHT_SIZE-1:0] Wgt_2_189,input [WEIGHT_SIZE-1:0] Wgt_2_190,input [WEIGHT_SIZE-1:0] Wgt_2_191,input [WEIGHT_SIZE-1:0] Wgt_2_192,input [WEIGHT_SIZE-1:0] Wgt_2_193,input [WEIGHT_SIZE-1:0] Wgt_2_194,input [WEIGHT_SIZE-1:0] Wgt_2_195,input [WEIGHT_SIZE-1:0] Wgt_2_196,input [WEIGHT_SIZE-1:0] Wgt_2_197,input [WEIGHT_SIZE-1:0] Wgt_2_198,input [WEIGHT_SIZE-1:0] Wgt_2_199,input [WEIGHT_SIZE-1:0] Wgt_2_200,input [WEIGHT_SIZE-1:0] Wgt_2_201,input [WEIGHT_SIZE-1:0] Wgt_2_202,input [WEIGHT_SIZE-1:0] Wgt_2_203,input [WEIGHT_SIZE-1:0] Wgt_2_204,input [WEIGHT_SIZE-1:0] Wgt_2_205,input [WEIGHT_SIZE-1:0] Wgt_2_206,input [WEIGHT_SIZE-1:0] Wgt_2_207,input [WEIGHT_SIZE-1:0] Wgt_2_208,input [WEIGHT_SIZE-1:0] Wgt_2_209,input [WEIGHT_SIZE-1:0] Wgt_2_210,input [WEIGHT_SIZE-1:0] Wgt_2_211,input [WEIGHT_SIZE-1:0] Wgt_2_212,input [WEIGHT_SIZE-1:0] Wgt_2_213,input [WEIGHT_SIZE-1:0] Wgt_2_214,input [WEIGHT_SIZE-1:0] Wgt_2_215,input [WEIGHT_SIZE-1:0] Wgt_2_216,input [WEIGHT_SIZE-1:0] Wgt_2_217,input [WEIGHT_SIZE-1:0] Wgt_2_218,input [WEIGHT_SIZE-1:0] Wgt_2_219,input [WEIGHT_SIZE-1:0] Wgt_2_220,input [WEIGHT_SIZE-1:0] Wgt_2_221,input [WEIGHT_SIZE-1:0] Wgt_2_222,input [WEIGHT_SIZE-1:0] Wgt_2_223,input [WEIGHT_SIZE-1:0] Wgt_2_224,input [WEIGHT_SIZE-1:0] Wgt_2_225,input [WEIGHT_SIZE-1:0] Wgt_2_226,input [WEIGHT_SIZE-1:0] Wgt_2_227,input [WEIGHT_SIZE-1:0] Wgt_2_228,input [WEIGHT_SIZE-1:0] Wgt_2_229,input [WEIGHT_SIZE-1:0] Wgt_2_230,input [WEIGHT_SIZE-1:0] Wgt_2_231,input [WEIGHT_SIZE-1:0] Wgt_2_232,input [WEIGHT_SIZE-1:0] Wgt_2_233,input [WEIGHT_SIZE-1:0] Wgt_2_234,input [WEIGHT_SIZE-1:0] Wgt_2_235,input [WEIGHT_SIZE-1:0] Wgt_2_236,input [WEIGHT_SIZE-1:0] Wgt_2_237,input [WEIGHT_SIZE-1:0] Wgt_2_238,input [WEIGHT_SIZE-1:0] Wgt_2_239,input [WEIGHT_SIZE-1:0] Wgt_2_240,input [WEIGHT_SIZE-1:0] Wgt_2_241,input [WEIGHT_SIZE-1:0] Wgt_2_242,input [WEIGHT_SIZE-1:0] Wgt_2_243,input [WEIGHT_SIZE-1:0] Wgt_2_244,input [WEIGHT_SIZE-1:0] Wgt_2_245,input [WEIGHT_SIZE-1:0] Wgt_2_246,input [WEIGHT_SIZE-1:0] Wgt_2_247,input [WEIGHT_SIZE-1:0] Wgt_2_248,input [WEIGHT_SIZE-1:0] Wgt_2_249,input [WEIGHT_SIZE-1:0] Wgt_2_250,input [WEIGHT_SIZE-1:0] Wgt_2_251,input [WEIGHT_SIZE-1:0] Wgt_2_252,input [WEIGHT_SIZE-1:0] Wgt_2_253,input [WEIGHT_SIZE-1:0] Wgt_2_254,input [WEIGHT_SIZE-1:0] Wgt_2_255,input [WEIGHT_SIZE-1:0] Wgt_2_256,input [WEIGHT_SIZE-1:0] Wgt_2_257,input [WEIGHT_SIZE-1:0] Wgt_2_258,input [WEIGHT_SIZE-1:0] Wgt_2_259,input [WEIGHT_SIZE-1:0] Wgt_2_260,input [WEIGHT_SIZE-1:0] Wgt_2_261,input [WEIGHT_SIZE-1:0] Wgt_2_262,input [WEIGHT_SIZE-1:0] Wgt_2_263,input [WEIGHT_SIZE-1:0] Wgt_2_264,input [WEIGHT_SIZE-1:0] Wgt_2_265,input [WEIGHT_SIZE-1:0] Wgt_2_266,input [WEIGHT_SIZE-1:0] Wgt_2_267,input [WEIGHT_SIZE-1:0] Wgt_2_268,input [WEIGHT_SIZE-1:0] Wgt_2_269,input [WEIGHT_SIZE-1:0] Wgt_2_270,input [WEIGHT_SIZE-1:0] Wgt_2_271,input [WEIGHT_SIZE-1:0] Wgt_2_272,input [WEIGHT_SIZE-1:0] Wgt_2_273,input [WEIGHT_SIZE-1:0] Wgt_2_274,input [WEIGHT_SIZE-1:0] Wgt_2_275,input [WEIGHT_SIZE-1:0] Wgt_2_276,input [WEIGHT_SIZE-1:0] Wgt_2_277,input [WEIGHT_SIZE-1:0] Wgt_2_278,input [WEIGHT_SIZE-1:0] Wgt_2_279,input [WEIGHT_SIZE-1:0] Wgt_2_280,input [WEIGHT_SIZE-1:0] Wgt_2_281,input [WEIGHT_SIZE-1:0] Wgt_2_282,input [WEIGHT_SIZE-1:0] Wgt_2_283,input [WEIGHT_SIZE-1:0] Wgt_2_284,input [WEIGHT_SIZE-1:0] Wgt_2_285,input [WEIGHT_SIZE-1:0] Wgt_2_286,input [WEIGHT_SIZE-1:0] Wgt_2_287,input [WEIGHT_SIZE-1:0] Wgt_2_288,input [WEIGHT_SIZE-1:0] Wgt_2_289,input [WEIGHT_SIZE-1:0] Wgt_2_290,input [WEIGHT_SIZE-1:0] Wgt_2_291,input [WEIGHT_SIZE-1:0] Wgt_2_292,input [WEIGHT_SIZE-1:0] Wgt_2_293,input [WEIGHT_SIZE-1:0] Wgt_2_294,input [WEIGHT_SIZE-1:0] Wgt_2_295,input [WEIGHT_SIZE-1:0] Wgt_2_296,input [WEIGHT_SIZE-1:0] Wgt_2_297,input [WEIGHT_SIZE-1:0] Wgt_2_298,input [WEIGHT_SIZE-1:0] Wgt_2_299,input [WEIGHT_SIZE-1:0] Wgt_2_300,input [WEIGHT_SIZE-1:0] Wgt_2_301,input [WEIGHT_SIZE-1:0] Wgt_2_302,input [WEIGHT_SIZE-1:0] Wgt_2_303,input [WEIGHT_SIZE-1:0] Wgt_2_304,input [WEIGHT_SIZE-1:0] Wgt_2_305,input [WEIGHT_SIZE-1:0] Wgt_2_306,input [WEIGHT_SIZE-1:0] Wgt_2_307,input [WEIGHT_SIZE-1:0] Wgt_2_308,input [WEIGHT_SIZE-1:0] Wgt_2_309,input [WEIGHT_SIZE-1:0] Wgt_2_310,input [WEIGHT_SIZE-1:0] Wgt_2_311,input [WEIGHT_SIZE-1:0] Wgt_2_312,input [WEIGHT_SIZE-1:0] Wgt_2_313,input [WEIGHT_SIZE-1:0] Wgt_2_314,input [WEIGHT_SIZE-1:0] Wgt_2_315,input [WEIGHT_SIZE-1:0] Wgt_2_316,input [WEIGHT_SIZE-1:0] Wgt_2_317,input [WEIGHT_SIZE-1:0] Wgt_2_318,input [WEIGHT_SIZE-1:0] Wgt_2_319,input [WEIGHT_SIZE-1:0] Wgt_2_320,input [WEIGHT_SIZE-1:0] Wgt_2_321,input [WEIGHT_SIZE-1:0] Wgt_2_322,input [WEIGHT_SIZE-1:0] Wgt_2_323,input [WEIGHT_SIZE-1:0] Wgt_2_324,input [WEIGHT_SIZE-1:0] Wgt_2_325,input [WEIGHT_SIZE-1:0] Wgt_2_326,input [WEIGHT_SIZE-1:0] Wgt_2_327,input [WEIGHT_SIZE-1:0] Wgt_2_328,input [WEIGHT_SIZE-1:0] Wgt_2_329,input [WEIGHT_SIZE-1:0] Wgt_2_330,input [WEIGHT_SIZE-1:0] Wgt_2_331,input [WEIGHT_SIZE-1:0] Wgt_2_332,input [WEIGHT_SIZE-1:0] Wgt_2_333,input [WEIGHT_SIZE-1:0] Wgt_2_334,input [WEIGHT_SIZE-1:0] Wgt_2_335,input [WEIGHT_SIZE-1:0] Wgt_2_336,input [WEIGHT_SIZE-1:0] Wgt_2_337,input [WEIGHT_SIZE-1:0] Wgt_2_338,input [WEIGHT_SIZE-1:0] Wgt_2_339,input [WEIGHT_SIZE-1:0] Wgt_2_340,input [WEIGHT_SIZE-1:0] Wgt_2_341,input [WEIGHT_SIZE-1:0] Wgt_2_342,input [WEIGHT_SIZE-1:0] Wgt_2_343,input [WEIGHT_SIZE-1:0] Wgt_2_344,input [WEIGHT_SIZE-1:0] Wgt_2_345,input [WEIGHT_SIZE-1:0] Wgt_2_346,input [WEIGHT_SIZE-1:0] Wgt_2_347,input [WEIGHT_SIZE-1:0] Wgt_2_348,input [WEIGHT_SIZE-1:0] Wgt_2_349,input [WEIGHT_SIZE-1:0] Wgt_2_350,input [WEIGHT_SIZE-1:0] Wgt_2_351,input [WEIGHT_SIZE-1:0] Wgt_2_352,input [WEIGHT_SIZE-1:0] Wgt_2_353,input [WEIGHT_SIZE-1:0] Wgt_2_354,input [WEIGHT_SIZE-1:0] Wgt_2_355,input [WEIGHT_SIZE-1:0] Wgt_2_356,input [WEIGHT_SIZE-1:0] Wgt_2_357,input [WEIGHT_SIZE-1:0] Wgt_2_358,input [WEIGHT_SIZE-1:0] Wgt_2_359,input [WEIGHT_SIZE-1:0] Wgt_2_360,input [WEIGHT_SIZE-1:0] Wgt_2_361,input [WEIGHT_SIZE-1:0] Wgt_2_362,input [WEIGHT_SIZE-1:0] Wgt_2_363,input [WEIGHT_SIZE-1:0] Wgt_2_364,input [WEIGHT_SIZE-1:0] Wgt_2_365,input [WEIGHT_SIZE-1:0] Wgt_2_366,input [WEIGHT_SIZE-1:0] Wgt_2_367,input [WEIGHT_SIZE-1:0] Wgt_2_368,input [WEIGHT_SIZE-1:0] Wgt_2_369,input [WEIGHT_SIZE-1:0] Wgt_2_370,input [WEIGHT_SIZE-1:0] Wgt_2_371,input [WEIGHT_SIZE-1:0] Wgt_2_372,input [WEIGHT_SIZE-1:0] Wgt_2_373,input [WEIGHT_SIZE-1:0] Wgt_2_374,input [WEIGHT_SIZE-1:0] Wgt_2_375,input [WEIGHT_SIZE-1:0] Wgt_2_376,input [WEIGHT_SIZE-1:0] Wgt_2_377,input [WEIGHT_SIZE-1:0] Wgt_2_378,input [WEIGHT_SIZE-1:0] Wgt_2_379,input [WEIGHT_SIZE-1:0] Wgt_2_380,input [WEIGHT_SIZE-1:0] Wgt_2_381,input [WEIGHT_SIZE-1:0] Wgt_2_382,input [WEIGHT_SIZE-1:0] Wgt_2_383,input [WEIGHT_SIZE-1:0] Wgt_2_384,input [WEIGHT_SIZE-1:0] Wgt_2_385,input [WEIGHT_SIZE-1:0] Wgt_2_386,input [WEIGHT_SIZE-1:0] Wgt_2_387,input [WEIGHT_SIZE-1:0] Wgt_2_388,input [WEIGHT_SIZE-1:0] Wgt_2_389,input [WEIGHT_SIZE-1:0] Wgt_2_390,input [WEIGHT_SIZE-1:0] Wgt_2_391,input [WEIGHT_SIZE-1:0] Wgt_2_392,input [WEIGHT_SIZE-1:0] Wgt_2_393,input [WEIGHT_SIZE-1:0] Wgt_2_394,input [WEIGHT_SIZE-1:0] Wgt_2_395,input [WEIGHT_SIZE-1:0] Wgt_2_396,input [WEIGHT_SIZE-1:0] Wgt_2_397,input [WEIGHT_SIZE-1:0] Wgt_2_398,input [WEIGHT_SIZE-1:0] Wgt_2_399,input [WEIGHT_SIZE-1:0] Wgt_2_400,input [WEIGHT_SIZE-1:0] Wgt_2_401,input [WEIGHT_SIZE-1:0] Wgt_2_402,input [WEIGHT_SIZE-1:0] Wgt_2_403,input [WEIGHT_SIZE-1:0] Wgt_2_404,input [WEIGHT_SIZE-1:0] Wgt_2_405,input [WEIGHT_SIZE-1:0] Wgt_2_406,input [WEIGHT_SIZE-1:0] Wgt_2_407,input [WEIGHT_SIZE-1:0] Wgt_2_408,input [WEIGHT_SIZE-1:0] Wgt_2_409,input [WEIGHT_SIZE-1:0] Wgt_2_410,input [WEIGHT_SIZE-1:0] Wgt_2_411,input [WEIGHT_SIZE-1:0] Wgt_2_412,input [WEIGHT_SIZE-1:0] Wgt_2_413,input [WEIGHT_SIZE-1:0] Wgt_2_414,input [WEIGHT_SIZE-1:0] Wgt_2_415,input [WEIGHT_SIZE-1:0] Wgt_2_416,input [WEIGHT_SIZE-1:0] Wgt_2_417,input [WEIGHT_SIZE-1:0] Wgt_2_418,input [WEIGHT_SIZE-1:0] Wgt_2_419,input [WEIGHT_SIZE-1:0] Wgt_2_420,input [WEIGHT_SIZE-1:0] Wgt_2_421,input [WEIGHT_SIZE-1:0] Wgt_2_422,input [WEIGHT_SIZE-1:0] Wgt_2_423,input [WEIGHT_SIZE-1:0] Wgt_2_424,input [WEIGHT_SIZE-1:0] Wgt_2_425,input [WEIGHT_SIZE-1:0] Wgt_2_426,input [WEIGHT_SIZE-1:0] Wgt_2_427,input [WEIGHT_SIZE-1:0] Wgt_2_428,input [WEIGHT_SIZE-1:0] Wgt_2_429,input [WEIGHT_SIZE-1:0] Wgt_2_430,input [WEIGHT_SIZE-1:0] Wgt_2_431,input [WEIGHT_SIZE-1:0] Wgt_2_432,input [WEIGHT_SIZE-1:0] Wgt_2_433,input [WEIGHT_SIZE-1:0] Wgt_2_434,input [WEIGHT_SIZE-1:0] Wgt_2_435,input [WEIGHT_SIZE-1:0] Wgt_2_436,input [WEIGHT_SIZE-1:0] Wgt_2_437,input [WEIGHT_SIZE-1:0] Wgt_2_438,input [WEIGHT_SIZE-1:0] Wgt_2_439,input [WEIGHT_SIZE-1:0] Wgt_2_440,input [WEIGHT_SIZE-1:0] Wgt_2_441,input [WEIGHT_SIZE-1:0] Wgt_2_442,input [WEIGHT_SIZE-1:0] Wgt_2_443,input [WEIGHT_SIZE-1:0] Wgt_2_444,input [WEIGHT_SIZE-1:0] Wgt_2_445,input [WEIGHT_SIZE-1:0] Wgt_2_446,input [WEIGHT_SIZE-1:0] Wgt_2_447,input [WEIGHT_SIZE-1:0] Wgt_2_448,input [WEIGHT_SIZE-1:0] Wgt_2_449,input [WEIGHT_SIZE-1:0] Wgt_2_450,input [WEIGHT_SIZE-1:0] Wgt_2_451,input [WEIGHT_SIZE-1:0] Wgt_2_452,input [WEIGHT_SIZE-1:0] Wgt_2_453,input [WEIGHT_SIZE-1:0] Wgt_2_454,input [WEIGHT_SIZE-1:0] Wgt_2_455,input [WEIGHT_SIZE-1:0] Wgt_2_456,input [WEIGHT_SIZE-1:0] Wgt_2_457,input [WEIGHT_SIZE-1:0] Wgt_2_458,input [WEIGHT_SIZE-1:0] Wgt_2_459,input [WEIGHT_SIZE-1:0] Wgt_2_460,input [WEIGHT_SIZE-1:0] Wgt_2_461,input [WEIGHT_SIZE-1:0] Wgt_2_462,input [WEIGHT_SIZE-1:0] Wgt_2_463,input [WEIGHT_SIZE-1:0] Wgt_2_464,input [WEIGHT_SIZE-1:0] Wgt_2_465,input [WEIGHT_SIZE-1:0] Wgt_2_466,input [WEIGHT_SIZE-1:0] Wgt_2_467,input [WEIGHT_SIZE-1:0] Wgt_2_468,input [WEIGHT_SIZE-1:0] Wgt_2_469,input [WEIGHT_SIZE-1:0] Wgt_2_470,input [WEIGHT_SIZE-1:0] Wgt_2_471,input [WEIGHT_SIZE-1:0] Wgt_2_472,input [WEIGHT_SIZE-1:0] Wgt_2_473,input [WEIGHT_SIZE-1:0] Wgt_2_474,input [WEIGHT_SIZE-1:0] Wgt_2_475,input [WEIGHT_SIZE-1:0] Wgt_2_476,input [WEIGHT_SIZE-1:0] Wgt_2_477,input [WEIGHT_SIZE-1:0] Wgt_2_478,input [WEIGHT_SIZE-1:0] Wgt_2_479,input [WEIGHT_SIZE-1:0] Wgt_2_480,input [WEIGHT_SIZE-1:0] Wgt_2_481,input [WEIGHT_SIZE-1:0] Wgt_2_482,input [WEIGHT_SIZE-1:0] Wgt_2_483,input [WEIGHT_SIZE-1:0] Wgt_2_484,input [WEIGHT_SIZE-1:0] Wgt_2_485,input [WEIGHT_SIZE-1:0] Wgt_2_486,input [WEIGHT_SIZE-1:0] Wgt_2_487,input [WEIGHT_SIZE-1:0] Wgt_2_488,input [WEIGHT_SIZE-1:0] Wgt_2_489,input [WEIGHT_SIZE-1:0] Wgt_2_490,input [WEIGHT_SIZE-1:0] Wgt_2_491,input [WEIGHT_SIZE-1:0] Wgt_2_492,input [WEIGHT_SIZE-1:0] Wgt_2_493,input [WEIGHT_SIZE-1:0] Wgt_2_494,input [WEIGHT_SIZE-1:0] Wgt_2_495,input [WEIGHT_SIZE-1:0] Wgt_2_496,input [WEIGHT_SIZE-1:0] Wgt_2_497,input [WEIGHT_SIZE-1:0] Wgt_2_498,input [WEIGHT_SIZE-1:0] Wgt_2_499,input [WEIGHT_SIZE-1:0] Wgt_2_500,input [WEIGHT_SIZE-1:0] Wgt_2_501,input [WEIGHT_SIZE-1:0] Wgt_2_502,input [WEIGHT_SIZE-1:0] Wgt_2_503,input [WEIGHT_SIZE-1:0] Wgt_2_504,input [WEIGHT_SIZE-1:0] Wgt_2_505,input [WEIGHT_SIZE-1:0] Wgt_2_506,input [WEIGHT_SIZE-1:0] Wgt_2_507,input [WEIGHT_SIZE-1:0] Wgt_2_508,input [WEIGHT_SIZE-1:0] Wgt_2_509,input [WEIGHT_SIZE-1:0] Wgt_2_510,input [WEIGHT_SIZE-1:0] Wgt_2_511,input [WEIGHT_SIZE-1:0] Wgt_2_512,input [WEIGHT_SIZE-1:0] Wgt_2_513,input [WEIGHT_SIZE-1:0] Wgt_2_514,input [WEIGHT_SIZE-1:0] Wgt_2_515,input [WEIGHT_SIZE-1:0] Wgt_2_516,input [WEIGHT_SIZE-1:0] Wgt_2_517,input [WEIGHT_SIZE-1:0] Wgt_2_518,input [WEIGHT_SIZE-1:0] Wgt_2_519,input [WEIGHT_SIZE-1:0] Wgt_2_520,input [WEIGHT_SIZE-1:0] Wgt_2_521,input [WEIGHT_SIZE-1:0] Wgt_2_522,input [WEIGHT_SIZE-1:0] Wgt_2_523,input [WEIGHT_SIZE-1:0] Wgt_2_524,input [WEIGHT_SIZE-1:0] Wgt_2_525,input [WEIGHT_SIZE-1:0] Wgt_2_526,input [WEIGHT_SIZE-1:0] Wgt_2_527,input [WEIGHT_SIZE-1:0] Wgt_2_528,input [WEIGHT_SIZE-1:0] Wgt_2_529,input [WEIGHT_SIZE-1:0] Wgt_2_530,input [WEIGHT_SIZE-1:0] Wgt_2_531,input [WEIGHT_SIZE-1:0] Wgt_2_532,input [WEIGHT_SIZE-1:0] Wgt_2_533,input [WEIGHT_SIZE-1:0] Wgt_2_534,input [WEIGHT_SIZE-1:0] Wgt_2_535,input [WEIGHT_SIZE-1:0] Wgt_2_536,input [WEIGHT_SIZE-1:0] Wgt_2_537,input [WEIGHT_SIZE-1:0] Wgt_2_538,input [WEIGHT_SIZE-1:0] Wgt_2_539,input [WEIGHT_SIZE-1:0] Wgt_2_540,input [WEIGHT_SIZE-1:0] Wgt_2_541,input [WEIGHT_SIZE-1:0] Wgt_2_542,input [WEIGHT_SIZE-1:0] Wgt_2_543,input [WEIGHT_SIZE-1:0] Wgt_2_544,input [WEIGHT_SIZE-1:0] Wgt_2_545,input [WEIGHT_SIZE-1:0] Wgt_2_546,input [WEIGHT_SIZE-1:0] Wgt_2_547,input [WEIGHT_SIZE-1:0] Wgt_2_548,input [WEIGHT_SIZE-1:0] Wgt_2_549,input [WEIGHT_SIZE-1:0] Wgt_2_550,input [WEIGHT_SIZE-1:0] Wgt_2_551,input [WEIGHT_SIZE-1:0] Wgt_2_552,input [WEIGHT_SIZE-1:0] Wgt_2_553,input [WEIGHT_SIZE-1:0] Wgt_2_554,input [WEIGHT_SIZE-1:0] Wgt_2_555,input [WEIGHT_SIZE-1:0] Wgt_2_556,input [WEIGHT_SIZE-1:0] Wgt_2_557,input [WEIGHT_SIZE-1:0] Wgt_2_558,input [WEIGHT_SIZE-1:0] Wgt_2_559,input [WEIGHT_SIZE-1:0] Wgt_2_560,input [WEIGHT_SIZE-1:0] Wgt_2_561,input [WEIGHT_SIZE-1:0] Wgt_2_562,input [WEIGHT_SIZE-1:0] Wgt_2_563,input [WEIGHT_SIZE-1:0] Wgt_2_564,input [WEIGHT_SIZE-1:0] Wgt_2_565,input [WEIGHT_SIZE-1:0] Wgt_2_566,input [WEIGHT_SIZE-1:0] Wgt_2_567,input [WEIGHT_SIZE-1:0] Wgt_2_568,input [WEIGHT_SIZE-1:0] Wgt_2_569,input [WEIGHT_SIZE-1:0] Wgt_2_570,input [WEIGHT_SIZE-1:0] Wgt_2_571,input [WEIGHT_SIZE-1:0] Wgt_2_572,input [WEIGHT_SIZE-1:0] Wgt_2_573,input [WEIGHT_SIZE-1:0] Wgt_2_574,input [WEIGHT_SIZE-1:0] Wgt_2_575,input [WEIGHT_SIZE-1:0] Wgt_2_576,input [WEIGHT_SIZE-1:0] Wgt_2_577,input [WEIGHT_SIZE-1:0] Wgt_2_578,input [WEIGHT_SIZE-1:0] Wgt_2_579,input [WEIGHT_SIZE-1:0] Wgt_2_580,input [WEIGHT_SIZE-1:0] Wgt_2_581,input [WEIGHT_SIZE-1:0] Wgt_2_582,input [WEIGHT_SIZE-1:0] Wgt_2_583,input [WEIGHT_SIZE-1:0] Wgt_2_584,input [WEIGHT_SIZE-1:0] Wgt_2_585,input [WEIGHT_SIZE-1:0] Wgt_2_586,input [WEIGHT_SIZE-1:0] Wgt_2_587,input [WEIGHT_SIZE-1:0] Wgt_2_588,input [WEIGHT_SIZE-1:0] Wgt_2_589,input [WEIGHT_SIZE-1:0] Wgt_2_590,input [WEIGHT_SIZE-1:0] Wgt_2_591,input [WEIGHT_SIZE-1:0] Wgt_2_592,input [WEIGHT_SIZE-1:0] Wgt_2_593,input [WEIGHT_SIZE-1:0] Wgt_2_594,input [WEIGHT_SIZE-1:0] Wgt_2_595,input [WEIGHT_SIZE-1:0] Wgt_2_596,input [WEIGHT_SIZE-1:0] Wgt_2_597,input [WEIGHT_SIZE-1:0] Wgt_2_598,input [WEIGHT_SIZE-1:0] Wgt_2_599,input [WEIGHT_SIZE-1:0] Wgt_2_600,input [WEIGHT_SIZE-1:0] Wgt_2_601,input [WEIGHT_SIZE-1:0] Wgt_2_602,input [WEIGHT_SIZE-1:0] Wgt_2_603,input [WEIGHT_SIZE-1:0] Wgt_2_604,input [WEIGHT_SIZE-1:0] Wgt_2_605,input [WEIGHT_SIZE-1:0] Wgt_2_606,input [WEIGHT_SIZE-1:0] Wgt_2_607,input [WEIGHT_SIZE-1:0] Wgt_2_608,input [WEIGHT_SIZE-1:0] Wgt_2_609,input [WEIGHT_SIZE-1:0] Wgt_2_610,input [WEIGHT_SIZE-1:0] Wgt_2_611,input [WEIGHT_SIZE-1:0] Wgt_2_612,input [WEIGHT_SIZE-1:0] Wgt_2_613,input [WEIGHT_SIZE-1:0] Wgt_2_614,input [WEIGHT_SIZE-1:0] Wgt_2_615,input [WEIGHT_SIZE-1:0] Wgt_2_616,input [WEIGHT_SIZE-1:0] Wgt_2_617,input [WEIGHT_SIZE-1:0] Wgt_2_618,input [WEIGHT_SIZE-1:0] Wgt_2_619,input [WEIGHT_SIZE-1:0] Wgt_2_620,input [WEIGHT_SIZE-1:0] Wgt_2_621,input [WEIGHT_SIZE-1:0] Wgt_2_622,input [WEIGHT_SIZE-1:0] Wgt_2_623,input [WEIGHT_SIZE-1:0] Wgt_2_624,input [WEIGHT_SIZE-1:0] Wgt_2_625,input [WEIGHT_SIZE-1:0] Wgt_2_626,input [WEIGHT_SIZE-1:0] Wgt_2_627,input [WEIGHT_SIZE-1:0] Wgt_2_628,input [WEIGHT_SIZE-1:0] Wgt_2_629,input [WEIGHT_SIZE-1:0] Wgt_2_630,input [WEIGHT_SIZE-1:0] Wgt_2_631,input [WEIGHT_SIZE-1:0] Wgt_2_632,input [WEIGHT_SIZE-1:0] Wgt_2_633,input [WEIGHT_SIZE-1:0] Wgt_2_634,input [WEIGHT_SIZE-1:0] Wgt_2_635,input [WEIGHT_SIZE-1:0] Wgt_2_636,input [WEIGHT_SIZE-1:0] Wgt_2_637,input [WEIGHT_SIZE-1:0] Wgt_2_638,input [WEIGHT_SIZE-1:0] Wgt_2_639,input [WEIGHT_SIZE-1:0] Wgt_2_640,input [WEIGHT_SIZE-1:0] Wgt_2_641,input [WEIGHT_SIZE-1:0] Wgt_2_642,input [WEIGHT_SIZE-1:0] Wgt_2_643,input [WEIGHT_SIZE-1:0] Wgt_2_644,input [WEIGHT_SIZE-1:0] Wgt_2_645,input [WEIGHT_SIZE-1:0] Wgt_2_646,input [WEIGHT_SIZE-1:0] Wgt_2_647,input [WEIGHT_SIZE-1:0] Wgt_2_648,input [WEIGHT_SIZE-1:0] Wgt_2_649,input [WEIGHT_SIZE-1:0] Wgt_2_650,input [WEIGHT_SIZE-1:0] Wgt_2_651,input [WEIGHT_SIZE-1:0] Wgt_2_652,input [WEIGHT_SIZE-1:0] Wgt_2_653,input [WEIGHT_SIZE-1:0] Wgt_2_654,input [WEIGHT_SIZE-1:0] Wgt_2_655,input [WEIGHT_SIZE-1:0] Wgt_2_656,input [WEIGHT_SIZE-1:0] Wgt_2_657,input [WEIGHT_SIZE-1:0] Wgt_2_658,input [WEIGHT_SIZE-1:0] Wgt_2_659,input [WEIGHT_SIZE-1:0] Wgt_2_660,input [WEIGHT_SIZE-1:0] Wgt_2_661,input [WEIGHT_SIZE-1:0] Wgt_2_662,input [WEIGHT_SIZE-1:0] Wgt_2_663,input [WEIGHT_SIZE-1:0] Wgt_2_664,input [WEIGHT_SIZE-1:0] Wgt_2_665,input [WEIGHT_SIZE-1:0] Wgt_2_666,input [WEIGHT_SIZE-1:0] Wgt_2_667,input [WEIGHT_SIZE-1:0] Wgt_2_668,input [WEIGHT_SIZE-1:0] Wgt_2_669,input [WEIGHT_SIZE-1:0] Wgt_2_670,input [WEIGHT_SIZE-1:0] Wgt_2_671,input [WEIGHT_SIZE-1:0] Wgt_2_672,input [WEIGHT_SIZE-1:0] Wgt_2_673,input [WEIGHT_SIZE-1:0] Wgt_2_674,input [WEIGHT_SIZE-1:0] Wgt_2_675,input [WEIGHT_SIZE-1:0] Wgt_2_676,input [WEIGHT_SIZE-1:0] Wgt_2_677,input [WEIGHT_SIZE-1:0] Wgt_2_678,input [WEIGHT_SIZE-1:0] Wgt_2_679,input [WEIGHT_SIZE-1:0] Wgt_2_680,input [WEIGHT_SIZE-1:0] Wgt_2_681,input [WEIGHT_SIZE-1:0] Wgt_2_682,input [WEIGHT_SIZE-1:0] Wgt_2_683,input [WEIGHT_SIZE-1:0] Wgt_2_684,input [WEIGHT_SIZE-1:0] Wgt_2_685,input [WEIGHT_SIZE-1:0] Wgt_2_686,input [WEIGHT_SIZE-1:0] Wgt_2_687,input [WEIGHT_SIZE-1:0] Wgt_2_688,input [WEIGHT_SIZE-1:0] Wgt_2_689,input [WEIGHT_SIZE-1:0] Wgt_2_690,input [WEIGHT_SIZE-1:0] Wgt_2_691,input [WEIGHT_SIZE-1:0] Wgt_2_692,input [WEIGHT_SIZE-1:0] Wgt_2_693,input [WEIGHT_SIZE-1:0] Wgt_2_694,input [WEIGHT_SIZE-1:0] Wgt_2_695,input [WEIGHT_SIZE-1:0] Wgt_2_696,input [WEIGHT_SIZE-1:0] Wgt_2_697,input [WEIGHT_SIZE-1:0] Wgt_2_698,input [WEIGHT_SIZE-1:0] Wgt_2_699,input [WEIGHT_SIZE-1:0] Wgt_2_700,input [WEIGHT_SIZE-1:0] Wgt_2_701,input [WEIGHT_SIZE-1:0] Wgt_2_702,input [WEIGHT_SIZE-1:0] Wgt_2_703,input [WEIGHT_SIZE-1:0] Wgt_2_704,input [WEIGHT_SIZE-1:0] Wgt_2_705,input [WEIGHT_SIZE-1:0] Wgt_2_706,input [WEIGHT_SIZE-1:0] Wgt_2_707,input [WEIGHT_SIZE-1:0] Wgt_2_708,input [WEIGHT_SIZE-1:0] Wgt_2_709,input [WEIGHT_SIZE-1:0] Wgt_2_710,input [WEIGHT_SIZE-1:0] Wgt_2_711,input [WEIGHT_SIZE-1:0] Wgt_2_712,input [WEIGHT_SIZE-1:0] Wgt_2_713,input [WEIGHT_SIZE-1:0] Wgt_2_714,input [WEIGHT_SIZE-1:0] Wgt_2_715,input [WEIGHT_SIZE-1:0] Wgt_2_716,input [WEIGHT_SIZE-1:0] Wgt_2_717,input [WEIGHT_SIZE-1:0] Wgt_2_718,input [WEIGHT_SIZE-1:0] Wgt_2_719,input [WEIGHT_SIZE-1:0] Wgt_2_720,input [WEIGHT_SIZE-1:0] Wgt_2_721,input [WEIGHT_SIZE-1:0] Wgt_2_722,input [WEIGHT_SIZE-1:0] Wgt_2_723,input [WEIGHT_SIZE-1:0] Wgt_2_724,input [WEIGHT_SIZE-1:0] Wgt_2_725,input [WEIGHT_SIZE-1:0] Wgt_2_726,input [WEIGHT_SIZE-1:0] Wgt_2_727,input [WEIGHT_SIZE-1:0] Wgt_2_728,input [WEIGHT_SIZE-1:0] Wgt_2_729,input [WEIGHT_SIZE-1:0] Wgt_2_730,input [WEIGHT_SIZE-1:0] Wgt_2_731,input [WEIGHT_SIZE-1:0] Wgt_2_732,input [WEIGHT_SIZE-1:0] Wgt_2_733,input [WEIGHT_SIZE-1:0] Wgt_2_734,input [WEIGHT_SIZE-1:0] Wgt_2_735,input [WEIGHT_SIZE-1:0] Wgt_2_736,input [WEIGHT_SIZE-1:0] Wgt_2_737,input [WEIGHT_SIZE-1:0] Wgt_2_738,input [WEIGHT_SIZE-1:0] Wgt_2_739,input [WEIGHT_SIZE-1:0] Wgt_2_740,input [WEIGHT_SIZE-1:0] Wgt_2_741,input [WEIGHT_SIZE-1:0] Wgt_2_742,input [WEIGHT_SIZE-1:0] Wgt_2_743,input [WEIGHT_SIZE-1:0] Wgt_2_744,input [WEIGHT_SIZE-1:0] Wgt_2_745,input [WEIGHT_SIZE-1:0] Wgt_2_746,input [WEIGHT_SIZE-1:0] Wgt_2_747,input [WEIGHT_SIZE-1:0] Wgt_2_748,input [WEIGHT_SIZE-1:0] Wgt_2_749,input [WEIGHT_SIZE-1:0] Wgt_2_750,input [WEIGHT_SIZE-1:0] Wgt_2_751,input [WEIGHT_SIZE-1:0] Wgt_2_752,input [WEIGHT_SIZE-1:0] Wgt_2_753,input [WEIGHT_SIZE-1:0] Wgt_2_754,input [WEIGHT_SIZE-1:0] Wgt_2_755,input [WEIGHT_SIZE-1:0] Wgt_2_756,input [WEIGHT_SIZE-1:0] Wgt_2_757,input [WEIGHT_SIZE-1:0] Wgt_2_758,input [WEIGHT_SIZE-1:0] Wgt_2_759,input [WEIGHT_SIZE-1:0] Wgt_2_760,input [WEIGHT_SIZE-1:0] Wgt_2_761,input [WEIGHT_SIZE-1:0] Wgt_2_762,input [WEIGHT_SIZE-1:0] Wgt_2_763,input [WEIGHT_SIZE-1:0] Wgt_2_764,input [WEIGHT_SIZE-1:0] Wgt_2_765,input [WEIGHT_SIZE-1:0] Wgt_2_766,input [WEIGHT_SIZE-1:0] Wgt_2_767,input [WEIGHT_SIZE-1:0] Wgt_2_768,input [WEIGHT_SIZE-1:0] Wgt_2_769,input [WEIGHT_SIZE-1:0] Wgt_2_770,input [WEIGHT_SIZE-1:0] Wgt_2_771,input [WEIGHT_SIZE-1:0] Wgt_2_772,input [WEIGHT_SIZE-1:0] Wgt_2_773,input [WEIGHT_SIZE-1:0] Wgt_2_774,input [WEIGHT_SIZE-1:0] Wgt_2_775,input [WEIGHT_SIZE-1:0] Wgt_2_776,input [WEIGHT_SIZE-1:0] Wgt_2_777,input [WEIGHT_SIZE-1:0] Wgt_2_778,input [WEIGHT_SIZE-1:0] Wgt_2_779,input [WEIGHT_SIZE-1:0] Wgt_2_780,input [WEIGHT_SIZE-1:0] Wgt_2_781,input [WEIGHT_SIZE-1:0] Wgt_2_782,input [WEIGHT_SIZE-1:0] Wgt_2_783,input [WEIGHT_SIZE-1:0] Wgt_2_784,input [WEIGHT_SIZE-1:0] Wgt_3_0,input [WEIGHT_SIZE-1:0] Wgt_3_1,input [WEIGHT_SIZE-1:0] Wgt_3_2,input [WEIGHT_SIZE-1:0] Wgt_3_3,input [WEIGHT_SIZE-1:0] Wgt_3_4,input [WEIGHT_SIZE-1:0] Wgt_3_5,input [WEIGHT_SIZE-1:0] Wgt_3_6,input [WEIGHT_SIZE-1:0] Wgt_3_7,input [WEIGHT_SIZE-1:0] Wgt_3_8,input [WEIGHT_SIZE-1:0] Wgt_3_9,input [WEIGHT_SIZE-1:0] Wgt_3_10,input [WEIGHT_SIZE-1:0] Wgt_3_11,input [WEIGHT_SIZE-1:0] Wgt_3_12,input [WEIGHT_SIZE-1:0] Wgt_3_13,input [WEIGHT_SIZE-1:0] Wgt_3_14,input [WEIGHT_SIZE-1:0] Wgt_3_15,input [WEIGHT_SIZE-1:0] Wgt_3_16,input [WEIGHT_SIZE-1:0] Wgt_3_17,input [WEIGHT_SIZE-1:0] Wgt_3_18,input [WEIGHT_SIZE-1:0] Wgt_3_19,input [WEIGHT_SIZE-1:0] Wgt_3_20,input [WEIGHT_SIZE-1:0] Wgt_3_21,input [WEIGHT_SIZE-1:0] Wgt_3_22,input [WEIGHT_SIZE-1:0] Wgt_3_23,input [WEIGHT_SIZE-1:0] Wgt_3_24,input [WEIGHT_SIZE-1:0] Wgt_3_25,input [WEIGHT_SIZE-1:0] Wgt_3_26,input [WEIGHT_SIZE-1:0] Wgt_3_27,input [WEIGHT_SIZE-1:0] Wgt_3_28,input [WEIGHT_SIZE-1:0] Wgt_3_29,input [WEIGHT_SIZE-1:0] Wgt_3_30,input [WEIGHT_SIZE-1:0] Wgt_3_31,input [WEIGHT_SIZE-1:0] Wgt_3_32,input [WEIGHT_SIZE-1:0] Wgt_3_33,input [WEIGHT_SIZE-1:0] Wgt_3_34,input [WEIGHT_SIZE-1:0] Wgt_3_35,input [WEIGHT_SIZE-1:0] Wgt_3_36,input [WEIGHT_SIZE-1:0] Wgt_3_37,input [WEIGHT_SIZE-1:0] Wgt_3_38,input [WEIGHT_SIZE-1:0] Wgt_3_39,input [WEIGHT_SIZE-1:0] Wgt_3_40,input [WEIGHT_SIZE-1:0] Wgt_3_41,input [WEIGHT_SIZE-1:0] Wgt_3_42,input [WEIGHT_SIZE-1:0] Wgt_3_43,input [WEIGHT_SIZE-1:0] Wgt_3_44,input [WEIGHT_SIZE-1:0] Wgt_3_45,input [WEIGHT_SIZE-1:0] Wgt_3_46,input [WEIGHT_SIZE-1:0] Wgt_3_47,input [WEIGHT_SIZE-1:0] Wgt_3_48,input [WEIGHT_SIZE-1:0] Wgt_3_49,input [WEIGHT_SIZE-1:0] Wgt_3_50,input [WEIGHT_SIZE-1:0] Wgt_3_51,input [WEIGHT_SIZE-1:0] Wgt_3_52,input [WEIGHT_SIZE-1:0] Wgt_3_53,input [WEIGHT_SIZE-1:0] Wgt_3_54,input [WEIGHT_SIZE-1:0] Wgt_3_55,input [WEIGHT_SIZE-1:0] Wgt_3_56,input [WEIGHT_SIZE-1:0] Wgt_3_57,input [WEIGHT_SIZE-1:0] Wgt_3_58,input [WEIGHT_SIZE-1:0] Wgt_3_59,input [WEIGHT_SIZE-1:0] Wgt_3_60,input [WEIGHT_SIZE-1:0] Wgt_3_61,input [WEIGHT_SIZE-1:0] Wgt_3_62,input [WEIGHT_SIZE-1:0] Wgt_3_63,input [WEIGHT_SIZE-1:0] Wgt_3_64,input [WEIGHT_SIZE-1:0] Wgt_3_65,input [WEIGHT_SIZE-1:0] Wgt_3_66,input [WEIGHT_SIZE-1:0] Wgt_3_67,input [WEIGHT_SIZE-1:0] Wgt_3_68,input [WEIGHT_SIZE-1:0] Wgt_3_69,input [WEIGHT_SIZE-1:0] Wgt_3_70,input [WEIGHT_SIZE-1:0] Wgt_3_71,input [WEIGHT_SIZE-1:0] Wgt_3_72,input [WEIGHT_SIZE-1:0] Wgt_3_73,input [WEIGHT_SIZE-1:0] Wgt_3_74,input [WEIGHT_SIZE-1:0] Wgt_3_75,input [WEIGHT_SIZE-1:0] Wgt_3_76,input [WEIGHT_SIZE-1:0] Wgt_3_77,input [WEIGHT_SIZE-1:0] Wgt_3_78,input [WEIGHT_SIZE-1:0] Wgt_3_79,input [WEIGHT_SIZE-1:0] Wgt_3_80,input [WEIGHT_SIZE-1:0] Wgt_3_81,input [WEIGHT_SIZE-1:0] Wgt_3_82,input [WEIGHT_SIZE-1:0] Wgt_3_83,input [WEIGHT_SIZE-1:0] Wgt_3_84,input [WEIGHT_SIZE-1:0] Wgt_3_85,input [WEIGHT_SIZE-1:0] Wgt_3_86,input [WEIGHT_SIZE-1:0] Wgt_3_87,input [WEIGHT_SIZE-1:0] Wgt_3_88,input [WEIGHT_SIZE-1:0] Wgt_3_89,input [WEIGHT_SIZE-1:0] Wgt_3_90,input [WEIGHT_SIZE-1:0] Wgt_3_91,input [WEIGHT_SIZE-1:0] Wgt_3_92,input [WEIGHT_SIZE-1:0] Wgt_3_93,input [WEIGHT_SIZE-1:0] Wgt_3_94,input [WEIGHT_SIZE-1:0] Wgt_3_95,input [WEIGHT_SIZE-1:0] Wgt_3_96,input [WEIGHT_SIZE-1:0] Wgt_3_97,input [WEIGHT_SIZE-1:0] Wgt_3_98,input [WEIGHT_SIZE-1:0] Wgt_3_99,input [WEIGHT_SIZE-1:0] Wgt_3_100,input [WEIGHT_SIZE-1:0] Wgt_3_101,input [WEIGHT_SIZE-1:0] Wgt_3_102,input [WEIGHT_SIZE-1:0] Wgt_3_103,input [WEIGHT_SIZE-1:0] Wgt_3_104,input [WEIGHT_SIZE-1:0] Wgt_3_105,input [WEIGHT_SIZE-1:0] Wgt_3_106,input [WEIGHT_SIZE-1:0] Wgt_3_107,input [WEIGHT_SIZE-1:0] Wgt_3_108,input [WEIGHT_SIZE-1:0] Wgt_3_109,input [WEIGHT_SIZE-1:0] Wgt_3_110,input [WEIGHT_SIZE-1:0] Wgt_3_111,input [WEIGHT_SIZE-1:0] Wgt_3_112,input [WEIGHT_SIZE-1:0] Wgt_3_113,input [WEIGHT_SIZE-1:0] Wgt_3_114,input [WEIGHT_SIZE-1:0] Wgt_3_115,input [WEIGHT_SIZE-1:0] Wgt_3_116,input [WEIGHT_SIZE-1:0] Wgt_3_117,input [WEIGHT_SIZE-1:0] Wgt_3_118,input [WEIGHT_SIZE-1:0] Wgt_3_119,input [WEIGHT_SIZE-1:0] Wgt_3_120,input [WEIGHT_SIZE-1:0] Wgt_3_121,input [WEIGHT_SIZE-1:0] Wgt_3_122,input [WEIGHT_SIZE-1:0] Wgt_3_123,input [WEIGHT_SIZE-1:0] Wgt_3_124,input [WEIGHT_SIZE-1:0] Wgt_3_125,input [WEIGHT_SIZE-1:0] Wgt_3_126,input [WEIGHT_SIZE-1:0] Wgt_3_127,input [WEIGHT_SIZE-1:0] Wgt_3_128,input [WEIGHT_SIZE-1:0] Wgt_3_129,input [WEIGHT_SIZE-1:0] Wgt_3_130,input [WEIGHT_SIZE-1:0] Wgt_3_131,input [WEIGHT_SIZE-1:0] Wgt_3_132,input [WEIGHT_SIZE-1:0] Wgt_3_133,input [WEIGHT_SIZE-1:0] Wgt_3_134,input [WEIGHT_SIZE-1:0] Wgt_3_135,input [WEIGHT_SIZE-1:0] Wgt_3_136,input [WEIGHT_SIZE-1:0] Wgt_3_137,input [WEIGHT_SIZE-1:0] Wgt_3_138,input [WEIGHT_SIZE-1:0] Wgt_3_139,input [WEIGHT_SIZE-1:0] Wgt_3_140,input [WEIGHT_SIZE-1:0] Wgt_3_141,input [WEIGHT_SIZE-1:0] Wgt_3_142,input [WEIGHT_SIZE-1:0] Wgt_3_143,input [WEIGHT_SIZE-1:0] Wgt_3_144,input [WEIGHT_SIZE-1:0] Wgt_3_145,input [WEIGHT_SIZE-1:0] Wgt_3_146,input [WEIGHT_SIZE-1:0] Wgt_3_147,input [WEIGHT_SIZE-1:0] Wgt_3_148,input [WEIGHT_SIZE-1:0] Wgt_3_149,input [WEIGHT_SIZE-1:0] Wgt_3_150,input [WEIGHT_SIZE-1:0] Wgt_3_151,input [WEIGHT_SIZE-1:0] Wgt_3_152,input [WEIGHT_SIZE-1:0] Wgt_3_153,input [WEIGHT_SIZE-1:0] Wgt_3_154,input [WEIGHT_SIZE-1:0] Wgt_3_155,input [WEIGHT_SIZE-1:0] Wgt_3_156,input [WEIGHT_SIZE-1:0] Wgt_3_157,input [WEIGHT_SIZE-1:0] Wgt_3_158,input [WEIGHT_SIZE-1:0] Wgt_3_159,input [WEIGHT_SIZE-1:0] Wgt_3_160,input [WEIGHT_SIZE-1:0] Wgt_3_161,input [WEIGHT_SIZE-1:0] Wgt_3_162,input [WEIGHT_SIZE-1:0] Wgt_3_163,input [WEIGHT_SIZE-1:0] Wgt_3_164,input [WEIGHT_SIZE-1:0] Wgt_3_165,input [WEIGHT_SIZE-1:0] Wgt_3_166,input [WEIGHT_SIZE-1:0] Wgt_3_167,input [WEIGHT_SIZE-1:0] Wgt_3_168,input [WEIGHT_SIZE-1:0] Wgt_3_169,input [WEIGHT_SIZE-1:0] Wgt_3_170,input [WEIGHT_SIZE-1:0] Wgt_3_171,input [WEIGHT_SIZE-1:0] Wgt_3_172,input [WEIGHT_SIZE-1:0] Wgt_3_173,input [WEIGHT_SIZE-1:0] Wgt_3_174,input [WEIGHT_SIZE-1:0] Wgt_3_175,input [WEIGHT_SIZE-1:0] Wgt_3_176,input [WEIGHT_SIZE-1:0] Wgt_3_177,input [WEIGHT_SIZE-1:0] Wgt_3_178,input [WEIGHT_SIZE-1:0] Wgt_3_179,input [WEIGHT_SIZE-1:0] Wgt_3_180,input [WEIGHT_SIZE-1:0] Wgt_3_181,input [WEIGHT_SIZE-1:0] Wgt_3_182,input [WEIGHT_SIZE-1:0] Wgt_3_183,input [WEIGHT_SIZE-1:0] Wgt_3_184,input [WEIGHT_SIZE-1:0] Wgt_3_185,input [WEIGHT_SIZE-1:0] Wgt_3_186,input [WEIGHT_SIZE-1:0] Wgt_3_187,input [WEIGHT_SIZE-1:0] Wgt_3_188,input [WEIGHT_SIZE-1:0] Wgt_3_189,input [WEIGHT_SIZE-1:0] Wgt_3_190,input [WEIGHT_SIZE-1:0] Wgt_3_191,input [WEIGHT_SIZE-1:0] Wgt_3_192,input [WEIGHT_SIZE-1:0] Wgt_3_193,input [WEIGHT_SIZE-1:0] Wgt_3_194,input [WEIGHT_SIZE-1:0] Wgt_3_195,input [WEIGHT_SIZE-1:0] Wgt_3_196,input [WEIGHT_SIZE-1:0] Wgt_3_197,input [WEIGHT_SIZE-1:0] Wgt_3_198,input [WEIGHT_SIZE-1:0] Wgt_3_199,input [WEIGHT_SIZE-1:0] Wgt_3_200,input [WEIGHT_SIZE-1:0] Wgt_3_201,input [WEIGHT_SIZE-1:0] Wgt_3_202,input [WEIGHT_SIZE-1:0] Wgt_3_203,input [WEIGHT_SIZE-1:0] Wgt_3_204,input [WEIGHT_SIZE-1:0] Wgt_3_205,input [WEIGHT_SIZE-1:0] Wgt_3_206,input [WEIGHT_SIZE-1:0] Wgt_3_207,input [WEIGHT_SIZE-1:0] Wgt_3_208,input [WEIGHT_SIZE-1:0] Wgt_3_209,input [WEIGHT_SIZE-1:0] Wgt_3_210,input [WEIGHT_SIZE-1:0] Wgt_3_211,input [WEIGHT_SIZE-1:0] Wgt_3_212,input [WEIGHT_SIZE-1:0] Wgt_3_213,input [WEIGHT_SIZE-1:0] Wgt_3_214,input [WEIGHT_SIZE-1:0] Wgt_3_215,input [WEIGHT_SIZE-1:0] Wgt_3_216,input [WEIGHT_SIZE-1:0] Wgt_3_217,input [WEIGHT_SIZE-1:0] Wgt_3_218,input [WEIGHT_SIZE-1:0] Wgt_3_219,input [WEIGHT_SIZE-1:0] Wgt_3_220,input [WEIGHT_SIZE-1:0] Wgt_3_221,input [WEIGHT_SIZE-1:0] Wgt_3_222,input [WEIGHT_SIZE-1:0] Wgt_3_223,input [WEIGHT_SIZE-1:0] Wgt_3_224,input [WEIGHT_SIZE-1:0] Wgt_3_225,input [WEIGHT_SIZE-1:0] Wgt_3_226,input [WEIGHT_SIZE-1:0] Wgt_3_227,input [WEIGHT_SIZE-1:0] Wgt_3_228,input [WEIGHT_SIZE-1:0] Wgt_3_229,input [WEIGHT_SIZE-1:0] Wgt_3_230,input [WEIGHT_SIZE-1:0] Wgt_3_231,input [WEIGHT_SIZE-1:0] Wgt_3_232,input [WEIGHT_SIZE-1:0] Wgt_3_233,input [WEIGHT_SIZE-1:0] Wgt_3_234,input [WEIGHT_SIZE-1:0] Wgt_3_235,input [WEIGHT_SIZE-1:0] Wgt_3_236,input [WEIGHT_SIZE-1:0] Wgt_3_237,input [WEIGHT_SIZE-1:0] Wgt_3_238,input [WEIGHT_SIZE-1:0] Wgt_3_239,input [WEIGHT_SIZE-1:0] Wgt_3_240,input [WEIGHT_SIZE-1:0] Wgt_3_241,input [WEIGHT_SIZE-1:0] Wgt_3_242,input [WEIGHT_SIZE-1:0] Wgt_3_243,input [WEIGHT_SIZE-1:0] Wgt_3_244,input [WEIGHT_SIZE-1:0] Wgt_3_245,input [WEIGHT_SIZE-1:0] Wgt_3_246,input [WEIGHT_SIZE-1:0] Wgt_3_247,input [WEIGHT_SIZE-1:0] Wgt_3_248,input [WEIGHT_SIZE-1:0] Wgt_3_249,input [WEIGHT_SIZE-1:0] Wgt_3_250,input [WEIGHT_SIZE-1:0] Wgt_3_251,input [WEIGHT_SIZE-1:0] Wgt_3_252,input [WEIGHT_SIZE-1:0] Wgt_3_253,input [WEIGHT_SIZE-1:0] Wgt_3_254,input [WEIGHT_SIZE-1:0] Wgt_3_255,input [WEIGHT_SIZE-1:0] Wgt_3_256,input [WEIGHT_SIZE-1:0] Wgt_3_257,input [WEIGHT_SIZE-1:0] Wgt_3_258,input [WEIGHT_SIZE-1:0] Wgt_3_259,input [WEIGHT_SIZE-1:0] Wgt_3_260,input [WEIGHT_SIZE-1:0] Wgt_3_261,input [WEIGHT_SIZE-1:0] Wgt_3_262,input [WEIGHT_SIZE-1:0] Wgt_3_263,input [WEIGHT_SIZE-1:0] Wgt_3_264,input [WEIGHT_SIZE-1:0] Wgt_3_265,input [WEIGHT_SIZE-1:0] Wgt_3_266,input [WEIGHT_SIZE-1:0] Wgt_3_267,input [WEIGHT_SIZE-1:0] Wgt_3_268,input [WEIGHT_SIZE-1:0] Wgt_3_269,input [WEIGHT_SIZE-1:0] Wgt_3_270,input [WEIGHT_SIZE-1:0] Wgt_3_271,input [WEIGHT_SIZE-1:0] Wgt_3_272,input [WEIGHT_SIZE-1:0] Wgt_3_273,input [WEIGHT_SIZE-1:0] Wgt_3_274,input [WEIGHT_SIZE-1:0] Wgt_3_275,input [WEIGHT_SIZE-1:0] Wgt_3_276,input [WEIGHT_SIZE-1:0] Wgt_3_277,input [WEIGHT_SIZE-1:0] Wgt_3_278,input [WEIGHT_SIZE-1:0] Wgt_3_279,input [WEIGHT_SIZE-1:0] Wgt_3_280,input [WEIGHT_SIZE-1:0] Wgt_3_281,input [WEIGHT_SIZE-1:0] Wgt_3_282,input [WEIGHT_SIZE-1:0] Wgt_3_283,input [WEIGHT_SIZE-1:0] Wgt_3_284,input [WEIGHT_SIZE-1:0] Wgt_3_285,input [WEIGHT_SIZE-1:0] Wgt_3_286,input [WEIGHT_SIZE-1:0] Wgt_3_287,input [WEIGHT_SIZE-1:0] Wgt_3_288,input [WEIGHT_SIZE-1:0] Wgt_3_289,input [WEIGHT_SIZE-1:0] Wgt_3_290,input [WEIGHT_SIZE-1:0] Wgt_3_291,input [WEIGHT_SIZE-1:0] Wgt_3_292,input [WEIGHT_SIZE-1:0] Wgt_3_293,input [WEIGHT_SIZE-1:0] Wgt_3_294,input [WEIGHT_SIZE-1:0] Wgt_3_295,input [WEIGHT_SIZE-1:0] Wgt_3_296,input [WEIGHT_SIZE-1:0] Wgt_3_297,input [WEIGHT_SIZE-1:0] Wgt_3_298,input [WEIGHT_SIZE-1:0] Wgt_3_299,input [WEIGHT_SIZE-1:0] Wgt_3_300,input [WEIGHT_SIZE-1:0] Wgt_3_301,input [WEIGHT_SIZE-1:0] Wgt_3_302,input [WEIGHT_SIZE-1:0] Wgt_3_303,input [WEIGHT_SIZE-1:0] Wgt_3_304,input [WEIGHT_SIZE-1:0] Wgt_3_305,input [WEIGHT_SIZE-1:0] Wgt_3_306,input [WEIGHT_SIZE-1:0] Wgt_3_307,input [WEIGHT_SIZE-1:0] Wgt_3_308,input [WEIGHT_SIZE-1:0] Wgt_3_309,input [WEIGHT_SIZE-1:0] Wgt_3_310,input [WEIGHT_SIZE-1:0] Wgt_3_311,input [WEIGHT_SIZE-1:0] Wgt_3_312,input [WEIGHT_SIZE-1:0] Wgt_3_313,input [WEIGHT_SIZE-1:0] Wgt_3_314,input [WEIGHT_SIZE-1:0] Wgt_3_315,input [WEIGHT_SIZE-1:0] Wgt_3_316,input [WEIGHT_SIZE-1:0] Wgt_3_317,input [WEIGHT_SIZE-1:0] Wgt_3_318,input [WEIGHT_SIZE-1:0] Wgt_3_319,input [WEIGHT_SIZE-1:0] Wgt_3_320,input [WEIGHT_SIZE-1:0] Wgt_3_321,input [WEIGHT_SIZE-1:0] Wgt_3_322,input [WEIGHT_SIZE-1:0] Wgt_3_323,input [WEIGHT_SIZE-1:0] Wgt_3_324,input [WEIGHT_SIZE-1:0] Wgt_3_325,input [WEIGHT_SIZE-1:0] Wgt_3_326,input [WEIGHT_SIZE-1:0] Wgt_3_327,input [WEIGHT_SIZE-1:0] Wgt_3_328,input [WEIGHT_SIZE-1:0] Wgt_3_329,input [WEIGHT_SIZE-1:0] Wgt_3_330,input [WEIGHT_SIZE-1:0] Wgt_3_331,input [WEIGHT_SIZE-1:0] Wgt_3_332,input [WEIGHT_SIZE-1:0] Wgt_3_333,input [WEIGHT_SIZE-1:0] Wgt_3_334,input [WEIGHT_SIZE-1:0] Wgt_3_335,input [WEIGHT_SIZE-1:0] Wgt_3_336,input [WEIGHT_SIZE-1:0] Wgt_3_337,input [WEIGHT_SIZE-1:0] Wgt_3_338,input [WEIGHT_SIZE-1:0] Wgt_3_339,input [WEIGHT_SIZE-1:0] Wgt_3_340,input [WEIGHT_SIZE-1:0] Wgt_3_341,input [WEIGHT_SIZE-1:0] Wgt_3_342,input [WEIGHT_SIZE-1:0] Wgt_3_343,input [WEIGHT_SIZE-1:0] Wgt_3_344,input [WEIGHT_SIZE-1:0] Wgt_3_345,input [WEIGHT_SIZE-1:0] Wgt_3_346,input [WEIGHT_SIZE-1:0] Wgt_3_347,input [WEIGHT_SIZE-1:0] Wgt_3_348,input [WEIGHT_SIZE-1:0] Wgt_3_349,input [WEIGHT_SIZE-1:0] Wgt_3_350,input [WEIGHT_SIZE-1:0] Wgt_3_351,input [WEIGHT_SIZE-1:0] Wgt_3_352,input [WEIGHT_SIZE-1:0] Wgt_3_353,input [WEIGHT_SIZE-1:0] Wgt_3_354,input [WEIGHT_SIZE-1:0] Wgt_3_355,input [WEIGHT_SIZE-1:0] Wgt_3_356,input [WEIGHT_SIZE-1:0] Wgt_3_357,input [WEIGHT_SIZE-1:0] Wgt_3_358,input [WEIGHT_SIZE-1:0] Wgt_3_359,input [WEIGHT_SIZE-1:0] Wgt_3_360,input [WEIGHT_SIZE-1:0] Wgt_3_361,input [WEIGHT_SIZE-1:0] Wgt_3_362,input [WEIGHT_SIZE-1:0] Wgt_3_363,input [WEIGHT_SIZE-1:0] Wgt_3_364,input [WEIGHT_SIZE-1:0] Wgt_3_365,input [WEIGHT_SIZE-1:0] Wgt_3_366,input [WEIGHT_SIZE-1:0] Wgt_3_367,input [WEIGHT_SIZE-1:0] Wgt_3_368,input [WEIGHT_SIZE-1:0] Wgt_3_369,input [WEIGHT_SIZE-1:0] Wgt_3_370,input [WEIGHT_SIZE-1:0] Wgt_3_371,input [WEIGHT_SIZE-1:0] Wgt_3_372,input [WEIGHT_SIZE-1:0] Wgt_3_373,input [WEIGHT_SIZE-1:0] Wgt_3_374,input [WEIGHT_SIZE-1:0] Wgt_3_375,input [WEIGHT_SIZE-1:0] Wgt_3_376,input [WEIGHT_SIZE-1:0] Wgt_3_377,input [WEIGHT_SIZE-1:0] Wgt_3_378,input [WEIGHT_SIZE-1:0] Wgt_3_379,input [WEIGHT_SIZE-1:0] Wgt_3_380,input [WEIGHT_SIZE-1:0] Wgt_3_381,input [WEIGHT_SIZE-1:0] Wgt_3_382,input [WEIGHT_SIZE-1:0] Wgt_3_383,input [WEIGHT_SIZE-1:0] Wgt_3_384,input [WEIGHT_SIZE-1:0] Wgt_3_385,input [WEIGHT_SIZE-1:0] Wgt_3_386,input [WEIGHT_SIZE-1:0] Wgt_3_387,input [WEIGHT_SIZE-1:0] Wgt_3_388,input [WEIGHT_SIZE-1:0] Wgt_3_389,input [WEIGHT_SIZE-1:0] Wgt_3_390,input [WEIGHT_SIZE-1:0] Wgt_3_391,input [WEIGHT_SIZE-1:0] Wgt_3_392,input [WEIGHT_SIZE-1:0] Wgt_3_393,input [WEIGHT_SIZE-1:0] Wgt_3_394,input [WEIGHT_SIZE-1:0] Wgt_3_395,input [WEIGHT_SIZE-1:0] Wgt_3_396,input [WEIGHT_SIZE-1:0] Wgt_3_397,input [WEIGHT_SIZE-1:0] Wgt_3_398,input [WEIGHT_SIZE-1:0] Wgt_3_399,input [WEIGHT_SIZE-1:0] Wgt_3_400,input [WEIGHT_SIZE-1:0] Wgt_3_401,input [WEIGHT_SIZE-1:0] Wgt_3_402,input [WEIGHT_SIZE-1:0] Wgt_3_403,input [WEIGHT_SIZE-1:0] Wgt_3_404,input [WEIGHT_SIZE-1:0] Wgt_3_405,input [WEIGHT_SIZE-1:0] Wgt_3_406,input [WEIGHT_SIZE-1:0] Wgt_3_407,input [WEIGHT_SIZE-1:0] Wgt_3_408,input [WEIGHT_SIZE-1:0] Wgt_3_409,input [WEIGHT_SIZE-1:0] Wgt_3_410,input [WEIGHT_SIZE-1:0] Wgt_3_411,input [WEIGHT_SIZE-1:0] Wgt_3_412,input [WEIGHT_SIZE-1:0] Wgt_3_413,input [WEIGHT_SIZE-1:0] Wgt_3_414,input [WEIGHT_SIZE-1:0] Wgt_3_415,input [WEIGHT_SIZE-1:0] Wgt_3_416,input [WEIGHT_SIZE-1:0] Wgt_3_417,input [WEIGHT_SIZE-1:0] Wgt_3_418,input [WEIGHT_SIZE-1:0] Wgt_3_419,input [WEIGHT_SIZE-1:0] Wgt_3_420,input [WEIGHT_SIZE-1:0] Wgt_3_421,input [WEIGHT_SIZE-1:0] Wgt_3_422,input [WEIGHT_SIZE-1:0] Wgt_3_423,input [WEIGHT_SIZE-1:0] Wgt_3_424,input [WEIGHT_SIZE-1:0] Wgt_3_425,input [WEIGHT_SIZE-1:0] Wgt_3_426,input [WEIGHT_SIZE-1:0] Wgt_3_427,input [WEIGHT_SIZE-1:0] Wgt_3_428,input [WEIGHT_SIZE-1:0] Wgt_3_429,input [WEIGHT_SIZE-1:0] Wgt_3_430,input [WEIGHT_SIZE-1:0] Wgt_3_431,input [WEIGHT_SIZE-1:0] Wgt_3_432,input [WEIGHT_SIZE-1:0] Wgt_3_433,input [WEIGHT_SIZE-1:0] Wgt_3_434,input [WEIGHT_SIZE-1:0] Wgt_3_435,input [WEIGHT_SIZE-1:0] Wgt_3_436,input [WEIGHT_SIZE-1:0] Wgt_3_437,input [WEIGHT_SIZE-1:0] Wgt_3_438,input [WEIGHT_SIZE-1:0] Wgt_3_439,input [WEIGHT_SIZE-1:0] Wgt_3_440,input [WEIGHT_SIZE-1:0] Wgt_3_441,input [WEIGHT_SIZE-1:0] Wgt_3_442,input [WEIGHT_SIZE-1:0] Wgt_3_443,input [WEIGHT_SIZE-1:0] Wgt_3_444,input [WEIGHT_SIZE-1:0] Wgt_3_445,input [WEIGHT_SIZE-1:0] Wgt_3_446,input [WEIGHT_SIZE-1:0] Wgt_3_447,input [WEIGHT_SIZE-1:0] Wgt_3_448,input [WEIGHT_SIZE-1:0] Wgt_3_449,input [WEIGHT_SIZE-1:0] Wgt_3_450,input [WEIGHT_SIZE-1:0] Wgt_3_451,input [WEIGHT_SIZE-1:0] Wgt_3_452,input [WEIGHT_SIZE-1:0] Wgt_3_453,input [WEIGHT_SIZE-1:0] Wgt_3_454,input [WEIGHT_SIZE-1:0] Wgt_3_455,input [WEIGHT_SIZE-1:0] Wgt_3_456,input [WEIGHT_SIZE-1:0] Wgt_3_457,input [WEIGHT_SIZE-1:0] Wgt_3_458,input [WEIGHT_SIZE-1:0] Wgt_3_459,input [WEIGHT_SIZE-1:0] Wgt_3_460,input [WEIGHT_SIZE-1:0] Wgt_3_461,input [WEIGHT_SIZE-1:0] Wgt_3_462,input [WEIGHT_SIZE-1:0] Wgt_3_463,input [WEIGHT_SIZE-1:0] Wgt_3_464,input [WEIGHT_SIZE-1:0] Wgt_3_465,input [WEIGHT_SIZE-1:0] Wgt_3_466,input [WEIGHT_SIZE-1:0] Wgt_3_467,input [WEIGHT_SIZE-1:0] Wgt_3_468,input [WEIGHT_SIZE-1:0] Wgt_3_469,input [WEIGHT_SIZE-1:0] Wgt_3_470,input [WEIGHT_SIZE-1:0] Wgt_3_471,input [WEIGHT_SIZE-1:0] Wgt_3_472,input [WEIGHT_SIZE-1:0] Wgt_3_473,input [WEIGHT_SIZE-1:0] Wgt_3_474,input [WEIGHT_SIZE-1:0] Wgt_3_475,input [WEIGHT_SIZE-1:0] Wgt_3_476,input [WEIGHT_SIZE-1:0] Wgt_3_477,input [WEIGHT_SIZE-1:0] Wgt_3_478,input [WEIGHT_SIZE-1:0] Wgt_3_479,input [WEIGHT_SIZE-1:0] Wgt_3_480,input [WEIGHT_SIZE-1:0] Wgt_3_481,input [WEIGHT_SIZE-1:0] Wgt_3_482,input [WEIGHT_SIZE-1:0] Wgt_3_483,input [WEIGHT_SIZE-1:0] Wgt_3_484,input [WEIGHT_SIZE-1:0] Wgt_3_485,input [WEIGHT_SIZE-1:0] Wgt_3_486,input [WEIGHT_SIZE-1:0] Wgt_3_487,input [WEIGHT_SIZE-1:0] Wgt_3_488,input [WEIGHT_SIZE-1:0] Wgt_3_489,input [WEIGHT_SIZE-1:0] Wgt_3_490,input [WEIGHT_SIZE-1:0] Wgt_3_491,input [WEIGHT_SIZE-1:0] Wgt_3_492,input [WEIGHT_SIZE-1:0] Wgt_3_493,input [WEIGHT_SIZE-1:0] Wgt_3_494,input [WEIGHT_SIZE-1:0] Wgt_3_495,input [WEIGHT_SIZE-1:0] Wgt_3_496,input [WEIGHT_SIZE-1:0] Wgt_3_497,input [WEIGHT_SIZE-1:0] Wgt_3_498,input [WEIGHT_SIZE-1:0] Wgt_3_499,input [WEIGHT_SIZE-1:0] Wgt_3_500,input [WEIGHT_SIZE-1:0] Wgt_3_501,input [WEIGHT_SIZE-1:0] Wgt_3_502,input [WEIGHT_SIZE-1:0] Wgt_3_503,input [WEIGHT_SIZE-1:0] Wgt_3_504,input [WEIGHT_SIZE-1:0] Wgt_3_505,input [WEIGHT_SIZE-1:0] Wgt_3_506,input [WEIGHT_SIZE-1:0] Wgt_3_507,input [WEIGHT_SIZE-1:0] Wgt_3_508,input [WEIGHT_SIZE-1:0] Wgt_3_509,input [WEIGHT_SIZE-1:0] Wgt_3_510,input [WEIGHT_SIZE-1:0] Wgt_3_511,input [WEIGHT_SIZE-1:0] Wgt_3_512,input [WEIGHT_SIZE-1:0] Wgt_3_513,input [WEIGHT_SIZE-1:0] Wgt_3_514,input [WEIGHT_SIZE-1:0] Wgt_3_515,input [WEIGHT_SIZE-1:0] Wgt_3_516,input [WEIGHT_SIZE-1:0] Wgt_3_517,input [WEIGHT_SIZE-1:0] Wgt_3_518,input [WEIGHT_SIZE-1:0] Wgt_3_519,input [WEIGHT_SIZE-1:0] Wgt_3_520,input [WEIGHT_SIZE-1:0] Wgt_3_521,input [WEIGHT_SIZE-1:0] Wgt_3_522,input [WEIGHT_SIZE-1:0] Wgt_3_523,input [WEIGHT_SIZE-1:0] Wgt_3_524,input [WEIGHT_SIZE-1:0] Wgt_3_525,input [WEIGHT_SIZE-1:0] Wgt_3_526,input [WEIGHT_SIZE-1:0] Wgt_3_527,input [WEIGHT_SIZE-1:0] Wgt_3_528,input [WEIGHT_SIZE-1:0] Wgt_3_529,input [WEIGHT_SIZE-1:0] Wgt_3_530,input [WEIGHT_SIZE-1:0] Wgt_3_531,input [WEIGHT_SIZE-1:0] Wgt_3_532,input [WEIGHT_SIZE-1:0] Wgt_3_533,input [WEIGHT_SIZE-1:0] Wgt_3_534,input [WEIGHT_SIZE-1:0] Wgt_3_535,input [WEIGHT_SIZE-1:0] Wgt_3_536,input [WEIGHT_SIZE-1:0] Wgt_3_537,input [WEIGHT_SIZE-1:0] Wgt_3_538,input [WEIGHT_SIZE-1:0] Wgt_3_539,input [WEIGHT_SIZE-1:0] Wgt_3_540,input [WEIGHT_SIZE-1:0] Wgt_3_541,input [WEIGHT_SIZE-1:0] Wgt_3_542,input [WEIGHT_SIZE-1:0] Wgt_3_543,input [WEIGHT_SIZE-1:0] Wgt_3_544,input [WEIGHT_SIZE-1:0] Wgt_3_545,input [WEIGHT_SIZE-1:0] Wgt_3_546,input [WEIGHT_SIZE-1:0] Wgt_3_547,input [WEIGHT_SIZE-1:0] Wgt_3_548,input [WEIGHT_SIZE-1:0] Wgt_3_549,input [WEIGHT_SIZE-1:0] Wgt_3_550,input [WEIGHT_SIZE-1:0] Wgt_3_551,input [WEIGHT_SIZE-1:0] Wgt_3_552,input [WEIGHT_SIZE-1:0] Wgt_3_553,input [WEIGHT_SIZE-1:0] Wgt_3_554,input [WEIGHT_SIZE-1:0] Wgt_3_555,input [WEIGHT_SIZE-1:0] Wgt_3_556,input [WEIGHT_SIZE-1:0] Wgt_3_557,input [WEIGHT_SIZE-1:0] Wgt_3_558,input [WEIGHT_SIZE-1:0] Wgt_3_559,input [WEIGHT_SIZE-1:0] Wgt_3_560,input [WEIGHT_SIZE-1:0] Wgt_3_561,input [WEIGHT_SIZE-1:0] Wgt_3_562,input [WEIGHT_SIZE-1:0] Wgt_3_563,input [WEIGHT_SIZE-1:0] Wgt_3_564,input [WEIGHT_SIZE-1:0] Wgt_3_565,input [WEIGHT_SIZE-1:0] Wgt_3_566,input [WEIGHT_SIZE-1:0] Wgt_3_567,input [WEIGHT_SIZE-1:0] Wgt_3_568,input [WEIGHT_SIZE-1:0] Wgt_3_569,input [WEIGHT_SIZE-1:0] Wgt_3_570,input [WEIGHT_SIZE-1:0] Wgt_3_571,input [WEIGHT_SIZE-1:0] Wgt_3_572,input [WEIGHT_SIZE-1:0] Wgt_3_573,input [WEIGHT_SIZE-1:0] Wgt_3_574,input [WEIGHT_SIZE-1:0] Wgt_3_575,input [WEIGHT_SIZE-1:0] Wgt_3_576,input [WEIGHT_SIZE-1:0] Wgt_3_577,input [WEIGHT_SIZE-1:0] Wgt_3_578,input [WEIGHT_SIZE-1:0] Wgt_3_579,input [WEIGHT_SIZE-1:0] Wgt_3_580,input [WEIGHT_SIZE-1:0] Wgt_3_581,input [WEIGHT_SIZE-1:0] Wgt_3_582,input [WEIGHT_SIZE-1:0] Wgt_3_583,input [WEIGHT_SIZE-1:0] Wgt_3_584,input [WEIGHT_SIZE-1:0] Wgt_3_585,input [WEIGHT_SIZE-1:0] Wgt_3_586,input [WEIGHT_SIZE-1:0] Wgt_3_587,input [WEIGHT_SIZE-1:0] Wgt_3_588,input [WEIGHT_SIZE-1:0] Wgt_3_589,input [WEIGHT_SIZE-1:0] Wgt_3_590,input [WEIGHT_SIZE-1:0] Wgt_3_591,input [WEIGHT_SIZE-1:0] Wgt_3_592,input [WEIGHT_SIZE-1:0] Wgt_3_593,input [WEIGHT_SIZE-1:0] Wgt_3_594,input [WEIGHT_SIZE-1:0] Wgt_3_595,input [WEIGHT_SIZE-1:0] Wgt_3_596,input [WEIGHT_SIZE-1:0] Wgt_3_597,input [WEIGHT_SIZE-1:0] Wgt_3_598,input [WEIGHT_SIZE-1:0] Wgt_3_599,input [WEIGHT_SIZE-1:0] Wgt_3_600,input [WEIGHT_SIZE-1:0] Wgt_3_601,input [WEIGHT_SIZE-1:0] Wgt_3_602,input [WEIGHT_SIZE-1:0] Wgt_3_603,input [WEIGHT_SIZE-1:0] Wgt_3_604,input [WEIGHT_SIZE-1:0] Wgt_3_605,input [WEIGHT_SIZE-1:0] Wgt_3_606,input [WEIGHT_SIZE-1:0] Wgt_3_607,input [WEIGHT_SIZE-1:0] Wgt_3_608,input [WEIGHT_SIZE-1:0] Wgt_3_609,input [WEIGHT_SIZE-1:0] Wgt_3_610,input [WEIGHT_SIZE-1:0] Wgt_3_611,input [WEIGHT_SIZE-1:0] Wgt_3_612,input [WEIGHT_SIZE-1:0] Wgt_3_613,input [WEIGHT_SIZE-1:0] Wgt_3_614,input [WEIGHT_SIZE-1:0] Wgt_3_615,input [WEIGHT_SIZE-1:0] Wgt_3_616,input [WEIGHT_SIZE-1:0] Wgt_3_617,input [WEIGHT_SIZE-1:0] Wgt_3_618,input [WEIGHT_SIZE-1:0] Wgt_3_619,input [WEIGHT_SIZE-1:0] Wgt_3_620,input [WEIGHT_SIZE-1:0] Wgt_3_621,input [WEIGHT_SIZE-1:0] Wgt_3_622,input [WEIGHT_SIZE-1:0] Wgt_3_623,input [WEIGHT_SIZE-1:0] Wgt_3_624,input [WEIGHT_SIZE-1:0] Wgt_3_625,input [WEIGHT_SIZE-1:0] Wgt_3_626,input [WEIGHT_SIZE-1:0] Wgt_3_627,input [WEIGHT_SIZE-1:0] Wgt_3_628,input [WEIGHT_SIZE-1:0] Wgt_3_629,input [WEIGHT_SIZE-1:0] Wgt_3_630,input [WEIGHT_SIZE-1:0] Wgt_3_631,input [WEIGHT_SIZE-1:0] Wgt_3_632,input [WEIGHT_SIZE-1:0] Wgt_3_633,input [WEIGHT_SIZE-1:0] Wgt_3_634,input [WEIGHT_SIZE-1:0] Wgt_3_635,input [WEIGHT_SIZE-1:0] Wgt_3_636,input [WEIGHT_SIZE-1:0] Wgt_3_637,input [WEIGHT_SIZE-1:0] Wgt_3_638,input [WEIGHT_SIZE-1:0] Wgt_3_639,input [WEIGHT_SIZE-1:0] Wgt_3_640,input [WEIGHT_SIZE-1:0] Wgt_3_641,input [WEIGHT_SIZE-1:0] Wgt_3_642,input [WEIGHT_SIZE-1:0] Wgt_3_643,input [WEIGHT_SIZE-1:0] Wgt_3_644,input [WEIGHT_SIZE-1:0] Wgt_3_645,input [WEIGHT_SIZE-1:0] Wgt_3_646,input [WEIGHT_SIZE-1:0] Wgt_3_647,input [WEIGHT_SIZE-1:0] Wgt_3_648,input [WEIGHT_SIZE-1:0] Wgt_3_649,input [WEIGHT_SIZE-1:0] Wgt_3_650,input [WEIGHT_SIZE-1:0] Wgt_3_651,input [WEIGHT_SIZE-1:0] Wgt_3_652,input [WEIGHT_SIZE-1:0] Wgt_3_653,input [WEIGHT_SIZE-1:0] Wgt_3_654,input [WEIGHT_SIZE-1:0] Wgt_3_655,input [WEIGHT_SIZE-1:0] Wgt_3_656,input [WEIGHT_SIZE-1:0] Wgt_3_657,input [WEIGHT_SIZE-1:0] Wgt_3_658,input [WEIGHT_SIZE-1:0] Wgt_3_659,input [WEIGHT_SIZE-1:0] Wgt_3_660,input [WEIGHT_SIZE-1:0] Wgt_3_661,input [WEIGHT_SIZE-1:0] Wgt_3_662,input [WEIGHT_SIZE-1:0] Wgt_3_663,input [WEIGHT_SIZE-1:0] Wgt_3_664,input [WEIGHT_SIZE-1:0] Wgt_3_665,input [WEIGHT_SIZE-1:0] Wgt_3_666,input [WEIGHT_SIZE-1:0] Wgt_3_667,input [WEIGHT_SIZE-1:0] Wgt_3_668,input [WEIGHT_SIZE-1:0] Wgt_3_669,input [WEIGHT_SIZE-1:0] Wgt_3_670,input [WEIGHT_SIZE-1:0] Wgt_3_671,input [WEIGHT_SIZE-1:0] Wgt_3_672,input [WEIGHT_SIZE-1:0] Wgt_3_673,input [WEIGHT_SIZE-1:0] Wgt_3_674,input [WEIGHT_SIZE-1:0] Wgt_3_675,input [WEIGHT_SIZE-1:0] Wgt_3_676,input [WEIGHT_SIZE-1:0] Wgt_3_677,input [WEIGHT_SIZE-1:0] Wgt_3_678,input [WEIGHT_SIZE-1:0] Wgt_3_679,input [WEIGHT_SIZE-1:0] Wgt_3_680,input [WEIGHT_SIZE-1:0] Wgt_3_681,input [WEIGHT_SIZE-1:0] Wgt_3_682,input [WEIGHT_SIZE-1:0] Wgt_3_683,input [WEIGHT_SIZE-1:0] Wgt_3_684,input [WEIGHT_SIZE-1:0] Wgt_3_685,input [WEIGHT_SIZE-1:0] Wgt_3_686,input [WEIGHT_SIZE-1:0] Wgt_3_687,input [WEIGHT_SIZE-1:0] Wgt_3_688,input [WEIGHT_SIZE-1:0] Wgt_3_689,input [WEIGHT_SIZE-1:0] Wgt_3_690,input [WEIGHT_SIZE-1:0] Wgt_3_691,input [WEIGHT_SIZE-1:0] Wgt_3_692,input [WEIGHT_SIZE-1:0] Wgt_3_693,input [WEIGHT_SIZE-1:0] Wgt_3_694,input [WEIGHT_SIZE-1:0] Wgt_3_695,input [WEIGHT_SIZE-1:0] Wgt_3_696,input [WEIGHT_SIZE-1:0] Wgt_3_697,input [WEIGHT_SIZE-1:0] Wgt_3_698,input [WEIGHT_SIZE-1:0] Wgt_3_699,input [WEIGHT_SIZE-1:0] Wgt_3_700,input [WEIGHT_SIZE-1:0] Wgt_3_701,input [WEIGHT_SIZE-1:0] Wgt_3_702,input [WEIGHT_SIZE-1:0] Wgt_3_703,input [WEIGHT_SIZE-1:0] Wgt_3_704,input [WEIGHT_SIZE-1:0] Wgt_3_705,input [WEIGHT_SIZE-1:0] Wgt_3_706,input [WEIGHT_SIZE-1:0] Wgt_3_707,input [WEIGHT_SIZE-1:0] Wgt_3_708,input [WEIGHT_SIZE-1:0] Wgt_3_709,input [WEIGHT_SIZE-1:0] Wgt_3_710,input [WEIGHT_SIZE-1:0] Wgt_3_711,input [WEIGHT_SIZE-1:0] Wgt_3_712,input [WEIGHT_SIZE-1:0] Wgt_3_713,input [WEIGHT_SIZE-1:0] Wgt_3_714,input [WEIGHT_SIZE-1:0] Wgt_3_715,input [WEIGHT_SIZE-1:0] Wgt_3_716,input [WEIGHT_SIZE-1:0] Wgt_3_717,input [WEIGHT_SIZE-1:0] Wgt_3_718,input [WEIGHT_SIZE-1:0] Wgt_3_719,input [WEIGHT_SIZE-1:0] Wgt_3_720,input [WEIGHT_SIZE-1:0] Wgt_3_721,input [WEIGHT_SIZE-1:0] Wgt_3_722,input [WEIGHT_SIZE-1:0] Wgt_3_723,input [WEIGHT_SIZE-1:0] Wgt_3_724,input [WEIGHT_SIZE-1:0] Wgt_3_725,input [WEIGHT_SIZE-1:0] Wgt_3_726,input [WEIGHT_SIZE-1:0] Wgt_3_727,input [WEIGHT_SIZE-1:0] Wgt_3_728,input [WEIGHT_SIZE-1:0] Wgt_3_729,input [WEIGHT_SIZE-1:0] Wgt_3_730,input [WEIGHT_SIZE-1:0] Wgt_3_731,input [WEIGHT_SIZE-1:0] Wgt_3_732,input [WEIGHT_SIZE-1:0] Wgt_3_733,input [WEIGHT_SIZE-1:0] Wgt_3_734,input [WEIGHT_SIZE-1:0] Wgt_3_735,input [WEIGHT_SIZE-1:0] Wgt_3_736,input [WEIGHT_SIZE-1:0] Wgt_3_737,input [WEIGHT_SIZE-1:0] Wgt_3_738,input [WEIGHT_SIZE-1:0] Wgt_3_739,input [WEIGHT_SIZE-1:0] Wgt_3_740,input [WEIGHT_SIZE-1:0] Wgt_3_741,input [WEIGHT_SIZE-1:0] Wgt_3_742,input [WEIGHT_SIZE-1:0] Wgt_3_743,input [WEIGHT_SIZE-1:0] Wgt_3_744,input [WEIGHT_SIZE-1:0] Wgt_3_745,input [WEIGHT_SIZE-1:0] Wgt_3_746,input [WEIGHT_SIZE-1:0] Wgt_3_747,input [WEIGHT_SIZE-1:0] Wgt_3_748,input [WEIGHT_SIZE-1:0] Wgt_3_749,input [WEIGHT_SIZE-1:0] Wgt_3_750,input [WEIGHT_SIZE-1:0] Wgt_3_751,input [WEIGHT_SIZE-1:0] Wgt_3_752,input [WEIGHT_SIZE-1:0] Wgt_3_753,input [WEIGHT_SIZE-1:0] Wgt_3_754,input [WEIGHT_SIZE-1:0] Wgt_3_755,input [WEIGHT_SIZE-1:0] Wgt_3_756,input [WEIGHT_SIZE-1:0] Wgt_3_757,input [WEIGHT_SIZE-1:0] Wgt_3_758,input [WEIGHT_SIZE-1:0] Wgt_3_759,input [WEIGHT_SIZE-1:0] Wgt_3_760,input [WEIGHT_SIZE-1:0] Wgt_3_761,input [WEIGHT_SIZE-1:0] Wgt_3_762,input [WEIGHT_SIZE-1:0] Wgt_3_763,input [WEIGHT_SIZE-1:0] Wgt_3_764,input [WEIGHT_SIZE-1:0] Wgt_3_765,input [WEIGHT_SIZE-1:0] Wgt_3_766,input [WEIGHT_SIZE-1:0] Wgt_3_767,input [WEIGHT_SIZE-1:0] Wgt_3_768,input [WEIGHT_SIZE-1:0] Wgt_3_769,input [WEIGHT_SIZE-1:0] Wgt_3_770,input [WEIGHT_SIZE-1:0] Wgt_3_771,input [WEIGHT_SIZE-1:0] Wgt_3_772,input [WEIGHT_SIZE-1:0] Wgt_3_773,input [WEIGHT_SIZE-1:0] Wgt_3_774,input [WEIGHT_SIZE-1:0] Wgt_3_775,input [WEIGHT_SIZE-1:0] Wgt_3_776,input [WEIGHT_SIZE-1:0] Wgt_3_777,input [WEIGHT_SIZE-1:0] Wgt_3_778,input [WEIGHT_SIZE-1:0] Wgt_3_779,input [WEIGHT_SIZE-1:0] Wgt_3_780,input [WEIGHT_SIZE-1:0] Wgt_3_781,input [WEIGHT_SIZE-1:0] Wgt_3_782,input [WEIGHT_SIZE-1:0] Wgt_3_783,input [WEIGHT_SIZE-1:0] Wgt_3_784,input [WEIGHT_SIZE-1:0] Wgt_4_0,input [WEIGHT_SIZE-1:0] Wgt_4_1,input [WEIGHT_SIZE-1:0] Wgt_4_2,input [WEIGHT_SIZE-1:0] Wgt_4_3,input [WEIGHT_SIZE-1:0] Wgt_4_4,input [WEIGHT_SIZE-1:0] Wgt_4_5,input [WEIGHT_SIZE-1:0] Wgt_4_6,input [WEIGHT_SIZE-1:0] Wgt_4_7,input [WEIGHT_SIZE-1:0] Wgt_4_8,input [WEIGHT_SIZE-1:0] Wgt_4_9,input [WEIGHT_SIZE-1:0] Wgt_4_10,input [WEIGHT_SIZE-1:0] Wgt_4_11,input [WEIGHT_SIZE-1:0] Wgt_4_12,input [WEIGHT_SIZE-1:0] Wgt_4_13,input [WEIGHT_SIZE-1:0] Wgt_4_14,input [WEIGHT_SIZE-1:0] Wgt_4_15,input [WEIGHT_SIZE-1:0] Wgt_4_16,input [WEIGHT_SIZE-1:0] Wgt_4_17,input [WEIGHT_SIZE-1:0] Wgt_4_18,input [WEIGHT_SIZE-1:0] Wgt_4_19,input [WEIGHT_SIZE-1:0] Wgt_4_20,input [WEIGHT_SIZE-1:0] Wgt_4_21,input [WEIGHT_SIZE-1:0] Wgt_4_22,input [WEIGHT_SIZE-1:0] Wgt_4_23,input [WEIGHT_SIZE-1:0] Wgt_4_24,input [WEIGHT_SIZE-1:0] Wgt_4_25,input [WEIGHT_SIZE-1:0] Wgt_4_26,input [WEIGHT_SIZE-1:0] Wgt_4_27,input [WEIGHT_SIZE-1:0] Wgt_4_28,input [WEIGHT_SIZE-1:0] Wgt_4_29,input [WEIGHT_SIZE-1:0] Wgt_4_30,input [WEIGHT_SIZE-1:0] Wgt_4_31,input [WEIGHT_SIZE-1:0] Wgt_4_32,input [WEIGHT_SIZE-1:0] Wgt_4_33,input [WEIGHT_SIZE-1:0] Wgt_4_34,input [WEIGHT_SIZE-1:0] Wgt_4_35,input [WEIGHT_SIZE-1:0] Wgt_4_36,input [WEIGHT_SIZE-1:0] Wgt_4_37,input [WEIGHT_SIZE-1:0] Wgt_4_38,input [WEIGHT_SIZE-1:0] Wgt_4_39,input [WEIGHT_SIZE-1:0] Wgt_4_40,input [WEIGHT_SIZE-1:0] Wgt_4_41,input [WEIGHT_SIZE-1:0] Wgt_4_42,input [WEIGHT_SIZE-1:0] Wgt_4_43,input [WEIGHT_SIZE-1:0] Wgt_4_44,input [WEIGHT_SIZE-1:0] Wgt_4_45,input [WEIGHT_SIZE-1:0] Wgt_4_46,input [WEIGHT_SIZE-1:0] Wgt_4_47,input [WEIGHT_SIZE-1:0] Wgt_4_48,input [WEIGHT_SIZE-1:0] Wgt_4_49,input [WEIGHT_SIZE-1:0] Wgt_4_50,input [WEIGHT_SIZE-1:0] Wgt_4_51,input [WEIGHT_SIZE-1:0] Wgt_4_52,input [WEIGHT_SIZE-1:0] Wgt_4_53,input [WEIGHT_SIZE-1:0] Wgt_4_54,input [WEIGHT_SIZE-1:0] Wgt_4_55,input [WEIGHT_SIZE-1:0] Wgt_4_56,input [WEIGHT_SIZE-1:0] Wgt_4_57,input [WEIGHT_SIZE-1:0] Wgt_4_58,input [WEIGHT_SIZE-1:0] Wgt_4_59,input [WEIGHT_SIZE-1:0] Wgt_4_60,input [WEIGHT_SIZE-1:0] Wgt_4_61,input [WEIGHT_SIZE-1:0] Wgt_4_62,input [WEIGHT_SIZE-1:0] Wgt_4_63,input [WEIGHT_SIZE-1:0] Wgt_4_64,input [WEIGHT_SIZE-1:0] Wgt_4_65,input [WEIGHT_SIZE-1:0] Wgt_4_66,input [WEIGHT_SIZE-1:0] Wgt_4_67,input [WEIGHT_SIZE-1:0] Wgt_4_68,input [WEIGHT_SIZE-1:0] Wgt_4_69,input [WEIGHT_SIZE-1:0] Wgt_4_70,input [WEIGHT_SIZE-1:0] Wgt_4_71,input [WEIGHT_SIZE-1:0] Wgt_4_72,input [WEIGHT_SIZE-1:0] Wgt_4_73,input [WEIGHT_SIZE-1:0] Wgt_4_74,input [WEIGHT_SIZE-1:0] Wgt_4_75,input [WEIGHT_SIZE-1:0] Wgt_4_76,input [WEIGHT_SIZE-1:0] Wgt_4_77,input [WEIGHT_SIZE-1:0] Wgt_4_78,input [WEIGHT_SIZE-1:0] Wgt_4_79,input [WEIGHT_SIZE-1:0] Wgt_4_80,input [WEIGHT_SIZE-1:0] Wgt_4_81,input [WEIGHT_SIZE-1:0] Wgt_4_82,input [WEIGHT_SIZE-1:0] Wgt_4_83,input [WEIGHT_SIZE-1:0] Wgt_4_84,input [WEIGHT_SIZE-1:0] Wgt_4_85,input [WEIGHT_SIZE-1:0] Wgt_4_86,input [WEIGHT_SIZE-1:0] Wgt_4_87,input [WEIGHT_SIZE-1:0] Wgt_4_88,input [WEIGHT_SIZE-1:0] Wgt_4_89,input [WEIGHT_SIZE-1:0] Wgt_4_90,input [WEIGHT_SIZE-1:0] Wgt_4_91,input [WEIGHT_SIZE-1:0] Wgt_4_92,input [WEIGHT_SIZE-1:0] Wgt_4_93,input [WEIGHT_SIZE-1:0] Wgt_4_94,input [WEIGHT_SIZE-1:0] Wgt_4_95,input [WEIGHT_SIZE-1:0] Wgt_4_96,input [WEIGHT_SIZE-1:0] Wgt_4_97,input [WEIGHT_SIZE-1:0] Wgt_4_98,input [WEIGHT_SIZE-1:0] Wgt_4_99,input [WEIGHT_SIZE-1:0] Wgt_4_100,input [WEIGHT_SIZE-1:0] Wgt_4_101,input [WEIGHT_SIZE-1:0] Wgt_4_102,input [WEIGHT_SIZE-1:0] Wgt_4_103,input [WEIGHT_SIZE-1:0] Wgt_4_104,input [WEIGHT_SIZE-1:0] Wgt_4_105,input [WEIGHT_SIZE-1:0] Wgt_4_106,input [WEIGHT_SIZE-1:0] Wgt_4_107,input [WEIGHT_SIZE-1:0] Wgt_4_108,input [WEIGHT_SIZE-1:0] Wgt_4_109,input [WEIGHT_SIZE-1:0] Wgt_4_110,input [WEIGHT_SIZE-1:0] Wgt_4_111,input [WEIGHT_SIZE-1:0] Wgt_4_112,input [WEIGHT_SIZE-1:0] Wgt_4_113,input [WEIGHT_SIZE-1:0] Wgt_4_114,input [WEIGHT_SIZE-1:0] Wgt_4_115,input [WEIGHT_SIZE-1:0] Wgt_4_116,input [WEIGHT_SIZE-1:0] Wgt_4_117,input [WEIGHT_SIZE-1:0] Wgt_4_118,input [WEIGHT_SIZE-1:0] Wgt_4_119,input [WEIGHT_SIZE-1:0] Wgt_4_120,input [WEIGHT_SIZE-1:0] Wgt_4_121,input [WEIGHT_SIZE-1:0] Wgt_4_122,input [WEIGHT_SIZE-1:0] Wgt_4_123,input [WEIGHT_SIZE-1:0] Wgt_4_124,input [WEIGHT_SIZE-1:0] Wgt_4_125,input [WEIGHT_SIZE-1:0] Wgt_4_126,input [WEIGHT_SIZE-1:0] Wgt_4_127,input [WEIGHT_SIZE-1:0] Wgt_4_128,input [WEIGHT_SIZE-1:0] Wgt_4_129,input [WEIGHT_SIZE-1:0] Wgt_4_130,input [WEIGHT_SIZE-1:0] Wgt_4_131,input [WEIGHT_SIZE-1:0] Wgt_4_132,input [WEIGHT_SIZE-1:0] Wgt_4_133,input [WEIGHT_SIZE-1:0] Wgt_4_134,input [WEIGHT_SIZE-1:0] Wgt_4_135,input [WEIGHT_SIZE-1:0] Wgt_4_136,input [WEIGHT_SIZE-1:0] Wgt_4_137,input [WEIGHT_SIZE-1:0] Wgt_4_138,input [WEIGHT_SIZE-1:0] Wgt_4_139,input [WEIGHT_SIZE-1:0] Wgt_4_140,input [WEIGHT_SIZE-1:0] Wgt_4_141,input [WEIGHT_SIZE-1:0] Wgt_4_142,input [WEIGHT_SIZE-1:0] Wgt_4_143,input [WEIGHT_SIZE-1:0] Wgt_4_144,input [WEIGHT_SIZE-1:0] Wgt_4_145,input [WEIGHT_SIZE-1:0] Wgt_4_146,input [WEIGHT_SIZE-1:0] Wgt_4_147,input [WEIGHT_SIZE-1:0] Wgt_4_148,input [WEIGHT_SIZE-1:0] Wgt_4_149,input [WEIGHT_SIZE-1:0] Wgt_4_150,input [WEIGHT_SIZE-1:0] Wgt_4_151,input [WEIGHT_SIZE-1:0] Wgt_4_152,input [WEIGHT_SIZE-1:0] Wgt_4_153,input [WEIGHT_SIZE-1:0] Wgt_4_154,input [WEIGHT_SIZE-1:0] Wgt_4_155,input [WEIGHT_SIZE-1:0] Wgt_4_156,input [WEIGHT_SIZE-1:0] Wgt_4_157,input [WEIGHT_SIZE-1:0] Wgt_4_158,input [WEIGHT_SIZE-1:0] Wgt_4_159,input [WEIGHT_SIZE-1:0] Wgt_4_160,input [WEIGHT_SIZE-1:0] Wgt_4_161,input [WEIGHT_SIZE-1:0] Wgt_4_162,input [WEIGHT_SIZE-1:0] Wgt_4_163,input [WEIGHT_SIZE-1:0] Wgt_4_164,input [WEIGHT_SIZE-1:0] Wgt_4_165,input [WEIGHT_SIZE-1:0] Wgt_4_166,input [WEIGHT_SIZE-1:0] Wgt_4_167,input [WEIGHT_SIZE-1:0] Wgt_4_168,input [WEIGHT_SIZE-1:0] Wgt_4_169,input [WEIGHT_SIZE-1:0] Wgt_4_170,input [WEIGHT_SIZE-1:0] Wgt_4_171,input [WEIGHT_SIZE-1:0] Wgt_4_172,input [WEIGHT_SIZE-1:0] Wgt_4_173,input [WEIGHT_SIZE-1:0] Wgt_4_174,input [WEIGHT_SIZE-1:0] Wgt_4_175,input [WEIGHT_SIZE-1:0] Wgt_4_176,input [WEIGHT_SIZE-1:0] Wgt_4_177,input [WEIGHT_SIZE-1:0] Wgt_4_178,input [WEIGHT_SIZE-1:0] Wgt_4_179,input [WEIGHT_SIZE-1:0] Wgt_4_180,input [WEIGHT_SIZE-1:0] Wgt_4_181,input [WEIGHT_SIZE-1:0] Wgt_4_182,input [WEIGHT_SIZE-1:0] Wgt_4_183,input [WEIGHT_SIZE-1:0] Wgt_4_184,input [WEIGHT_SIZE-1:0] Wgt_4_185,input [WEIGHT_SIZE-1:0] Wgt_4_186,input [WEIGHT_SIZE-1:0] Wgt_4_187,input [WEIGHT_SIZE-1:0] Wgt_4_188,input [WEIGHT_SIZE-1:0] Wgt_4_189,input [WEIGHT_SIZE-1:0] Wgt_4_190,input [WEIGHT_SIZE-1:0] Wgt_4_191,input [WEIGHT_SIZE-1:0] Wgt_4_192,input [WEIGHT_SIZE-1:0] Wgt_4_193,input [WEIGHT_SIZE-1:0] Wgt_4_194,input [WEIGHT_SIZE-1:0] Wgt_4_195,input [WEIGHT_SIZE-1:0] Wgt_4_196,input [WEIGHT_SIZE-1:0] Wgt_4_197,input [WEIGHT_SIZE-1:0] Wgt_4_198,input [WEIGHT_SIZE-1:0] Wgt_4_199,input [WEIGHT_SIZE-1:0] Wgt_4_200,input [WEIGHT_SIZE-1:0] Wgt_4_201,input [WEIGHT_SIZE-1:0] Wgt_4_202,input [WEIGHT_SIZE-1:0] Wgt_4_203,input [WEIGHT_SIZE-1:0] Wgt_4_204,input [WEIGHT_SIZE-1:0] Wgt_4_205,input [WEIGHT_SIZE-1:0] Wgt_4_206,input [WEIGHT_SIZE-1:0] Wgt_4_207,input [WEIGHT_SIZE-1:0] Wgt_4_208,input [WEIGHT_SIZE-1:0] Wgt_4_209,input [WEIGHT_SIZE-1:0] Wgt_4_210,input [WEIGHT_SIZE-1:0] Wgt_4_211,input [WEIGHT_SIZE-1:0] Wgt_4_212,input [WEIGHT_SIZE-1:0] Wgt_4_213,input [WEIGHT_SIZE-1:0] Wgt_4_214,input [WEIGHT_SIZE-1:0] Wgt_4_215,input [WEIGHT_SIZE-1:0] Wgt_4_216,input [WEIGHT_SIZE-1:0] Wgt_4_217,input [WEIGHT_SIZE-1:0] Wgt_4_218,input [WEIGHT_SIZE-1:0] Wgt_4_219,input [WEIGHT_SIZE-1:0] Wgt_4_220,input [WEIGHT_SIZE-1:0] Wgt_4_221,input [WEIGHT_SIZE-1:0] Wgt_4_222,input [WEIGHT_SIZE-1:0] Wgt_4_223,input [WEIGHT_SIZE-1:0] Wgt_4_224,input [WEIGHT_SIZE-1:0] Wgt_4_225,input [WEIGHT_SIZE-1:0] Wgt_4_226,input [WEIGHT_SIZE-1:0] Wgt_4_227,input [WEIGHT_SIZE-1:0] Wgt_4_228,input [WEIGHT_SIZE-1:0] Wgt_4_229,input [WEIGHT_SIZE-1:0] Wgt_4_230,input [WEIGHT_SIZE-1:0] Wgt_4_231,input [WEIGHT_SIZE-1:0] Wgt_4_232,input [WEIGHT_SIZE-1:0] Wgt_4_233,input [WEIGHT_SIZE-1:0] Wgt_4_234,input [WEIGHT_SIZE-1:0] Wgt_4_235,input [WEIGHT_SIZE-1:0] Wgt_4_236,input [WEIGHT_SIZE-1:0] Wgt_4_237,input [WEIGHT_SIZE-1:0] Wgt_4_238,input [WEIGHT_SIZE-1:0] Wgt_4_239,input [WEIGHT_SIZE-1:0] Wgt_4_240,input [WEIGHT_SIZE-1:0] Wgt_4_241,input [WEIGHT_SIZE-1:0] Wgt_4_242,input [WEIGHT_SIZE-1:0] Wgt_4_243,input [WEIGHT_SIZE-1:0] Wgt_4_244,input [WEIGHT_SIZE-1:0] Wgt_4_245,input [WEIGHT_SIZE-1:0] Wgt_4_246,input [WEIGHT_SIZE-1:0] Wgt_4_247,input [WEIGHT_SIZE-1:0] Wgt_4_248,input [WEIGHT_SIZE-1:0] Wgt_4_249,input [WEIGHT_SIZE-1:0] Wgt_4_250,input [WEIGHT_SIZE-1:0] Wgt_4_251,input [WEIGHT_SIZE-1:0] Wgt_4_252,input [WEIGHT_SIZE-1:0] Wgt_4_253,input [WEIGHT_SIZE-1:0] Wgt_4_254,input [WEIGHT_SIZE-1:0] Wgt_4_255,input [WEIGHT_SIZE-1:0] Wgt_4_256,input [WEIGHT_SIZE-1:0] Wgt_4_257,input [WEIGHT_SIZE-1:0] Wgt_4_258,input [WEIGHT_SIZE-1:0] Wgt_4_259,input [WEIGHT_SIZE-1:0] Wgt_4_260,input [WEIGHT_SIZE-1:0] Wgt_4_261,input [WEIGHT_SIZE-1:0] Wgt_4_262,input [WEIGHT_SIZE-1:0] Wgt_4_263,input [WEIGHT_SIZE-1:0] Wgt_4_264,input [WEIGHT_SIZE-1:0] Wgt_4_265,input [WEIGHT_SIZE-1:0] Wgt_4_266,input [WEIGHT_SIZE-1:0] Wgt_4_267,input [WEIGHT_SIZE-1:0] Wgt_4_268,input [WEIGHT_SIZE-1:0] Wgt_4_269,input [WEIGHT_SIZE-1:0] Wgt_4_270,input [WEIGHT_SIZE-1:0] Wgt_4_271,input [WEIGHT_SIZE-1:0] Wgt_4_272,input [WEIGHT_SIZE-1:0] Wgt_4_273,input [WEIGHT_SIZE-1:0] Wgt_4_274,input [WEIGHT_SIZE-1:0] Wgt_4_275,input [WEIGHT_SIZE-1:0] Wgt_4_276,input [WEIGHT_SIZE-1:0] Wgt_4_277,input [WEIGHT_SIZE-1:0] Wgt_4_278,input [WEIGHT_SIZE-1:0] Wgt_4_279,input [WEIGHT_SIZE-1:0] Wgt_4_280,input [WEIGHT_SIZE-1:0] Wgt_4_281,input [WEIGHT_SIZE-1:0] Wgt_4_282,input [WEIGHT_SIZE-1:0] Wgt_4_283,input [WEIGHT_SIZE-1:0] Wgt_4_284,input [WEIGHT_SIZE-1:0] Wgt_4_285,input [WEIGHT_SIZE-1:0] Wgt_4_286,input [WEIGHT_SIZE-1:0] Wgt_4_287,input [WEIGHT_SIZE-1:0] Wgt_4_288,input [WEIGHT_SIZE-1:0] Wgt_4_289,input [WEIGHT_SIZE-1:0] Wgt_4_290,input [WEIGHT_SIZE-1:0] Wgt_4_291,input [WEIGHT_SIZE-1:0] Wgt_4_292,input [WEIGHT_SIZE-1:0] Wgt_4_293,input [WEIGHT_SIZE-1:0] Wgt_4_294,input [WEIGHT_SIZE-1:0] Wgt_4_295,input [WEIGHT_SIZE-1:0] Wgt_4_296,input [WEIGHT_SIZE-1:0] Wgt_4_297,input [WEIGHT_SIZE-1:0] Wgt_4_298,input [WEIGHT_SIZE-1:0] Wgt_4_299,input [WEIGHT_SIZE-1:0] Wgt_4_300,input [WEIGHT_SIZE-1:0] Wgt_4_301,input [WEIGHT_SIZE-1:0] Wgt_4_302,input [WEIGHT_SIZE-1:0] Wgt_4_303,input [WEIGHT_SIZE-1:0] Wgt_4_304,input [WEIGHT_SIZE-1:0] Wgt_4_305,input [WEIGHT_SIZE-1:0] Wgt_4_306,input [WEIGHT_SIZE-1:0] Wgt_4_307,input [WEIGHT_SIZE-1:0] Wgt_4_308,input [WEIGHT_SIZE-1:0] Wgt_4_309,input [WEIGHT_SIZE-1:0] Wgt_4_310,input [WEIGHT_SIZE-1:0] Wgt_4_311,input [WEIGHT_SIZE-1:0] Wgt_4_312,input [WEIGHT_SIZE-1:0] Wgt_4_313,input [WEIGHT_SIZE-1:0] Wgt_4_314,input [WEIGHT_SIZE-1:0] Wgt_4_315,input [WEIGHT_SIZE-1:0] Wgt_4_316,input [WEIGHT_SIZE-1:0] Wgt_4_317,input [WEIGHT_SIZE-1:0] Wgt_4_318,input [WEIGHT_SIZE-1:0] Wgt_4_319,input [WEIGHT_SIZE-1:0] Wgt_4_320,input [WEIGHT_SIZE-1:0] Wgt_4_321,input [WEIGHT_SIZE-1:0] Wgt_4_322,input [WEIGHT_SIZE-1:0] Wgt_4_323,input [WEIGHT_SIZE-1:0] Wgt_4_324,input [WEIGHT_SIZE-1:0] Wgt_4_325,input [WEIGHT_SIZE-1:0] Wgt_4_326,input [WEIGHT_SIZE-1:0] Wgt_4_327,input [WEIGHT_SIZE-1:0] Wgt_4_328,input [WEIGHT_SIZE-1:0] Wgt_4_329,input [WEIGHT_SIZE-1:0] Wgt_4_330,input [WEIGHT_SIZE-1:0] Wgt_4_331,input [WEIGHT_SIZE-1:0] Wgt_4_332,input [WEIGHT_SIZE-1:0] Wgt_4_333,input [WEIGHT_SIZE-1:0] Wgt_4_334,input [WEIGHT_SIZE-1:0] Wgt_4_335,input [WEIGHT_SIZE-1:0] Wgt_4_336,input [WEIGHT_SIZE-1:0] Wgt_4_337,input [WEIGHT_SIZE-1:0] Wgt_4_338,input [WEIGHT_SIZE-1:0] Wgt_4_339,input [WEIGHT_SIZE-1:0] Wgt_4_340,input [WEIGHT_SIZE-1:0] Wgt_4_341,input [WEIGHT_SIZE-1:0] Wgt_4_342,input [WEIGHT_SIZE-1:0] Wgt_4_343,input [WEIGHT_SIZE-1:0] Wgt_4_344,input [WEIGHT_SIZE-1:0] Wgt_4_345,input [WEIGHT_SIZE-1:0] Wgt_4_346,input [WEIGHT_SIZE-1:0] Wgt_4_347,input [WEIGHT_SIZE-1:0] Wgt_4_348,input [WEIGHT_SIZE-1:0] Wgt_4_349,input [WEIGHT_SIZE-1:0] Wgt_4_350,input [WEIGHT_SIZE-1:0] Wgt_4_351,input [WEIGHT_SIZE-1:0] Wgt_4_352,input [WEIGHT_SIZE-1:0] Wgt_4_353,input [WEIGHT_SIZE-1:0] Wgt_4_354,input [WEIGHT_SIZE-1:0] Wgt_4_355,input [WEIGHT_SIZE-1:0] Wgt_4_356,input [WEIGHT_SIZE-1:0] Wgt_4_357,input [WEIGHT_SIZE-1:0] Wgt_4_358,input [WEIGHT_SIZE-1:0] Wgt_4_359,input [WEIGHT_SIZE-1:0] Wgt_4_360,input [WEIGHT_SIZE-1:0] Wgt_4_361,input [WEIGHT_SIZE-1:0] Wgt_4_362,input [WEIGHT_SIZE-1:0] Wgt_4_363,input [WEIGHT_SIZE-1:0] Wgt_4_364,input [WEIGHT_SIZE-1:0] Wgt_4_365,input [WEIGHT_SIZE-1:0] Wgt_4_366,input [WEIGHT_SIZE-1:0] Wgt_4_367,input [WEIGHT_SIZE-1:0] Wgt_4_368,input [WEIGHT_SIZE-1:0] Wgt_4_369,input [WEIGHT_SIZE-1:0] Wgt_4_370,input [WEIGHT_SIZE-1:0] Wgt_4_371,input [WEIGHT_SIZE-1:0] Wgt_4_372,input [WEIGHT_SIZE-1:0] Wgt_4_373,input [WEIGHT_SIZE-1:0] Wgt_4_374,input [WEIGHT_SIZE-1:0] Wgt_4_375,input [WEIGHT_SIZE-1:0] Wgt_4_376,input [WEIGHT_SIZE-1:0] Wgt_4_377,input [WEIGHT_SIZE-1:0] Wgt_4_378,input [WEIGHT_SIZE-1:0] Wgt_4_379,input [WEIGHT_SIZE-1:0] Wgt_4_380,input [WEIGHT_SIZE-1:0] Wgt_4_381,input [WEIGHT_SIZE-1:0] Wgt_4_382,input [WEIGHT_SIZE-1:0] Wgt_4_383,input [WEIGHT_SIZE-1:0] Wgt_4_384,input [WEIGHT_SIZE-1:0] Wgt_4_385,input [WEIGHT_SIZE-1:0] Wgt_4_386,input [WEIGHT_SIZE-1:0] Wgt_4_387,input [WEIGHT_SIZE-1:0] Wgt_4_388,input [WEIGHT_SIZE-1:0] Wgt_4_389,input [WEIGHT_SIZE-1:0] Wgt_4_390,input [WEIGHT_SIZE-1:0] Wgt_4_391,input [WEIGHT_SIZE-1:0] Wgt_4_392,input [WEIGHT_SIZE-1:0] Wgt_4_393,input [WEIGHT_SIZE-1:0] Wgt_4_394,input [WEIGHT_SIZE-1:0] Wgt_4_395,input [WEIGHT_SIZE-1:0] Wgt_4_396,input [WEIGHT_SIZE-1:0] Wgt_4_397,input [WEIGHT_SIZE-1:0] Wgt_4_398,input [WEIGHT_SIZE-1:0] Wgt_4_399,input [WEIGHT_SIZE-1:0] Wgt_4_400,input [WEIGHT_SIZE-1:0] Wgt_4_401,input [WEIGHT_SIZE-1:0] Wgt_4_402,input [WEIGHT_SIZE-1:0] Wgt_4_403,input [WEIGHT_SIZE-1:0] Wgt_4_404,input [WEIGHT_SIZE-1:0] Wgt_4_405,input [WEIGHT_SIZE-1:0] Wgt_4_406,input [WEIGHT_SIZE-1:0] Wgt_4_407,input [WEIGHT_SIZE-1:0] Wgt_4_408,input [WEIGHT_SIZE-1:0] Wgt_4_409,input [WEIGHT_SIZE-1:0] Wgt_4_410,input [WEIGHT_SIZE-1:0] Wgt_4_411,input [WEIGHT_SIZE-1:0] Wgt_4_412,input [WEIGHT_SIZE-1:0] Wgt_4_413,input [WEIGHT_SIZE-1:0] Wgt_4_414,input [WEIGHT_SIZE-1:0] Wgt_4_415,input [WEIGHT_SIZE-1:0] Wgt_4_416,input [WEIGHT_SIZE-1:0] Wgt_4_417,input [WEIGHT_SIZE-1:0] Wgt_4_418,input [WEIGHT_SIZE-1:0] Wgt_4_419,input [WEIGHT_SIZE-1:0] Wgt_4_420,input [WEIGHT_SIZE-1:0] Wgt_4_421,input [WEIGHT_SIZE-1:0] Wgt_4_422,input [WEIGHT_SIZE-1:0] Wgt_4_423,input [WEIGHT_SIZE-1:0] Wgt_4_424,input [WEIGHT_SIZE-1:0] Wgt_4_425,input [WEIGHT_SIZE-1:0] Wgt_4_426,input [WEIGHT_SIZE-1:0] Wgt_4_427,input [WEIGHT_SIZE-1:0] Wgt_4_428,input [WEIGHT_SIZE-1:0] Wgt_4_429,input [WEIGHT_SIZE-1:0] Wgt_4_430,input [WEIGHT_SIZE-1:0] Wgt_4_431,input [WEIGHT_SIZE-1:0] Wgt_4_432,input [WEIGHT_SIZE-1:0] Wgt_4_433,input [WEIGHT_SIZE-1:0] Wgt_4_434,input [WEIGHT_SIZE-1:0] Wgt_4_435,input [WEIGHT_SIZE-1:0] Wgt_4_436,input [WEIGHT_SIZE-1:0] Wgt_4_437,input [WEIGHT_SIZE-1:0] Wgt_4_438,input [WEIGHT_SIZE-1:0] Wgt_4_439,input [WEIGHT_SIZE-1:0] Wgt_4_440,input [WEIGHT_SIZE-1:0] Wgt_4_441,input [WEIGHT_SIZE-1:0] Wgt_4_442,input [WEIGHT_SIZE-1:0] Wgt_4_443,input [WEIGHT_SIZE-1:0] Wgt_4_444,input [WEIGHT_SIZE-1:0] Wgt_4_445,input [WEIGHT_SIZE-1:0] Wgt_4_446,input [WEIGHT_SIZE-1:0] Wgt_4_447,input [WEIGHT_SIZE-1:0] Wgt_4_448,input [WEIGHT_SIZE-1:0] Wgt_4_449,input [WEIGHT_SIZE-1:0] Wgt_4_450,input [WEIGHT_SIZE-1:0] Wgt_4_451,input [WEIGHT_SIZE-1:0] Wgt_4_452,input [WEIGHT_SIZE-1:0] Wgt_4_453,input [WEIGHT_SIZE-1:0] Wgt_4_454,input [WEIGHT_SIZE-1:0] Wgt_4_455,input [WEIGHT_SIZE-1:0] Wgt_4_456,input [WEIGHT_SIZE-1:0] Wgt_4_457,input [WEIGHT_SIZE-1:0] Wgt_4_458,input [WEIGHT_SIZE-1:0] Wgt_4_459,input [WEIGHT_SIZE-1:0] Wgt_4_460,input [WEIGHT_SIZE-1:0] Wgt_4_461,input [WEIGHT_SIZE-1:0] Wgt_4_462,input [WEIGHT_SIZE-1:0] Wgt_4_463,input [WEIGHT_SIZE-1:0] Wgt_4_464,input [WEIGHT_SIZE-1:0] Wgt_4_465,input [WEIGHT_SIZE-1:0] Wgt_4_466,input [WEIGHT_SIZE-1:0] Wgt_4_467,input [WEIGHT_SIZE-1:0] Wgt_4_468,input [WEIGHT_SIZE-1:0] Wgt_4_469,input [WEIGHT_SIZE-1:0] Wgt_4_470,input [WEIGHT_SIZE-1:0] Wgt_4_471,input [WEIGHT_SIZE-1:0] Wgt_4_472,input [WEIGHT_SIZE-1:0] Wgt_4_473,input [WEIGHT_SIZE-1:0] Wgt_4_474,input [WEIGHT_SIZE-1:0] Wgt_4_475,input [WEIGHT_SIZE-1:0] Wgt_4_476,input [WEIGHT_SIZE-1:0] Wgt_4_477,input [WEIGHT_SIZE-1:0] Wgt_4_478,input [WEIGHT_SIZE-1:0] Wgt_4_479,input [WEIGHT_SIZE-1:0] Wgt_4_480,input [WEIGHT_SIZE-1:0] Wgt_4_481,input [WEIGHT_SIZE-1:0] Wgt_4_482,input [WEIGHT_SIZE-1:0] Wgt_4_483,input [WEIGHT_SIZE-1:0] Wgt_4_484,input [WEIGHT_SIZE-1:0] Wgt_4_485,input [WEIGHT_SIZE-1:0] Wgt_4_486,input [WEIGHT_SIZE-1:0] Wgt_4_487,input [WEIGHT_SIZE-1:0] Wgt_4_488,input [WEIGHT_SIZE-1:0] Wgt_4_489,input [WEIGHT_SIZE-1:0] Wgt_4_490,input [WEIGHT_SIZE-1:0] Wgt_4_491,input [WEIGHT_SIZE-1:0] Wgt_4_492,input [WEIGHT_SIZE-1:0] Wgt_4_493,input [WEIGHT_SIZE-1:0] Wgt_4_494,input [WEIGHT_SIZE-1:0] Wgt_4_495,input [WEIGHT_SIZE-1:0] Wgt_4_496,input [WEIGHT_SIZE-1:0] Wgt_4_497,input [WEIGHT_SIZE-1:0] Wgt_4_498,input [WEIGHT_SIZE-1:0] Wgt_4_499,input [WEIGHT_SIZE-1:0] Wgt_4_500,input [WEIGHT_SIZE-1:0] Wgt_4_501,input [WEIGHT_SIZE-1:0] Wgt_4_502,input [WEIGHT_SIZE-1:0] Wgt_4_503,input [WEIGHT_SIZE-1:0] Wgt_4_504,input [WEIGHT_SIZE-1:0] Wgt_4_505,input [WEIGHT_SIZE-1:0] Wgt_4_506,input [WEIGHT_SIZE-1:0] Wgt_4_507,input [WEIGHT_SIZE-1:0] Wgt_4_508,input [WEIGHT_SIZE-1:0] Wgt_4_509,input [WEIGHT_SIZE-1:0] Wgt_4_510,input [WEIGHT_SIZE-1:0] Wgt_4_511,input [WEIGHT_SIZE-1:0] Wgt_4_512,input [WEIGHT_SIZE-1:0] Wgt_4_513,input [WEIGHT_SIZE-1:0] Wgt_4_514,input [WEIGHT_SIZE-1:0] Wgt_4_515,input [WEIGHT_SIZE-1:0] Wgt_4_516,input [WEIGHT_SIZE-1:0] Wgt_4_517,input [WEIGHT_SIZE-1:0] Wgt_4_518,input [WEIGHT_SIZE-1:0] Wgt_4_519,input [WEIGHT_SIZE-1:0] Wgt_4_520,input [WEIGHT_SIZE-1:0] Wgt_4_521,input [WEIGHT_SIZE-1:0] Wgt_4_522,input [WEIGHT_SIZE-1:0] Wgt_4_523,input [WEIGHT_SIZE-1:0] Wgt_4_524,input [WEIGHT_SIZE-1:0] Wgt_4_525,input [WEIGHT_SIZE-1:0] Wgt_4_526,input [WEIGHT_SIZE-1:0] Wgt_4_527,input [WEIGHT_SIZE-1:0] Wgt_4_528,input [WEIGHT_SIZE-1:0] Wgt_4_529,input [WEIGHT_SIZE-1:0] Wgt_4_530,input [WEIGHT_SIZE-1:0] Wgt_4_531,input [WEIGHT_SIZE-1:0] Wgt_4_532,input [WEIGHT_SIZE-1:0] Wgt_4_533,input [WEIGHT_SIZE-1:0] Wgt_4_534,input [WEIGHT_SIZE-1:0] Wgt_4_535,input [WEIGHT_SIZE-1:0] Wgt_4_536,input [WEIGHT_SIZE-1:0] Wgt_4_537,input [WEIGHT_SIZE-1:0] Wgt_4_538,input [WEIGHT_SIZE-1:0] Wgt_4_539,input [WEIGHT_SIZE-1:0] Wgt_4_540,input [WEIGHT_SIZE-1:0] Wgt_4_541,input [WEIGHT_SIZE-1:0] Wgt_4_542,input [WEIGHT_SIZE-1:0] Wgt_4_543,input [WEIGHT_SIZE-1:0] Wgt_4_544,input [WEIGHT_SIZE-1:0] Wgt_4_545,input [WEIGHT_SIZE-1:0] Wgt_4_546,input [WEIGHT_SIZE-1:0] Wgt_4_547,input [WEIGHT_SIZE-1:0] Wgt_4_548,input [WEIGHT_SIZE-1:0] Wgt_4_549,input [WEIGHT_SIZE-1:0] Wgt_4_550,input [WEIGHT_SIZE-1:0] Wgt_4_551,input [WEIGHT_SIZE-1:0] Wgt_4_552,input [WEIGHT_SIZE-1:0] Wgt_4_553,input [WEIGHT_SIZE-1:0] Wgt_4_554,input [WEIGHT_SIZE-1:0] Wgt_4_555,input [WEIGHT_SIZE-1:0] Wgt_4_556,input [WEIGHT_SIZE-1:0] Wgt_4_557,input [WEIGHT_SIZE-1:0] Wgt_4_558,input [WEIGHT_SIZE-1:0] Wgt_4_559,input [WEIGHT_SIZE-1:0] Wgt_4_560,input [WEIGHT_SIZE-1:0] Wgt_4_561,input [WEIGHT_SIZE-1:0] Wgt_4_562,input [WEIGHT_SIZE-1:0] Wgt_4_563,input [WEIGHT_SIZE-1:0] Wgt_4_564,input [WEIGHT_SIZE-1:0] Wgt_4_565,input [WEIGHT_SIZE-1:0] Wgt_4_566,input [WEIGHT_SIZE-1:0] Wgt_4_567,input [WEIGHT_SIZE-1:0] Wgt_4_568,input [WEIGHT_SIZE-1:0] Wgt_4_569,input [WEIGHT_SIZE-1:0] Wgt_4_570,input [WEIGHT_SIZE-1:0] Wgt_4_571,input [WEIGHT_SIZE-1:0] Wgt_4_572,input [WEIGHT_SIZE-1:0] Wgt_4_573,input [WEIGHT_SIZE-1:0] Wgt_4_574,input [WEIGHT_SIZE-1:0] Wgt_4_575,input [WEIGHT_SIZE-1:0] Wgt_4_576,input [WEIGHT_SIZE-1:0] Wgt_4_577,input [WEIGHT_SIZE-1:0] Wgt_4_578,input [WEIGHT_SIZE-1:0] Wgt_4_579,input [WEIGHT_SIZE-1:0] Wgt_4_580,input [WEIGHT_SIZE-1:0] Wgt_4_581,input [WEIGHT_SIZE-1:0] Wgt_4_582,input [WEIGHT_SIZE-1:0] Wgt_4_583,input [WEIGHT_SIZE-1:0] Wgt_4_584,input [WEIGHT_SIZE-1:0] Wgt_4_585,input [WEIGHT_SIZE-1:0] Wgt_4_586,input [WEIGHT_SIZE-1:0] Wgt_4_587,input [WEIGHT_SIZE-1:0] Wgt_4_588,input [WEIGHT_SIZE-1:0] Wgt_4_589,input [WEIGHT_SIZE-1:0] Wgt_4_590,input [WEIGHT_SIZE-1:0] Wgt_4_591,input [WEIGHT_SIZE-1:0] Wgt_4_592,input [WEIGHT_SIZE-1:0] Wgt_4_593,input [WEIGHT_SIZE-1:0] Wgt_4_594,input [WEIGHT_SIZE-1:0] Wgt_4_595,input [WEIGHT_SIZE-1:0] Wgt_4_596,input [WEIGHT_SIZE-1:0] Wgt_4_597,input [WEIGHT_SIZE-1:0] Wgt_4_598,input [WEIGHT_SIZE-1:0] Wgt_4_599,input [WEIGHT_SIZE-1:0] Wgt_4_600,input [WEIGHT_SIZE-1:0] Wgt_4_601,input [WEIGHT_SIZE-1:0] Wgt_4_602,input [WEIGHT_SIZE-1:0] Wgt_4_603,input [WEIGHT_SIZE-1:0] Wgt_4_604,input [WEIGHT_SIZE-1:0] Wgt_4_605,input [WEIGHT_SIZE-1:0] Wgt_4_606,input [WEIGHT_SIZE-1:0] Wgt_4_607,input [WEIGHT_SIZE-1:0] Wgt_4_608,input [WEIGHT_SIZE-1:0] Wgt_4_609,input [WEIGHT_SIZE-1:0] Wgt_4_610,input [WEIGHT_SIZE-1:0] Wgt_4_611,input [WEIGHT_SIZE-1:0] Wgt_4_612,input [WEIGHT_SIZE-1:0] Wgt_4_613,input [WEIGHT_SIZE-1:0] Wgt_4_614,input [WEIGHT_SIZE-1:0] Wgt_4_615,input [WEIGHT_SIZE-1:0] Wgt_4_616,input [WEIGHT_SIZE-1:0] Wgt_4_617,input [WEIGHT_SIZE-1:0] Wgt_4_618,input [WEIGHT_SIZE-1:0] Wgt_4_619,input [WEIGHT_SIZE-1:0] Wgt_4_620,input [WEIGHT_SIZE-1:0] Wgt_4_621,input [WEIGHT_SIZE-1:0] Wgt_4_622,input [WEIGHT_SIZE-1:0] Wgt_4_623,input [WEIGHT_SIZE-1:0] Wgt_4_624,input [WEIGHT_SIZE-1:0] Wgt_4_625,input [WEIGHT_SIZE-1:0] Wgt_4_626,input [WEIGHT_SIZE-1:0] Wgt_4_627,input [WEIGHT_SIZE-1:0] Wgt_4_628,input [WEIGHT_SIZE-1:0] Wgt_4_629,input [WEIGHT_SIZE-1:0] Wgt_4_630,input [WEIGHT_SIZE-1:0] Wgt_4_631,input [WEIGHT_SIZE-1:0] Wgt_4_632,input [WEIGHT_SIZE-1:0] Wgt_4_633,input [WEIGHT_SIZE-1:0] Wgt_4_634,input [WEIGHT_SIZE-1:0] Wgt_4_635,input [WEIGHT_SIZE-1:0] Wgt_4_636,input [WEIGHT_SIZE-1:0] Wgt_4_637,input [WEIGHT_SIZE-1:0] Wgt_4_638,input [WEIGHT_SIZE-1:0] Wgt_4_639,input [WEIGHT_SIZE-1:0] Wgt_4_640,input [WEIGHT_SIZE-1:0] Wgt_4_641,input [WEIGHT_SIZE-1:0] Wgt_4_642,input [WEIGHT_SIZE-1:0] Wgt_4_643,input [WEIGHT_SIZE-1:0] Wgt_4_644,input [WEIGHT_SIZE-1:0] Wgt_4_645,input [WEIGHT_SIZE-1:0] Wgt_4_646,input [WEIGHT_SIZE-1:0] Wgt_4_647,input [WEIGHT_SIZE-1:0] Wgt_4_648,input [WEIGHT_SIZE-1:0] Wgt_4_649,input [WEIGHT_SIZE-1:0] Wgt_4_650,input [WEIGHT_SIZE-1:0] Wgt_4_651,input [WEIGHT_SIZE-1:0] Wgt_4_652,input [WEIGHT_SIZE-1:0] Wgt_4_653,input [WEIGHT_SIZE-1:0] Wgt_4_654,input [WEIGHT_SIZE-1:0] Wgt_4_655,input [WEIGHT_SIZE-1:0] Wgt_4_656,input [WEIGHT_SIZE-1:0] Wgt_4_657,input [WEIGHT_SIZE-1:0] Wgt_4_658,input [WEIGHT_SIZE-1:0] Wgt_4_659,input [WEIGHT_SIZE-1:0] Wgt_4_660,input [WEIGHT_SIZE-1:0] Wgt_4_661,input [WEIGHT_SIZE-1:0] Wgt_4_662,input [WEIGHT_SIZE-1:0] Wgt_4_663,input [WEIGHT_SIZE-1:0] Wgt_4_664,input [WEIGHT_SIZE-1:0] Wgt_4_665,input [WEIGHT_SIZE-1:0] Wgt_4_666,input [WEIGHT_SIZE-1:0] Wgt_4_667,input [WEIGHT_SIZE-1:0] Wgt_4_668,input [WEIGHT_SIZE-1:0] Wgt_4_669,input [WEIGHT_SIZE-1:0] Wgt_4_670,input [WEIGHT_SIZE-1:0] Wgt_4_671,input [WEIGHT_SIZE-1:0] Wgt_4_672,input [WEIGHT_SIZE-1:0] Wgt_4_673,input [WEIGHT_SIZE-1:0] Wgt_4_674,input [WEIGHT_SIZE-1:0] Wgt_4_675,input [WEIGHT_SIZE-1:0] Wgt_4_676,input [WEIGHT_SIZE-1:0] Wgt_4_677,input [WEIGHT_SIZE-1:0] Wgt_4_678,input [WEIGHT_SIZE-1:0] Wgt_4_679,input [WEIGHT_SIZE-1:0] Wgt_4_680,input [WEIGHT_SIZE-1:0] Wgt_4_681,input [WEIGHT_SIZE-1:0] Wgt_4_682,input [WEIGHT_SIZE-1:0] Wgt_4_683,input [WEIGHT_SIZE-1:0] Wgt_4_684,input [WEIGHT_SIZE-1:0] Wgt_4_685,input [WEIGHT_SIZE-1:0] Wgt_4_686,input [WEIGHT_SIZE-1:0] Wgt_4_687,input [WEIGHT_SIZE-1:0] Wgt_4_688,input [WEIGHT_SIZE-1:0] Wgt_4_689,input [WEIGHT_SIZE-1:0] Wgt_4_690,input [WEIGHT_SIZE-1:0] Wgt_4_691,input [WEIGHT_SIZE-1:0] Wgt_4_692,input [WEIGHT_SIZE-1:0] Wgt_4_693,input [WEIGHT_SIZE-1:0] Wgt_4_694,input [WEIGHT_SIZE-1:0] Wgt_4_695,input [WEIGHT_SIZE-1:0] Wgt_4_696,input [WEIGHT_SIZE-1:0] Wgt_4_697,input [WEIGHT_SIZE-1:0] Wgt_4_698,input [WEIGHT_SIZE-1:0] Wgt_4_699,input [WEIGHT_SIZE-1:0] Wgt_4_700,input [WEIGHT_SIZE-1:0] Wgt_4_701,input [WEIGHT_SIZE-1:0] Wgt_4_702,input [WEIGHT_SIZE-1:0] Wgt_4_703,input [WEIGHT_SIZE-1:0] Wgt_4_704,input [WEIGHT_SIZE-1:0] Wgt_4_705,input [WEIGHT_SIZE-1:0] Wgt_4_706,input [WEIGHT_SIZE-1:0] Wgt_4_707,input [WEIGHT_SIZE-1:0] Wgt_4_708,input [WEIGHT_SIZE-1:0] Wgt_4_709,input [WEIGHT_SIZE-1:0] Wgt_4_710,input [WEIGHT_SIZE-1:0] Wgt_4_711,input [WEIGHT_SIZE-1:0] Wgt_4_712,input [WEIGHT_SIZE-1:0] Wgt_4_713,input [WEIGHT_SIZE-1:0] Wgt_4_714,input [WEIGHT_SIZE-1:0] Wgt_4_715,input [WEIGHT_SIZE-1:0] Wgt_4_716,input [WEIGHT_SIZE-1:0] Wgt_4_717,input [WEIGHT_SIZE-1:0] Wgt_4_718,input [WEIGHT_SIZE-1:0] Wgt_4_719,input [WEIGHT_SIZE-1:0] Wgt_4_720,input [WEIGHT_SIZE-1:0] Wgt_4_721,input [WEIGHT_SIZE-1:0] Wgt_4_722,input [WEIGHT_SIZE-1:0] Wgt_4_723,input [WEIGHT_SIZE-1:0] Wgt_4_724,input [WEIGHT_SIZE-1:0] Wgt_4_725,input [WEIGHT_SIZE-1:0] Wgt_4_726,input [WEIGHT_SIZE-1:0] Wgt_4_727,input [WEIGHT_SIZE-1:0] Wgt_4_728,input [WEIGHT_SIZE-1:0] Wgt_4_729,input [WEIGHT_SIZE-1:0] Wgt_4_730,input [WEIGHT_SIZE-1:0] Wgt_4_731,input [WEIGHT_SIZE-1:0] Wgt_4_732,input [WEIGHT_SIZE-1:0] Wgt_4_733,input [WEIGHT_SIZE-1:0] Wgt_4_734,input [WEIGHT_SIZE-1:0] Wgt_4_735,input [WEIGHT_SIZE-1:0] Wgt_4_736,input [WEIGHT_SIZE-1:0] Wgt_4_737,input [WEIGHT_SIZE-1:0] Wgt_4_738,input [WEIGHT_SIZE-1:0] Wgt_4_739,input [WEIGHT_SIZE-1:0] Wgt_4_740,input [WEIGHT_SIZE-1:0] Wgt_4_741,input [WEIGHT_SIZE-1:0] Wgt_4_742,input [WEIGHT_SIZE-1:0] Wgt_4_743,input [WEIGHT_SIZE-1:0] Wgt_4_744,input [WEIGHT_SIZE-1:0] Wgt_4_745,input [WEIGHT_SIZE-1:0] Wgt_4_746,input [WEIGHT_SIZE-1:0] Wgt_4_747,input [WEIGHT_SIZE-1:0] Wgt_4_748,input [WEIGHT_SIZE-1:0] Wgt_4_749,input [WEIGHT_SIZE-1:0] Wgt_4_750,input [WEIGHT_SIZE-1:0] Wgt_4_751,input [WEIGHT_SIZE-1:0] Wgt_4_752,input [WEIGHT_SIZE-1:0] Wgt_4_753,input [WEIGHT_SIZE-1:0] Wgt_4_754,input [WEIGHT_SIZE-1:0] Wgt_4_755,input [WEIGHT_SIZE-1:0] Wgt_4_756,input [WEIGHT_SIZE-1:0] Wgt_4_757,input [WEIGHT_SIZE-1:0] Wgt_4_758,input [WEIGHT_SIZE-1:0] Wgt_4_759,input [WEIGHT_SIZE-1:0] Wgt_4_760,input [WEIGHT_SIZE-1:0] Wgt_4_761,input [WEIGHT_SIZE-1:0] Wgt_4_762,input [WEIGHT_SIZE-1:0] Wgt_4_763,input [WEIGHT_SIZE-1:0] Wgt_4_764,input [WEIGHT_SIZE-1:0] Wgt_4_765,input [WEIGHT_SIZE-1:0] Wgt_4_766,input [WEIGHT_SIZE-1:0] Wgt_4_767,input [WEIGHT_SIZE-1:0] Wgt_4_768,input [WEIGHT_SIZE-1:0] Wgt_4_769,input [WEIGHT_SIZE-1:0] Wgt_4_770,input [WEIGHT_SIZE-1:0] Wgt_4_771,input [WEIGHT_SIZE-1:0] Wgt_4_772,input [WEIGHT_SIZE-1:0] Wgt_4_773,input [WEIGHT_SIZE-1:0] Wgt_4_774,input [WEIGHT_SIZE-1:0] Wgt_4_775,input [WEIGHT_SIZE-1:0] Wgt_4_776,input [WEIGHT_SIZE-1:0] Wgt_4_777,input [WEIGHT_SIZE-1:0] Wgt_4_778,input [WEIGHT_SIZE-1:0] Wgt_4_779,input [WEIGHT_SIZE-1:0] Wgt_4_780,input [WEIGHT_SIZE-1:0] Wgt_4_781,input [WEIGHT_SIZE-1:0] Wgt_4_782,input [WEIGHT_SIZE-1:0] Wgt_4_783,input [WEIGHT_SIZE-1:0] Wgt_4_784,input [WEIGHT_SIZE-1:0] Wgt_5_0,input [WEIGHT_SIZE-1:0] Wgt_5_1,input [WEIGHT_SIZE-1:0] Wgt_5_2,input [WEIGHT_SIZE-1:0] Wgt_5_3,input [WEIGHT_SIZE-1:0] Wgt_5_4,input [WEIGHT_SIZE-1:0] Wgt_5_5,input [WEIGHT_SIZE-1:0] Wgt_5_6,input [WEIGHT_SIZE-1:0] Wgt_5_7,input [WEIGHT_SIZE-1:0] Wgt_5_8,input [WEIGHT_SIZE-1:0] Wgt_5_9,input [WEIGHT_SIZE-1:0] Wgt_5_10,input [WEIGHT_SIZE-1:0] Wgt_5_11,input [WEIGHT_SIZE-1:0] Wgt_5_12,input [WEIGHT_SIZE-1:0] Wgt_5_13,input [WEIGHT_SIZE-1:0] Wgt_5_14,input [WEIGHT_SIZE-1:0] Wgt_5_15,input [WEIGHT_SIZE-1:0] Wgt_5_16,input [WEIGHT_SIZE-1:0] Wgt_5_17,input [WEIGHT_SIZE-1:0] Wgt_5_18,input [WEIGHT_SIZE-1:0] Wgt_5_19,input [WEIGHT_SIZE-1:0] Wgt_5_20,input [WEIGHT_SIZE-1:0] Wgt_5_21,input [WEIGHT_SIZE-1:0] Wgt_5_22,input [WEIGHT_SIZE-1:0] Wgt_5_23,input [WEIGHT_SIZE-1:0] Wgt_5_24,input [WEIGHT_SIZE-1:0] Wgt_5_25,input [WEIGHT_SIZE-1:0] Wgt_5_26,input [WEIGHT_SIZE-1:0] Wgt_5_27,input [WEIGHT_SIZE-1:0] Wgt_5_28,input [WEIGHT_SIZE-1:0] Wgt_5_29,input [WEIGHT_SIZE-1:0] Wgt_5_30,input [WEIGHT_SIZE-1:0] Wgt_5_31,input [WEIGHT_SIZE-1:0] Wgt_5_32,input [WEIGHT_SIZE-1:0] Wgt_5_33,input [WEIGHT_SIZE-1:0] Wgt_5_34,input [WEIGHT_SIZE-1:0] Wgt_5_35,input [WEIGHT_SIZE-1:0] Wgt_5_36,input [WEIGHT_SIZE-1:0] Wgt_5_37,input [WEIGHT_SIZE-1:0] Wgt_5_38,input [WEIGHT_SIZE-1:0] Wgt_5_39,input [WEIGHT_SIZE-1:0] Wgt_5_40,input [WEIGHT_SIZE-1:0] Wgt_5_41,input [WEIGHT_SIZE-1:0] Wgt_5_42,input [WEIGHT_SIZE-1:0] Wgt_5_43,input [WEIGHT_SIZE-1:0] Wgt_5_44,input [WEIGHT_SIZE-1:0] Wgt_5_45,input [WEIGHT_SIZE-1:0] Wgt_5_46,input [WEIGHT_SIZE-1:0] Wgt_5_47,input [WEIGHT_SIZE-1:0] Wgt_5_48,input [WEIGHT_SIZE-1:0] Wgt_5_49,input [WEIGHT_SIZE-1:0] Wgt_5_50,input [WEIGHT_SIZE-1:0] Wgt_5_51,input [WEIGHT_SIZE-1:0] Wgt_5_52,input [WEIGHT_SIZE-1:0] Wgt_5_53,input [WEIGHT_SIZE-1:0] Wgt_5_54,input [WEIGHT_SIZE-1:0] Wgt_5_55,input [WEIGHT_SIZE-1:0] Wgt_5_56,input [WEIGHT_SIZE-1:0] Wgt_5_57,input [WEIGHT_SIZE-1:0] Wgt_5_58,input [WEIGHT_SIZE-1:0] Wgt_5_59,input [WEIGHT_SIZE-1:0] Wgt_5_60,input [WEIGHT_SIZE-1:0] Wgt_5_61,input [WEIGHT_SIZE-1:0] Wgt_5_62,input [WEIGHT_SIZE-1:0] Wgt_5_63,input [WEIGHT_SIZE-1:0] Wgt_5_64,input [WEIGHT_SIZE-1:0] Wgt_5_65,input [WEIGHT_SIZE-1:0] Wgt_5_66,input [WEIGHT_SIZE-1:0] Wgt_5_67,input [WEIGHT_SIZE-1:0] Wgt_5_68,input [WEIGHT_SIZE-1:0] Wgt_5_69,input [WEIGHT_SIZE-1:0] Wgt_5_70,input [WEIGHT_SIZE-1:0] Wgt_5_71,input [WEIGHT_SIZE-1:0] Wgt_5_72,input [WEIGHT_SIZE-1:0] Wgt_5_73,input [WEIGHT_SIZE-1:0] Wgt_5_74,input [WEIGHT_SIZE-1:0] Wgt_5_75,input [WEIGHT_SIZE-1:0] Wgt_5_76,input [WEIGHT_SIZE-1:0] Wgt_5_77,input [WEIGHT_SIZE-1:0] Wgt_5_78,input [WEIGHT_SIZE-1:0] Wgt_5_79,input [WEIGHT_SIZE-1:0] Wgt_5_80,input [WEIGHT_SIZE-1:0] Wgt_5_81,input [WEIGHT_SIZE-1:0] Wgt_5_82,input [WEIGHT_SIZE-1:0] Wgt_5_83,input [WEIGHT_SIZE-1:0] Wgt_5_84,input [WEIGHT_SIZE-1:0] Wgt_5_85,input [WEIGHT_SIZE-1:0] Wgt_5_86,input [WEIGHT_SIZE-1:0] Wgt_5_87,input [WEIGHT_SIZE-1:0] Wgt_5_88,input [WEIGHT_SIZE-1:0] Wgt_5_89,input [WEIGHT_SIZE-1:0] Wgt_5_90,input [WEIGHT_SIZE-1:0] Wgt_5_91,input [WEIGHT_SIZE-1:0] Wgt_5_92,input [WEIGHT_SIZE-1:0] Wgt_5_93,input [WEIGHT_SIZE-1:0] Wgt_5_94,input [WEIGHT_SIZE-1:0] Wgt_5_95,input [WEIGHT_SIZE-1:0] Wgt_5_96,input [WEIGHT_SIZE-1:0] Wgt_5_97,input [WEIGHT_SIZE-1:0] Wgt_5_98,input [WEIGHT_SIZE-1:0] Wgt_5_99,input [WEIGHT_SIZE-1:0] Wgt_5_100,input [WEIGHT_SIZE-1:0] Wgt_5_101,input [WEIGHT_SIZE-1:0] Wgt_5_102,input [WEIGHT_SIZE-1:0] Wgt_5_103,input [WEIGHT_SIZE-1:0] Wgt_5_104,input [WEIGHT_SIZE-1:0] Wgt_5_105,input [WEIGHT_SIZE-1:0] Wgt_5_106,input [WEIGHT_SIZE-1:0] Wgt_5_107,input [WEIGHT_SIZE-1:0] Wgt_5_108,input [WEIGHT_SIZE-1:0] Wgt_5_109,input [WEIGHT_SIZE-1:0] Wgt_5_110,input [WEIGHT_SIZE-1:0] Wgt_5_111,input [WEIGHT_SIZE-1:0] Wgt_5_112,input [WEIGHT_SIZE-1:0] Wgt_5_113,input [WEIGHT_SIZE-1:0] Wgt_5_114,input [WEIGHT_SIZE-1:0] Wgt_5_115,input [WEIGHT_SIZE-1:0] Wgt_5_116,input [WEIGHT_SIZE-1:0] Wgt_5_117,input [WEIGHT_SIZE-1:0] Wgt_5_118,input [WEIGHT_SIZE-1:0] Wgt_5_119,input [WEIGHT_SIZE-1:0] Wgt_5_120,input [WEIGHT_SIZE-1:0] Wgt_5_121,input [WEIGHT_SIZE-1:0] Wgt_5_122,input [WEIGHT_SIZE-1:0] Wgt_5_123,input [WEIGHT_SIZE-1:0] Wgt_5_124,input [WEIGHT_SIZE-1:0] Wgt_5_125,input [WEIGHT_SIZE-1:0] Wgt_5_126,input [WEIGHT_SIZE-1:0] Wgt_5_127,input [WEIGHT_SIZE-1:0] Wgt_5_128,input [WEIGHT_SIZE-1:0] Wgt_5_129,input [WEIGHT_SIZE-1:0] Wgt_5_130,input [WEIGHT_SIZE-1:0] Wgt_5_131,input [WEIGHT_SIZE-1:0] Wgt_5_132,input [WEIGHT_SIZE-1:0] Wgt_5_133,input [WEIGHT_SIZE-1:0] Wgt_5_134,input [WEIGHT_SIZE-1:0] Wgt_5_135,input [WEIGHT_SIZE-1:0] Wgt_5_136,input [WEIGHT_SIZE-1:0] Wgt_5_137,input [WEIGHT_SIZE-1:0] Wgt_5_138,input [WEIGHT_SIZE-1:0] Wgt_5_139,input [WEIGHT_SIZE-1:0] Wgt_5_140,input [WEIGHT_SIZE-1:0] Wgt_5_141,input [WEIGHT_SIZE-1:0] Wgt_5_142,input [WEIGHT_SIZE-1:0] Wgt_5_143,input [WEIGHT_SIZE-1:0] Wgt_5_144,input [WEIGHT_SIZE-1:0] Wgt_5_145,input [WEIGHT_SIZE-1:0] Wgt_5_146,input [WEIGHT_SIZE-1:0] Wgt_5_147,input [WEIGHT_SIZE-1:0] Wgt_5_148,input [WEIGHT_SIZE-1:0] Wgt_5_149,input [WEIGHT_SIZE-1:0] Wgt_5_150,input [WEIGHT_SIZE-1:0] Wgt_5_151,input [WEIGHT_SIZE-1:0] Wgt_5_152,input [WEIGHT_SIZE-1:0] Wgt_5_153,input [WEIGHT_SIZE-1:0] Wgt_5_154,input [WEIGHT_SIZE-1:0] Wgt_5_155,input [WEIGHT_SIZE-1:0] Wgt_5_156,input [WEIGHT_SIZE-1:0] Wgt_5_157,input [WEIGHT_SIZE-1:0] Wgt_5_158,input [WEIGHT_SIZE-1:0] Wgt_5_159,input [WEIGHT_SIZE-1:0] Wgt_5_160,input [WEIGHT_SIZE-1:0] Wgt_5_161,input [WEIGHT_SIZE-1:0] Wgt_5_162,input [WEIGHT_SIZE-1:0] Wgt_5_163,input [WEIGHT_SIZE-1:0] Wgt_5_164,input [WEIGHT_SIZE-1:0] Wgt_5_165,input [WEIGHT_SIZE-1:0] Wgt_5_166,input [WEIGHT_SIZE-1:0] Wgt_5_167,input [WEIGHT_SIZE-1:0] Wgt_5_168,input [WEIGHT_SIZE-1:0] Wgt_5_169,input [WEIGHT_SIZE-1:0] Wgt_5_170,input [WEIGHT_SIZE-1:0] Wgt_5_171,input [WEIGHT_SIZE-1:0] Wgt_5_172,input [WEIGHT_SIZE-1:0] Wgt_5_173,input [WEIGHT_SIZE-1:0] Wgt_5_174,input [WEIGHT_SIZE-1:0] Wgt_5_175,input [WEIGHT_SIZE-1:0] Wgt_5_176,input [WEIGHT_SIZE-1:0] Wgt_5_177,input [WEIGHT_SIZE-1:0] Wgt_5_178,input [WEIGHT_SIZE-1:0] Wgt_5_179,input [WEIGHT_SIZE-1:0] Wgt_5_180,input [WEIGHT_SIZE-1:0] Wgt_5_181,input [WEIGHT_SIZE-1:0] Wgt_5_182,input [WEIGHT_SIZE-1:0] Wgt_5_183,input [WEIGHT_SIZE-1:0] Wgt_5_184,input [WEIGHT_SIZE-1:0] Wgt_5_185,input [WEIGHT_SIZE-1:0] Wgt_5_186,input [WEIGHT_SIZE-1:0] Wgt_5_187,input [WEIGHT_SIZE-1:0] Wgt_5_188,input [WEIGHT_SIZE-1:0] Wgt_5_189,input [WEIGHT_SIZE-1:0] Wgt_5_190,input [WEIGHT_SIZE-1:0] Wgt_5_191,input [WEIGHT_SIZE-1:0] Wgt_5_192,input [WEIGHT_SIZE-1:0] Wgt_5_193,input [WEIGHT_SIZE-1:0] Wgt_5_194,input [WEIGHT_SIZE-1:0] Wgt_5_195,input [WEIGHT_SIZE-1:0] Wgt_5_196,input [WEIGHT_SIZE-1:0] Wgt_5_197,input [WEIGHT_SIZE-1:0] Wgt_5_198,input [WEIGHT_SIZE-1:0] Wgt_5_199,input [WEIGHT_SIZE-1:0] Wgt_5_200,input [WEIGHT_SIZE-1:0] Wgt_5_201,input [WEIGHT_SIZE-1:0] Wgt_5_202,input [WEIGHT_SIZE-1:0] Wgt_5_203,input [WEIGHT_SIZE-1:0] Wgt_5_204,input [WEIGHT_SIZE-1:0] Wgt_5_205,input [WEIGHT_SIZE-1:0] Wgt_5_206,input [WEIGHT_SIZE-1:0] Wgt_5_207,input [WEIGHT_SIZE-1:0] Wgt_5_208,input [WEIGHT_SIZE-1:0] Wgt_5_209,input [WEIGHT_SIZE-1:0] Wgt_5_210,input [WEIGHT_SIZE-1:0] Wgt_5_211,input [WEIGHT_SIZE-1:0] Wgt_5_212,input [WEIGHT_SIZE-1:0] Wgt_5_213,input [WEIGHT_SIZE-1:0] Wgt_5_214,input [WEIGHT_SIZE-1:0] Wgt_5_215,input [WEIGHT_SIZE-1:0] Wgt_5_216,input [WEIGHT_SIZE-1:0] Wgt_5_217,input [WEIGHT_SIZE-1:0] Wgt_5_218,input [WEIGHT_SIZE-1:0] Wgt_5_219,input [WEIGHT_SIZE-1:0] Wgt_5_220,input [WEIGHT_SIZE-1:0] Wgt_5_221,input [WEIGHT_SIZE-1:0] Wgt_5_222,input [WEIGHT_SIZE-1:0] Wgt_5_223,input [WEIGHT_SIZE-1:0] Wgt_5_224,input [WEIGHT_SIZE-1:0] Wgt_5_225,input [WEIGHT_SIZE-1:0] Wgt_5_226,input [WEIGHT_SIZE-1:0] Wgt_5_227,input [WEIGHT_SIZE-1:0] Wgt_5_228,input [WEIGHT_SIZE-1:0] Wgt_5_229,input [WEIGHT_SIZE-1:0] Wgt_5_230,input [WEIGHT_SIZE-1:0] Wgt_5_231,input [WEIGHT_SIZE-1:0] Wgt_5_232,input [WEIGHT_SIZE-1:0] Wgt_5_233,input [WEIGHT_SIZE-1:0] Wgt_5_234,input [WEIGHT_SIZE-1:0] Wgt_5_235,input [WEIGHT_SIZE-1:0] Wgt_5_236,input [WEIGHT_SIZE-1:0] Wgt_5_237,input [WEIGHT_SIZE-1:0] Wgt_5_238,input [WEIGHT_SIZE-1:0] Wgt_5_239,input [WEIGHT_SIZE-1:0] Wgt_5_240,input [WEIGHT_SIZE-1:0] Wgt_5_241,input [WEIGHT_SIZE-1:0] Wgt_5_242,input [WEIGHT_SIZE-1:0] Wgt_5_243,input [WEIGHT_SIZE-1:0] Wgt_5_244,input [WEIGHT_SIZE-1:0] Wgt_5_245,input [WEIGHT_SIZE-1:0] Wgt_5_246,input [WEIGHT_SIZE-1:0] Wgt_5_247,input [WEIGHT_SIZE-1:0] Wgt_5_248,input [WEIGHT_SIZE-1:0] Wgt_5_249,input [WEIGHT_SIZE-1:0] Wgt_5_250,input [WEIGHT_SIZE-1:0] Wgt_5_251,input [WEIGHT_SIZE-1:0] Wgt_5_252,input [WEIGHT_SIZE-1:0] Wgt_5_253,input [WEIGHT_SIZE-1:0] Wgt_5_254,input [WEIGHT_SIZE-1:0] Wgt_5_255,input [WEIGHT_SIZE-1:0] Wgt_5_256,input [WEIGHT_SIZE-1:0] Wgt_5_257,input [WEIGHT_SIZE-1:0] Wgt_5_258,input [WEIGHT_SIZE-1:0] Wgt_5_259,input [WEIGHT_SIZE-1:0] Wgt_5_260,input [WEIGHT_SIZE-1:0] Wgt_5_261,input [WEIGHT_SIZE-1:0] Wgt_5_262,input [WEIGHT_SIZE-1:0] Wgt_5_263,input [WEIGHT_SIZE-1:0] Wgt_5_264,input [WEIGHT_SIZE-1:0] Wgt_5_265,input [WEIGHT_SIZE-1:0] Wgt_5_266,input [WEIGHT_SIZE-1:0] Wgt_5_267,input [WEIGHT_SIZE-1:0] Wgt_5_268,input [WEIGHT_SIZE-1:0] Wgt_5_269,input [WEIGHT_SIZE-1:0] Wgt_5_270,input [WEIGHT_SIZE-1:0] Wgt_5_271,input [WEIGHT_SIZE-1:0] Wgt_5_272,input [WEIGHT_SIZE-1:0] Wgt_5_273,input [WEIGHT_SIZE-1:0] Wgt_5_274,input [WEIGHT_SIZE-1:0] Wgt_5_275,input [WEIGHT_SIZE-1:0] Wgt_5_276,input [WEIGHT_SIZE-1:0] Wgt_5_277,input [WEIGHT_SIZE-1:0] Wgt_5_278,input [WEIGHT_SIZE-1:0] Wgt_5_279,input [WEIGHT_SIZE-1:0] Wgt_5_280,input [WEIGHT_SIZE-1:0] Wgt_5_281,input [WEIGHT_SIZE-1:0] Wgt_5_282,input [WEIGHT_SIZE-1:0] Wgt_5_283,input [WEIGHT_SIZE-1:0] Wgt_5_284,input [WEIGHT_SIZE-1:0] Wgt_5_285,input [WEIGHT_SIZE-1:0] Wgt_5_286,input [WEIGHT_SIZE-1:0] Wgt_5_287,input [WEIGHT_SIZE-1:0] Wgt_5_288,input [WEIGHT_SIZE-1:0] Wgt_5_289,input [WEIGHT_SIZE-1:0] Wgt_5_290,input [WEIGHT_SIZE-1:0] Wgt_5_291,input [WEIGHT_SIZE-1:0] Wgt_5_292,input [WEIGHT_SIZE-1:0] Wgt_5_293,input [WEIGHT_SIZE-1:0] Wgt_5_294,input [WEIGHT_SIZE-1:0] Wgt_5_295,input [WEIGHT_SIZE-1:0] Wgt_5_296,input [WEIGHT_SIZE-1:0] Wgt_5_297,input [WEIGHT_SIZE-1:0] Wgt_5_298,input [WEIGHT_SIZE-1:0] Wgt_5_299,input [WEIGHT_SIZE-1:0] Wgt_5_300,input [WEIGHT_SIZE-1:0] Wgt_5_301,input [WEIGHT_SIZE-1:0] Wgt_5_302,input [WEIGHT_SIZE-1:0] Wgt_5_303,input [WEIGHT_SIZE-1:0] Wgt_5_304,input [WEIGHT_SIZE-1:0] Wgt_5_305,input [WEIGHT_SIZE-1:0] Wgt_5_306,input [WEIGHT_SIZE-1:0] Wgt_5_307,input [WEIGHT_SIZE-1:0] Wgt_5_308,input [WEIGHT_SIZE-1:0] Wgt_5_309,input [WEIGHT_SIZE-1:0] Wgt_5_310,input [WEIGHT_SIZE-1:0] Wgt_5_311,input [WEIGHT_SIZE-1:0] Wgt_5_312,input [WEIGHT_SIZE-1:0] Wgt_5_313,input [WEIGHT_SIZE-1:0] Wgt_5_314,input [WEIGHT_SIZE-1:0] Wgt_5_315,input [WEIGHT_SIZE-1:0] Wgt_5_316,input [WEIGHT_SIZE-1:0] Wgt_5_317,input [WEIGHT_SIZE-1:0] Wgt_5_318,input [WEIGHT_SIZE-1:0] Wgt_5_319,input [WEIGHT_SIZE-1:0] Wgt_5_320,input [WEIGHT_SIZE-1:0] Wgt_5_321,input [WEIGHT_SIZE-1:0] Wgt_5_322,input [WEIGHT_SIZE-1:0] Wgt_5_323,input [WEIGHT_SIZE-1:0] Wgt_5_324,input [WEIGHT_SIZE-1:0] Wgt_5_325,input [WEIGHT_SIZE-1:0] Wgt_5_326,input [WEIGHT_SIZE-1:0] Wgt_5_327,input [WEIGHT_SIZE-1:0] Wgt_5_328,input [WEIGHT_SIZE-1:0] Wgt_5_329,input [WEIGHT_SIZE-1:0] Wgt_5_330,input [WEIGHT_SIZE-1:0] Wgt_5_331,input [WEIGHT_SIZE-1:0] Wgt_5_332,input [WEIGHT_SIZE-1:0] Wgt_5_333,input [WEIGHT_SIZE-1:0] Wgt_5_334,input [WEIGHT_SIZE-1:0] Wgt_5_335,input [WEIGHT_SIZE-1:0] Wgt_5_336,input [WEIGHT_SIZE-1:0] Wgt_5_337,input [WEIGHT_SIZE-1:0] Wgt_5_338,input [WEIGHT_SIZE-1:0] Wgt_5_339,input [WEIGHT_SIZE-1:0] Wgt_5_340,input [WEIGHT_SIZE-1:0] Wgt_5_341,input [WEIGHT_SIZE-1:0] Wgt_5_342,input [WEIGHT_SIZE-1:0] Wgt_5_343,input [WEIGHT_SIZE-1:0] Wgt_5_344,input [WEIGHT_SIZE-1:0] Wgt_5_345,input [WEIGHT_SIZE-1:0] Wgt_5_346,input [WEIGHT_SIZE-1:0] Wgt_5_347,input [WEIGHT_SIZE-1:0] Wgt_5_348,input [WEIGHT_SIZE-1:0] Wgt_5_349,input [WEIGHT_SIZE-1:0] Wgt_5_350,input [WEIGHT_SIZE-1:0] Wgt_5_351,input [WEIGHT_SIZE-1:0] Wgt_5_352,input [WEIGHT_SIZE-1:0] Wgt_5_353,input [WEIGHT_SIZE-1:0] Wgt_5_354,input [WEIGHT_SIZE-1:0] Wgt_5_355,input [WEIGHT_SIZE-1:0] Wgt_5_356,input [WEIGHT_SIZE-1:0] Wgt_5_357,input [WEIGHT_SIZE-1:0] Wgt_5_358,input [WEIGHT_SIZE-1:0] Wgt_5_359,input [WEIGHT_SIZE-1:0] Wgt_5_360,input [WEIGHT_SIZE-1:0] Wgt_5_361,input [WEIGHT_SIZE-1:0] Wgt_5_362,input [WEIGHT_SIZE-1:0] Wgt_5_363,input [WEIGHT_SIZE-1:0] Wgt_5_364,input [WEIGHT_SIZE-1:0] Wgt_5_365,input [WEIGHT_SIZE-1:0] Wgt_5_366,input [WEIGHT_SIZE-1:0] Wgt_5_367,input [WEIGHT_SIZE-1:0] Wgt_5_368,input [WEIGHT_SIZE-1:0] Wgt_5_369,input [WEIGHT_SIZE-1:0] Wgt_5_370,input [WEIGHT_SIZE-1:0] Wgt_5_371,input [WEIGHT_SIZE-1:0] Wgt_5_372,input [WEIGHT_SIZE-1:0] Wgt_5_373,input [WEIGHT_SIZE-1:0] Wgt_5_374,input [WEIGHT_SIZE-1:0] Wgt_5_375,input [WEIGHT_SIZE-1:0] Wgt_5_376,input [WEIGHT_SIZE-1:0] Wgt_5_377,input [WEIGHT_SIZE-1:0] Wgt_5_378,input [WEIGHT_SIZE-1:0] Wgt_5_379,input [WEIGHT_SIZE-1:0] Wgt_5_380,input [WEIGHT_SIZE-1:0] Wgt_5_381,input [WEIGHT_SIZE-1:0] Wgt_5_382,input [WEIGHT_SIZE-1:0] Wgt_5_383,input [WEIGHT_SIZE-1:0] Wgt_5_384,input [WEIGHT_SIZE-1:0] Wgt_5_385,input [WEIGHT_SIZE-1:0] Wgt_5_386,input [WEIGHT_SIZE-1:0] Wgt_5_387,input [WEIGHT_SIZE-1:0] Wgt_5_388,input [WEIGHT_SIZE-1:0] Wgt_5_389,input [WEIGHT_SIZE-1:0] Wgt_5_390,input [WEIGHT_SIZE-1:0] Wgt_5_391,input [WEIGHT_SIZE-1:0] Wgt_5_392,input [WEIGHT_SIZE-1:0] Wgt_5_393,input [WEIGHT_SIZE-1:0] Wgt_5_394,input [WEIGHT_SIZE-1:0] Wgt_5_395,input [WEIGHT_SIZE-1:0] Wgt_5_396,input [WEIGHT_SIZE-1:0] Wgt_5_397,input [WEIGHT_SIZE-1:0] Wgt_5_398,input [WEIGHT_SIZE-1:0] Wgt_5_399,input [WEIGHT_SIZE-1:0] Wgt_5_400,input [WEIGHT_SIZE-1:0] Wgt_5_401,input [WEIGHT_SIZE-1:0] Wgt_5_402,input [WEIGHT_SIZE-1:0] Wgt_5_403,input [WEIGHT_SIZE-1:0] Wgt_5_404,input [WEIGHT_SIZE-1:0] Wgt_5_405,input [WEIGHT_SIZE-1:0] Wgt_5_406,input [WEIGHT_SIZE-1:0] Wgt_5_407,input [WEIGHT_SIZE-1:0] Wgt_5_408,input [WEIGHT_SIZE-1:0] Wgt_5_409,input [WEIGHT_SIZE-1:0] Wgt_5_410,input [WEIGHT_SIZE-1:0] Wgt_5_411,input [WEIGHT_SIZE-1:0] Wgt_5_412,input [WEIGHT_SIZE-1:0] Wgt_5_413,input [WEIGHT_SIZE-1:0] Wgt_5_414,input [WEIGHT_SIZE-1:0] Wgt_5_415,input [WEIGHT_SIZE-1:0] Wgt_5_416,input [WEIGHT_SIZE-1:0] Wgt_5_417,input [WEIGHT_SIZE-1:0] Wgt_5_418,input [WEIGHT_SIZE-1:0] Wgt_5_419,input [WEIGHT_SIZE-1:0] Wgt_5_420,input [WEIGHT_SIZE-1:0] Wgt_5_421,input [WEIGHT_SIZE-1:0] Wgt_5_422,input [WEIGHT_SIZE-1:0] Wgt_5_423,input [WEIGHT_SIZE-1:0] Wgt_5_424,input [WEIGHT_SIZE-1:0] Wgt_5_425,input [WEIGHT_SIZE-1:0] Wgt_5_426,input [WEIGHT_SIZE-1:0] Wgt_5_427,input [WEIGHT_SIZE-1:0] Wgt_5_428,input [WEIGHT_SIZE-1:0] Wgt_5_429,input [WEIGHT_SIZE-1:0] Wgt_5_430,input [WEIGHT_SIZE-1:0] Wgt_5_431,input [WEIGHT_SIZE-1:0] Wgt_5_432,input [WEIGHT_SIZE-1:0] Wgt_5_433,input [WEIGHT_SIZE-1:0] Wgt_5_434,input [WEIGHT_SIZE-1:0] Wgt_5_435,input [WEIGHT_SIZE-1:0] Wgt_5_436,input [WEIGHT_SIZE-1:0] Wgt_5_437,input [WEIGHT_SIZE-1:0] Wgt_5_438,input [WEIGHT_SIZE-1:0] Wgt_5_439,input [WEIGHT_SIZE-1:0] Wgt_5_440,input [WEIGHT_SIZE-1:0] Wgt_5_441,input [WEIGHT_SIZE-1:0] Wgt_5_442,input [WEIGHT_SIZE-1:0] Wgt_5_443,input [WEIGHT_SIZE-1:0] Wgt_5_444,input [WEIGHT_SIZE-1:0] Wgt_5_445,input [WEIGHT_SIZE-1:0] Wgt_5_446,input [WEIGHT_SIZE-1:0] Wgt_5_447,input [WEIGHT_SIZE-1:0] Wgt_5_448,input [WEIGHT_SIZE-1:0] Wgt_5_449,input [WEIGHT_SIZE-1:0] Wgt_5_450,input [WEIGHT_SIZE-1:0] Wgt_5_451,input [WEIGHT_SIZE-1:0] Wgt_5_452,input [WEIGHT_SIZE-1:0] Wgt_5_453,input [WEIGHT_SIZE-1:0] Wgt_5_454,input [WEIGHT_SIZE-1:0] Wgt_5_455,input [WEIGHT_SIZE-1:0] Wgt_5_456,input [WEIGHT_SIZE-1:0] Wgt_5_457,input [WEIGHT_SIZE-1:0] Wgt_5_458,input [WEIGHT_SIZE-1:0] Wgt_5_459,input [WEIGHT_SIZE-1:0] Wgt_5_460,input [WEIGHT_SIZE-1:0] Wgt_5_461,input [WEIGHT_SIZE-1:0] Wgt_5_462,input [WEIGHT_SIZE-1:0] Wgt_5_463,input [WEIGHT_SIZE-1:0] Wgt_5_464,input [WEIGHT_SIZE-1:0] Wgt_5_465,input [WEIGHT_SIZE-1:0] Wgt_5_466,input [WEIGHT_SIZE-1:0] Wgt_5_467,input [WEIGHT_SIZE-1:0] Wgt_5_468,input [WEIGHT_SIZE-1:0] Wgt_5_469,input [WEIGHT_SIZE-1:0] Wgt_5_470,input [WEIGHT_SIZE-1:0] Wgt_5_471,input [WEIGHT_SIZE-1:0] Wgt_5_472,input [WEIGHT_SIZE-1:0] Wgt_5_473,input [WEIGHT_SIZE-1:0] Wgt_5_474,input [WEIGHT_SIZE-1:0] Wgt_5_475,input [WEIGHT_SIZE-1:0] Wgt_5_476,input [WEIGHT_SIZE-1:0] Wgt_5_477,input [WEIGHT_SIZE-1:0] Wgt_5_478,input [WEIGHT_SIZE-1:0] Wgt_5_479,input [WEIGHT_SIZE-1:0] Wgt_5_480,input [WEIGHT_SIZE-1:0] Wgt_5_481,input [WEIGHT_SIZE-1:0] Wgt_5_482,input [WEIGHT_SIZE-1:0] Wgt_5_483,input [WEIGHT_SIZE-1:0] Wgt_5_484,input [WEIGHT_SIZE-1:0] Wgt_5_485,input [WEIGHT_SIZE-1:0] Wgt_5_486,input [WEIGHT_SIZE-1:0] Wgt_5_487,input [WEIGHT_SIZE-1:0] Wgt_5_488,input [WEIGHT_SIZE-1:0] Wgt_5_489,input [WEIGHT_SIZE-1:0] Wgt_5_490,input [WEIGHT_SIZE-1:0] Wgt_5_491,input [WEIGHT_SIZE-1:0] Wgt_5_492,input [WEIGHT_SIZE-1:0] Wgt_5_493,input [WEIGHT_SIZE-1:0] Wgt_5_494,input [WEIGHT_SIZE-1:0] Wgt_5_495,input [WEIGHT_SIZE-1:0] Wgt_5_496,input [WEIGHT_SIZE-1:0] Wgt_5_497,input [WEIGHT_SIZE-1:0] Wgt_5_498,input [WEIGHT_SIZE-1:0] Wgt_5_499,input [WEIGHT_SIZE-1:0] Wgt_5_500,input [WEIGHT_SIZE-1:0] Wgt_5_501,input [WEIGHT_SIZE-1:0] Wgt_5_502,input [WEIGHT_SIZE-1:0] Wgt_5_503,input [WEIGHT_SIZE-1:0] Wgt_5_504,input [WEIGHT_SIZE-1:0] Wgt_5_505,input [WEIGHT_SIZE-1:0] Wgt_5_506,input [WEIGHT_SIZE-1:0] Wgt_5_507,input [WEIGHT_SIZE-1:0] Wgt_5_508,input [WEIGHT_SIZE-1:0] Wgt_5_509,input [WEIGHT_SIZE-1:0] Wgt_5_510,input [WEIGHT_SIZE-1:0] Wgt_5_511,input [WEIGHT_SIZE-1:0] Wgt_5_512,input [WEIGHT_SIZE-1:0] Wgt_5_513,input [WEIGHT_SIZE-1:0] Wgt_5_514,input [WEIGHT_SIZE-1:0] Wgt_5_515,input [WEIGHT_SIZE-1:0] Wgt_5_516,input [WEIGHT_SIZE-1:0] Wgt_5_517,input [WEIGHT_SIZE-1:0] Wgt_5_518,input [WEIGHT_SIZE-1:0] Wgt_5_519,input [WEIGHT_SIZE-1:0] Wgt_5_520,input [WEIGHT_SIZE-1:0] Wgt_5_521,input [WEIGHT_SIZE-1:0] Wgt_5_522,input [WEIGHT_SIZE-1:0] Wgt_5_523,input [WEIGHT_SIZE-1:0] Wgt_5_524,input [WEIGHT_SIZE-1:0] Wgt_5_525,input [WEIGHT_SIZE-1:0] Wgt_5_526,input [WEIGHT_SIZE-1:0] Wgt_5_527,input [WEIGHT_SIZE-1:0] Wgt_5_528,input [WEIGHT_SIZE-1:0] Wgt_5_529,input [WEIGHT_SIZE-1:0] Wgt_5_530,input [WEIGHT_SIZE-1:0] Wgt_5_531,input [WEIGHT_SIZE-1:0] Wgt_5_532,input [WEIGHT_SIZE-1:0] Wgt_5_533,input [WEIGHT_SIZE-1:0] Wgt_5_534,input [WEIGHT_SIZE-1:0] Wgt_5_535,input [WEIGHT_SIZE-1:0] Wgt_5_536,input [WEIGHT_SIZE-1:0] Wgt_5_537,input [WEIGHT_SIZE-1:0] Wgt_5_538,input [WEIGHT_SIZE-1:0] Wgt_5_539,input [WEIGHT_SIZE-1:0] Wgt_5_540,input [WEIGHT_SIZE-1:0] Wgt_5_541,input [WEIGHT_SIZE-1:0] Wgt_5_542,input [WEIGHT_SIZE-1:0] Wgt_5_543,input [WEIGHT_SIZE-1:0] Wgt_5_544,input [WEIGHT_SIZE-1:0] Wgt_5_545,input [WEIGHT_SIZE-1:0] Wgt_5_546,input [WEIGHT_SIZE-1:0] Wgt_5_547,input [WEIGHT_SIZE-1:0] Wgt_5_548,input [WEIGHT_SIZE-1:0] Wgt_5_549,input [WEIGHT_SIZE-1:0] Wgt_5_550,input [WEIGHT_SIZE-1:0] Wgt_5_551,input [WEIGHT_SIZE-1:0] Wgt_5_552,input [WEIGHT_SIZE-1:0] Wgt_5_553,input [WEIGHT_SIZE-1:0] Wgt_5_554,input [WEIGHT_SIZE-1:0] Wgt_5_555,input [WEIGHT_SIZE-1:0] Wgt_5_556,input [WEIGHT_SIZE-1:0] Wgt_5_557,input [WEIGHT_SIZE-1:0] Wgt_5_558,input [WEIGHT_SIZE-1:0] Wgt_5_559,input [WEIGHT_SIZE-1:0] Wgt_5_560,input [WEIGHT_SIZE-1:0] Wgt_5_561,input [WEIGHT_SIZE-1:0] Wgt_5_562,input [WEIGHT_SIZE-1:0] Wgt_5_563,input [WEIGHT_SIZE-1:0] Wgt_5_564,input [WEIGHT_SIZE-1:0] Wgt_5_565,input [WEIGHT_SIZE-1:0] Wgt_5_566,input [WEIGHT_SIZE-1:0] Wgt_5_567,input [WEIGHT_SIZE-1:0] Wgt_5_568,input [WEIGHT_SIZE-1:0] Wgt_5_569,input [WEIGHT_SIZE-1:0] Wgt_5_570,input [WEIGHT_SIZE-1:0] Wgt_5_571,input [WEIGHT_SIZE-1:0] Wgt_5_572,input [WEIGHT_SIZE-1:0] Wgt_5_573,input [WEIGHT_SIZE-1:0] Wgt_5_574,input [WEIGHT_SIZE-1:0] Wgt_5_575,input [WEIGHT_SIZE-1:0] Wgt_5_576,input [WEIGHT_SIZE-1:0] Wgt_5_577,input [WEIGHT_SIZE-1:0] Wgt_5_578,input [WEIGHT_SIZE-1:0] Wgt_5_579,input [WEIGHT_SIZE-1:0] Wgt_5_580,input [WEIGHT_SIZE-1:0] Wgt_5_581,input [WEIGHT_SIZE-1:0] Wgt_5_582,input [WEIGHT_SIZE-1:0] Wgt_5_583,input [WEIGHT_SIZE-1:0] Wgt_5_584,input [WEIGHT_SIZE-1:0] Wgt_5_585,input [WEIGHT_SIZE-1:0] Wgt_5_586,input [WEIGHT_SIZE-1:0] Wgt_5_587,input [WEIGHT_SIZE-1:0] Wgt_5_588,input [WEIGHT_SIZE-1:0] Wgt_5_589,input [WEIGHT_SIZE-1:0] Wgt_5_590,input [WEIGHT_SIZE-1:0] Wgt_5_591,input [WEIGHT_SIZE-1:0] Wgt_5_592,input [WEIGHT_SIZE-1:0] Wgt_5_593,input [WEIGHT_SIZE-1:0] Wgt_5_594,input [WEIGHT_SIZE-1:0] Wgt_5_595,input [WEIGHT_SIZE-1:0] Wgt_5_596,input [WEIGHT_SIZE-1:0] Wgt_5_597,input [WEIGHT_SIZE-1:0] Wgt_5_598,input [WEIGHT_SIZE-1:0] Wgt_5_599,input [WEIGHT_SIZE-1:0] Wgt_5_600,input [WEIGHT_SIZE-1:0] Wgt_5_601,input [WEIGHT_SIZE-1:0] Wgt_5_602,input [WEIGHT_SIZE-1:0] Wgt_5_603,input [WEIGHT_SIZE-1:0] Wgt_5_604,input [WEIGHT_SIZE-1:0] Wgt_5_605,input [WEIGHT_SIZE-1:0] Wgt_5_606,input [WEIGHT_SIZE-1:0] Wgt_5_607,input [WEIGHT_SIZE-1:0] Wgt_5_608,input [WEIGHT_SIZE-1:0] Wgt_5_609,input [WEIGHT_SIZE-1:0] Wgt_5_610,input [WEIGHT_SIZE-1:0] Wgt_5_611,input [WEIGHT_SIZE-1:0] Wgt_5_612,input [WEIGHT_SIZE-1:0] Wgt_5_613,input [WEIGHT_SIZE-1:0] Wgt_5_614,input [WEIGHT_SIZE-1:0] Wgt_5_615,input [WEIGHT_SIZE-1:0] Wgt_5_616,input [WEIGHT_SIZE-1:0] Wgt_5_617,input [WEIGHT_SIZE-1:0] Wgt_5_618,input [WEIGHT_SIZE-1:0] Wgt_5_619,input [WEIGHT_SIZE-1:0] Wgt_5_620,input [WEIGHT_SIZE-1:0] Wgt_5_621,input [WEIGHT_SIZE-1:0] Wgt_5_622,input [WEIGHT_SIZE-1:0] Wgt_5_623,input [WEIGHT_SIZE-1:0] Wgt_5_624,input [WEIGHT_SIZE-1:0] Wgt_5_625,input [WEIGHT_SIZE-1:0] Wgt_5_626,input [WEIGHT_SIZE-1:0] Wgt_5_627,input [WEIGHT_SIZE-1:0] Wgt_5_628,input [WEIGHT_SIZE-1:0] Wgt_5_629,input [WEIGHT_SIZE-1:0] Wgt_5_630,input [WEIGHT_SIZE-1:0] Wgt_5_631,input [WEIGHT_SIZE-1:0] Wgt_5_632,input [WEIGHT_SIZE-1:0] Wgt_5_633,input [WEIGHT_SIZE-1:0] Wgt_5_634,input [WEIGHT_SIZE-1:0] Wgt_5_635,input [WEIGHT_SIZE-1:0] Wgt_5_636,input [WEIGHT_SIZE-1:0] Wgt_5_637,input [WEIGHT_SIZE-1:0] Wgt_5_638,input [WEIGHT_SIZE-1:0] Wgt_5_639,input [WEIGHT_SIZE-1:0] Wgt_5_640,input [WEIGHT_SIZE-1:0] Wgt_5_641,input [WEIGHT_SIZE-1:0] Wgt_5_642,input [WEIGHT_SIZE-1:0] Wgt_5_643,input [WEIGHT_SIZE-1:0] Wgt_5_644,input [WEIGHT_SIZE-1:0] Wgt_5_645,input [WEIGHT_SIZE-1:0] Wgt_5_646,input [WEIGHT_SIZE-1:0] Wgt_5_647,input [WEIGHT_SIZE-1:0] Wgt_5_648,input [WEIGHT_SIZE-1:0] Wgt_5_649,input [WEIGHT_SIZE-1:0] Wgt_5_650,input [WEIGHT_SIZE-1:0] Wgt_5_651,input [WEIGHT_SIZE-1:0] Wgt_5_652,input [WEIGHT_SIZE-1:0] Wgt_5_653,input [WEIGHT_SIZE-1:0] Wgt_5_654,input [WEIGHT_SIZE-1:0] Wgt_5_655,input [WEIGHT_SIZE-1:0] Wgt_5_656,input [WEIGHT_SIZE-1:0] Wgt_5_657,input [WEIGHT_SIZE-1:0] Wgt_5_658,input [WEIGHT_SIZE-1:0] Wgt_5_659,input [WEIGHT_SIZE-1:0] Wgt_5_660,input [WEIGHT_SIZE-1:0] Wgt_5_661,input [WEIGHT_SIZE-1:0] Wgt_5_662,input [WEIGHT_SIZE-1:0] Wgt_5_663,input [WEIGHT_SIZE-1:0] Wgt_5_664,input [WEIGHT_SIZE-1:0] Wgt_5_665,input [WEIGHT_SIZE-1:0] Wgt_5_666,input [WEIGHT_SIZE-1:0] Wgt_5_667,input [WEIGHT_SIZE-1:0] Wgt_5_668,input [WEIGHT_SIZE-1:0] Wgt_5_669,input [WEIGHT_SIZE-1:0] Wgt_5_670,input [WEIGHT_SIZE-1:0] Wgt_5_671,input [WEIGHT_SIZE-1:0] Wgt_5_672,input [WEIGHT_SIZE-1:0] Wgt_5_673,input [WEIGHT_SIZE-1:0] Wgt_5_674,input [WEIGHT_SIZE-1:0] Wgt_5_675,input [WEIGHT_SIZE-1:0] Wgt_5_676,input [WEIGHT_SIZE-1:0] Wgt_5_677,input [WEIGHT_SIZE-1:0] Wgt_5_678,input [WEIGHT_SIZE-1:0] Wgt_5_679,input [WEIGHT_SIZE-1:0] Wgt_5_680,input [WEIGHT_SIZE-1:0] Wgt_5_681,input [WEIGHT_SIZE-1:0] Wgt_5_682,input [WEIGHT_SIZE-1:0] Wgt_5_683,input [WEIGHT_SIZE-1:0] Wgt_5_684,input [WEIGHT_SIZE-1:0] Wgt_5_685,input [WEIGHT_SIZE-1:0] Wgt_5_686,input [WEIGHT_SIZE-1:0] Wgt_5_687,input [WEIGHT_SIZE-1:0] Wgt_5_688,input [WEIGHT_SIZE-1:0] Wgt_5_689,input [WEIGHT_SIZE-1:0] Wgt_5_690,input [WEIGHT_SIZE-1:0] Wgt_5_691,input [WEIGHT_SIZE-1:0] Wgt_5_692,input [WEIGHT_SIZE-1:0] Wgt_5_693,input [WEIGHT_SIZE-1:0] Wgt_5_694,input [WEIGHT_SIZE-1:0] Wgt_5_695,input [WEIGHT_SIZE-1:0] Wgt_5_696,input [WEIGHT_SIZE-1:0] Wgt_5_697,input [WEIGHT_SIZE-1:0] Wgt_5_698,input [WEIGHT_SIZE-1:0] Wgt_5_699,input [WEIGHT_SIZE-1:0] Wgt_5_700,input [WEIGHT_SIZE-1:0] Wgt_5_701,input [WEIGHT_SIZE-1:0] Wgt_5_702,input [WEIGHT_SIZE-1:0] Wgt_5_703,input [WEIGHT_SIZE-1:0] Wgt_5_704,input [WEIGHT_SIZE-1:0] Wgt_5_705,input [WEIGHT_SIZE-1:0] Wgt_5_706,input [WEIGHT_SIZE-1:0] Wgt_5_707,input [WEIGHT_SIZE-1:0] Wgt_5_708,input [WEIGHT_SIZE-1:0] Wgt_5_709,input [WEIGHT_SIZE-1:0] Wgt_5_710,input [WEIGHT_SIZE-1:0] Wgt_5_711,input [WEIGHT_SIZE-1:0] Wgt_5_712,input [WEIGHT_SIZE-1:0] Wgt_5_713,input [WEIGHT_SIZE-1:0] Wgt_5_714,input [WEIGHT_SIZE-1:0] Wgt_5_715,input [WEIGHT_SIZE-1:0] Wgt_5_716,input [WEIGHT_SIZE-1:0] Wgt_5_717,input [WEIGHT_SIZE-1:0] Wgt_5_718,input [WEIGHT_SIZE-1:0] Wgt_5_719,input [WEIGHT_SIZE-1:0] Wgt_5_720,input [WEIGHT_SIZE-1:0] Wgt_5_721,input [WEIGHT_SIZE-1:0] Wgt_5_722,input [WEIGHT_SIZE-1:0] Wgt_5_723,input [WEIGHT_SIZE-1:0] Wgt_5_724,input [WEIGHT_SIZE-1:0] Wgt_5_725,input [WEIGHT_SIZE-1:0] Wgt_5_726,input [WEIGHT_SIZE-1:0] Wgt_5_727,input [WEIGHT_SIZE-1:0] Wgt_5_728,input [WEIGHT_SIZE-1:0] Wgt_5_729,input [WEIGHT_SIZE-1:0] Wgt_5_730,input [WEIGHT_SIZE-1:0] Wgt_5_731,input [WEIGHT_SIZE-1:0] Wgt_5_732,input [WEIGHT_SIZE-1:0] Wgt_5_733,input [WEIGHT_SIZE-1:0] Wgt_5_734,input [WEIGHT_SIZE-1:0] Wgt_5_735,input [WEIGHT_SIZE-1:0] Wgt_5_736,input [WEIGHT_SIZE-1:0] Wgt_5_737,input [WEIGHT_SIZE-1:0] Wgt_5_738,input [WEIGHT_SIZE-1:0] Wgt_5_739,input [WEIGHT_SIZE-1:0] Wgt_5_740,input [WEIGHT_SIZE-1:0] Wgt_5_741,input [WEIGHT_SIZE-1:0] Wgt_5_742,input [WEIGHT_SIZE-1:0] Wgt_5_743,input [WEIGHT_SIZE-1:0] Wgt_5_744,input [WEIGHT_SIZE-1:0] Wgt_5_745,input [WEIGHT_SIZE-1:0] Wgt_5_746,input [WEIGHT_SIZE-1:0] Wgt_5_747,input [WEIGHT_SIZE-1:0] Wgt_5_748,input [WEIGHT_SIZE-1:0] Wgt_5_749,input [WEIGHT_SIZE-1:0] Wgt_5_750,input [WEIGHT_SIZE-1:0] Wgt_5_751,input [WEIGHT_SIZE-1:0] Wgt_5_752,input [WEIGHT_SIZE-1:0] Wgt_5_753,input [WEIGHT_SIZE-1:0] Wgt_5_754,input [WEIGHT_SIZE-1:0] Wgt_5_755,input [WEIGHT_SIZE-1:0] Wgt_5_756,input [WEIGHT_SIZE-1:0] Wgt_5_757,input [WEIGHT_SIZE-1:0] Wgt_5_758,input [WEIGHT_SIZE-1:0] Wgt_5_759,input [WEIGHT_SIZE-1:0] Wgt_5_760,input [WEIGHT_SIZE-1:0] Wgt_5_761,input [WEIGHT_SIZE-1:0] Wgt_5_762,input [WEIGHT_SIZE-1:0] Wgt_5_763,input [WEIGHT_SIZE-1:0] Wgt_5_764,input [WEIGHT_SIZE-1:0] Wgt_5_765,input [WEIGHT_SIZE-1:0] Wgt_5_766,input [WEIGHT_SIZE-1:0] Wgt_5_767,input [WEIGHT_SIZE-1:0] Wgt_5_768,input [WEIGHT_SIZE-1:0] Wgt_5_769,input [WEIGHT_SIZE-1:0] Wgt_5_770,input [WEIGHT_SIZE-1:0] Wgt_5_771,input [WEIGHT_SIZE-1:0] Wgt_5_772,input [WEIGHT_SIZE-1:0] Wgt_5_773,input [WEIGHT_SIZE-1:0] Wgt_5_774,input [WEIGHT_SIZE-1:0] Wgt_5_775,input [WEIGHT_SIZE-1:0] Wgt_5_776,input [WEIGHT_SIZE-1:0] Wgt_5_777,input [WEIGHT_SIZE-1:0] Wgt_5_778,input [WEIGHT_SIZE-1:0] Wgt_5_779,input [WEIGHT_SIZE-1:0] Wgt_5_780,input [WEIGHT_SIZE-1:0] Wgt_5_781,input [WEIGHT_SIZE-1:0] Wgt_5_782,input [WEIGHT_SIZE-1:0] Wgt_5_783,input [WEIGHT_SIZE-1:0] Wgt_5_784,input [WEIGHT_SIZE-1:0] Wgt_6_0,input [WEIGHT_SIZE-1:0] Wgt_6_1,input [WEIGHT_SIZE-1:0] Wgt_6_2,input [WEIGHT_SIZE-1:0] Wgt_6_3,input [WEIGHT_SIZE-1:0] Wgt_6_4,input [WEIGHT_SIZE-1:0] Wgt_6_5,input [WEIGHT_SIZE-1:0] Wgt_6_6,input [WEIGHT_SIZE-1:0] Wgt_6_7,input [WEIGHT_SIZE-1:0] Wgt_6_8,input [WEIGHT_SIZE-1:0] Wgt_6_9,input [WEIGHT_SIZE-1:0] Wgt_6_10,input [WEIGHT_SIZE-1:0] Wgt_6_11,input [WEIGHT_SIZE-1:0] Wgt_6_12,input [WEIGHT_SIZE-1:0] Wgt_6_13,input [WEIGHT_SIZE-1:0] Wgt_6_14,input [WEIGHT_SIZE-1:0] Wgt_6_15,input [WEIGHT_SIZE-1:0] Wgt_6_16,input [WEIGHT_SIZE-1:0] Wgt_6_17,input [WEIGHT_SIZE-1:0] Wgt_6_18,input [WEIGHT_SIZE-1:0] Wgt_6_19,input [WEIGHT_SIZE-1:0] Wgt_6_20,input [WEIGHT_SIZE-1:0] Wgt_6_21,input [WEIGHT_SIZE-1:0] Wgt_6_22,input [WEIGHT_SIZE-1:0] Wgt_6_23,input [WEIGHT_SIZE-1:0] Wgt_6_24,input [WEIGHT_SIZE-1:0] Wgt_6_25,input [WEIGHT_SIZE-1:0] Wgt_6_26,input [WEIGHT_SIZE-1:0] Wgt_6_27,input [WEIGHT_SIZE-1:0] Wgt_6_28,input [WEIGHT_SIZE-1:0] Wgt_6_29,input [WEIGHT_SIZE-1:0] Wgt_6_30,input [WEIGHT_SIZE-1:0] Wgt_6_31,input [WEIGHT_SIZE-1:0] Wgt_6_32,input [WEIGHT_SIZE-1:0] Wgt_6_33,input [WEIGHT_SIZE-1:0] Wgt_6_34,input [WEIGHT_SIZE-1:0] Wgt_6_35,input [WEIGHT_SIZE-1:0] Wgt_6_36,input [WEIGHT_SIZE-1:0] Wgt_6_37,input [WEIGHT_SIZE-1:0] Wgt_6_38,input [WEIGHT_SIZE-1:0] Wgt_6_39,input [WEIGHT_SIZE-1:0] Wgt_6_40,input [WEIGHT_SIZE-1:0] Wgt_6_41,input [WEIGHT_SIZE-1:0] Wgt_6_42,input [WEIGHT_SIZE-1:0] Wgt_6_43,input [WEIGHT_SIZE-1:0] Wgt_6_44,input [WEIGHT_SIZE-1:0] Wgt_6_45,input [WEIGHT_SIZE-1:0] Wgt_6_46,input [WEIGHT_SIZE-1:0] Wgt_6_47,input [WEIGHT_SIZE-1:0] Wgt_6_48,input [WEIGHT_SIZE-1:0] Wgt_6_49,input [WEIGHT_SIZE-1:0] Wgt_6_50,input [WEIGHT_SIZE-1:0] Wgt_6_51,input [WEIGHT_SIZE-1:0] Wgt_6_52,input [WEIGHT_SIZE-1:0] Wgt_6_53,input [WEIGHT_SIZE-1:0] Wgt_6_54,input [WEIGHT_SIZE-1:0] Wgt_6_55,input [WEIGHT_SIZE-1:0] Wgt_6_56,input [WEIGHT_SIZE-1:0] Wgt_6_57,input [WEIGHT_SIZE-1:0] Wgt_6_58,input [WEIGHT_SIZE-1:0] Wgt_6_59,input [WEIGHT_SIZE-1:0] Wgt_6_60,input [WEIGHT_SIZE-1:0] Wgt_6_61,input [WEIGHT_SIZE-1:0] Wgt_6_62,input [WEIGHT_SIZE-1:0] Wgt_6_63,input [WEIGHT_SIZE-1:0] Wgt_6_64,input [WEIGHT_SIZE-1:0] Wgt_6_65,input [WEIGHT_SIZE-1:0] Wgt_6_66,input [WEIGHT_SIZE-1:0] Wgt_6_67,input [WEIGHT_SIZE-1:0] Wgt_6_68,input [WEIGHT_SIZE-1:0] Wgt_6_69,input [WEIGHT_SIZE-1:0] Wgt_6_70,input [WEIGHT_SIZE-1:0] Wgt_6_71,input [WEIGHT_SIZE-1:0] Wgt_6_72,input [WEIGHT_SIZE-1:0] Wgt_6_73,input [WEIGHT_SIZE-1:0] Wgt_6_74,input [WEIGHT_SIZE-1:0] Wgt_6_75,input [WEIGHT_SIZE-1:0] Wgt_6_76,input [WEIGHT_SIZE-1:0] Wgt_6_77,input [WEIGHT_SIZE-1:0] Wgt_6_78,input [WEIGHT_SIZE-1:0] Wgt_6_79,input [WEIGHT_SIZE-1:0] Wgt_6_80,input [WEIGHT_SIZE-1:0] Wgt_6_81,input [WEIGHT_SIZE-1:0] Wgt_6_82,input [WEIGHT_SIZE-1:0] Wgt_6_83,input [WEIGHT_SIZE-1:0] Wgt_6_84,input [WEIGHT_SIZE-1:0] Wgt_6_85,input [WEIGHT_SIZE-1:0] Wgt_6_86,input [WEIGHT_SIZE-1:0] Wgt_6_87,input [WEIGHT_SIZE-1:0] Wgt_6_88,input [WEIGHT_SIZE-1:0] Wgt_6_89,input [WEIGHT_SIZE-1:0] Wgt_6_90,input [WEIGHT_SIZE-1:0] Wgt_6_91,input [WEIGHT_SIZE-1:0] Wgt_6_92,input [WEIGHT_SIZE-1:0] Wgt_6_93,input [WEIGHT_SIZE-1:0] Wgt_6_94,input [WEIGHT_SIZE-1:0] Wgt_6_95,input [WEIGHT_SIZE-1:0] Wgt_6_96,input [WEIGHT_SIZE-1:0] Wgt_6_97,input [WEIGHT_SIZE-1:0] Wgt_6_98,input [WEIGHT_SIZE-1:0] Wgt_6_99,input [WEIGHT_SIZE-1:0] Wgt_6_100,input [WEIGHT_SIZE-1:0] Wgt_6_101,input [WEIGHT_SIZE-1:0] Wgt_6_102,input [WEIGHT_SIZE-1:0] Wgt_6_103,input [WEIGHT_SIZE-1:0] Wgt_6_104,input [WEIGHT_SIZE-1:0] Wgt_6_105,input [WEIGHT_SIZE-1:0] Wgt_6_106,input [WEIGHT_SIZE-1:0] Wgt_6_107,input [WEIGHT_SIZE-1:0] Wgt_6_108,input [WEIGHT_SIZE-1:0] Wgt_6_109,input [WEIGHT_SIZE-1:0] Wgt_6_110,input [WEIGHT_SIZE-1:0] Wgt_6_111,input [WEIGHT_SIZE-1:0] Wgt_6_112,input [WEIGHT_SIZE-1:0] Wgt_6_113,input [WEIGHT_SIZE-1:0] Wgt_6_114,input [WEIGHT_SIZE-1:0] Wgt_6_115,input [WEIGHT_SIZE-1:0] Wgt_6_116,input [WEIGHT_SIZE-1:0] Wgt_6_117,input [WEIGHT_SIZE-1:0] Wgt_6_118,input [WEIGHT_SIZE-1:0] Wgt_6_119,input [WEIGHT_SIZE-1:0] Wgt_6_120,input [WEIGHT_SIZE-1:0] Wgt_6_121,input [WEIGHT_SIZE-1:0] Wgt_6_122,input [WEIGHT_SIZE-1:0] Wgt_6_123,input [WEIGHT_SIZE-1:0] Wgt_6_124,input [WEIGHT_SIZE-1:0] Wgt_6_125,input [WEIGHT_SIZE-1:0] Wgt_6_126,input [WEIGHT_SIZE-1:0] Wgt_6_127,input [WEIGHT_SIZE-1:0] Wgt_6_128,input [WEIGHT_SIZE-1:0] Wgt_6_129,input [WEIGHT_SIZE-1:0] Wgt_6_130,input [WEIGHT_SIZE-1:0] Wgt_6_131,input [WEIGHT_SIZE-1:0] Wgt_6_132,input [WEIGHT_SIZE-1:0] Wgt_6_133,input [WEIGHT_SIZE-1:0] Wgt_6_134,input [WEIGHT_SIZE-1:0] Wgt_6_135,input [WEIGHT_SIZE-1:0] Wgt_6_136,input [WEIGHT_SIZE-1:0] Wgt_6_137,input [WEIGHT_SIZE-1:0] Wgt_6_138,input [WEIGHT_SIZE-1:0] Wgt_6_139,input [WEIGHT_SIZE-1:0] Wgt_6_140,input [WEIGHT_SIZE-1:0] Wgt_6_141,input [WEIGHT_SIZE-1:0] Wgt_6_142,input [WEIGHT_SIZE-1:0] Wgt_6_143,input [WEIGHT_SIZE-1:0] Wgt_6_144,input [WEIGHT_SIZE-1:0] Wgt_6_145,input [WEIGHT_SIZE-1:0] Wgt_6_146,input [WEIGHT_SIZE-1:0] Wgt_6_147,input [WEIGHT_SIZE-1:0] Wgt_6_148,input [WEIGHT_SIZE-1:0] Wgt_6_149,input [WEIGHT_SIZE-1:0] Wgt_6_150,input [WEIGHT_SIZE-1:0] Wgt_6_151,input [WEIGHT_SIZE-1:0] Wgt_6_152,input [WEIGHT_SIZE-1:0] Wgt_6_153,input [WEIGHT_SIZE-1:0] Wgt_6_154,input [WEIGHT_SIZE-1:0] Wgt_6_155,input [WEIGHT_SIZE-1:0] Wgt_6_156,input [WEIGHT_SIZE-1:0] Wgt_6_157,input [WEIGHT_SIZE-1:0] Wgt_6_158,input [WEIGHT_SIZE-1:0] Wgt_6_159,input [WEIGHT_SIZE-1:0] Wgt_6_160,input [WEIGHT_SIZE-1:0] Wgt_6_161,input [WEIGHT_SIZE-1:0] Wgt_6_162,input [WEIGHT_SIZE-1:0] Wgt_6_163,input [WEIGHT_SIZE-1:0] Wgt_6_164,input [WEIGHT_SIZE-1:0] Wgt_6_165,input [WEIGHT_SIZE-1:0] Wgt_6_166,input [WEIGHT_SIZE-1:0] Wgt_6_167,input [WEIGHT_SIZE-1:0] Wgt_6_168,input [WEIGHT_SIZE-1:0] Wgt_6_169,input [WEIGHT_SIZE-1:0] Wgt_6_170,input [WEIGHT_SIZE-1:0] Wgt_6_171,input [WEIGHT_SIZE-1:0] Wgt_6_172,input [WEIGHT_SIZE-1:0] Wgt_6_173,input [WEIGHT_SIZE-1:0] Wgt_6_174,input [WEIGHT_SIZE-1:0] Wgt_6_175,input [WEIGHT_SIZE-1:0] Wgt_6_176,input [WEIGHT_SIZE-1:0] Wgt_6_177,input [WEIGHT_SIZE-1:0] Wgt_6_178,input [WEIGHT_SIZE-1:0] Wgt_6_179,input [WEIGHT_SIZE-1:0] Wgt_6_180,input [WEIGHT_SIZE-1:0] Wgt_6_181,input [WEIGHT_SIZE-1:0] Wgt_6_182,input [WEIGHT_SIZE-1:0] Wgt_6_183,input [WEIGHT_SIZE-1:0] Wgt_6_184,input [WEIGHT_SIZE-1:0] Wgt_6_185,input [WEIGHT_SIZE-1:0] Wgt_6_186,input [WEIGHT_SIZE-1:0] Wgt_6_187,input [WEIGHT_SIZE-1:0] Wgt_6_188,input [WEIGHT_SIZE-1:0] Wgt_6_189,input [WEIGHT_SIZE-1:0] Wgt_6_190,input [WEIGHT_SIZE-1:0] Wgt_6_191,input [WEIGHT_SIZE-1:0] Wgt_6_192,input [WEIGHT_SIZE-1:0] Wgt_6_193,input [WEIGHT_SIZE-1:0] Wgt_6_194,input [WEIGHT_SIZE-1:0] Wgt_6_195,input [WEIGHT_SIZE-1:0] Wgt_6_196,input [WEIGHT_SIZE-1:0] Wgt_6_197,input [WEIGHT_SIZE-1:0] Wgt_6_198,input [WEIGHT_SIZE-1:0] Wgt_6_199,input [WEIGHT_SIZE-1:0] Wgt_6_200,input [WEIGHT_SIZE-1:0] Wgt_6_201,input [WEIGHT_SIZE-1:0] Wgt_6_202,input [WEIGHT_SIZE-1:0] Wgt_6_203,input [WEIGHT_SIZE-1:0] Wgt_6_204,input [WEIGHT_SIZE-1:0] Wgt_6_205,input [WEIGHT_SIZE-1:0] Wgt_6_206,input [WEIGHT_SIZE-1:0] Wgt_6_207,input [WEIGHT_SIZE-1:0] Wgt_6_208,input [WEIGHT_SIZE-1:0] Wgt_6_209,input [WEIGHT_SIZE-1:0] Wgt_6_210,input [WEIGHT_SIZE-1:0] Wgt_6_211,input [WEIGHT_SIZE-1:0] Wgt_6_212,input [WEIGHT_SIZE-1:0] Wgt_6_213,input [WEIGHT_SIZE-1:0] Wgt_6_214,input [WEIGHT_SIZE-1:0] Wgt_6_215,input [WEIGHT_SIZE-1:0] Wgt_6_216,input [WEIGHT_SIZE-1:0] Wgt_6_217,input [WEIGHT_SIZE-1:0] Wgt_6_218,input [WEIGHT_SIZE-1:0] Wgt_6_219,input [WEIGHT_SIZE-1:0] Wgt_6_220,input [WEIGHT_SIZE-1:0] Wgt_6_221,input [WEIGHT_SIZE-1:0] Wgt_6_222,input [WEIGHT_SIZE-1:0] Wgt_6_223,input [WEIGHT_SIZE-1:0] Wgt_6_224,input [WEIGHT_SIZE-1:0] Wgt_6_225,input [WEIGHT_SIZE-1:0] Wgt_6_226,input [WEIGHT_SIZE-1:0] Wgt_6_227,input [WEIGHT_SIZE-1:0] Wgt_6_228,input [WEIGHT_SIZE-1:0] Wgt_6_229,input [WEIGHT_SIZE-1:0] Wgt_6_230,input [WEIGHT_SIZE-1:0] Wgt_6_231,input [WEIGHT_SIZE-1:0] Wgt_6_232,input [WEIGHT_SIZE-1:0] Wgt_6_233,input [WEIGHT_SIZE-1:0] Wgt_6_234,input [WEIGHT_SIZE-1:0] Wgt_6_235,input [WEIGHT_SIZE-1:0] Wgt_6_236,input [WEIGHT_SIZE-1:0] Wgt_6_237,input [WEIGHT_SIZE-1:0] Wgt_6_238,input [WEIGHT_SIZE-1:0] Wgt_6_239,input [WEIGHT_SIZE-1:0] Wgt_6_240,input [WEIGHT_SIZE-1:0] Wgt_6_241,input [WEIGHT_SIZE-1:0] Wgt_6_242,input [WEIGHT_SIZE-1:0] Wgt_6_243,input [WEIGHT_SIZE-1:0] Wgt_6_244,input [WEIGHT_SIZE-1:0] Wgt_6_245,input [WEIGHT_SIZE-1:0] Wgt_6_246,input [WEIGHT_SIZE-1:0] Wgt_6_247,input [WEIGHT_SIZE-1:0] Wgt_6_248,input [WEIGHT_SIZE-1:0] Wgt_6_249,input [WEIGHT_SIZE-1:0] Wgt_6_250,input [WEIGHT_SIZE-1:0] Wgt_6_251,input [WEIGHT_SIZE-1:0] Wgt_6_252,input [WEIGHT_SIZE-1:0] Wgt_6_253,input [WEIGHT_SIZE-1:0] Wgt_6_254,input [WEIGHT_SIZE-1:0] Wgt_6_255,input [WEIGHT_SIZE-1:0] Wgt_6_256,input [WEIGHT_SIZE-1:0] Wgt_6_257,input [WEIGHT_SIZE-1:0] Wgt_6_258,input [WEIGHT_SIZE-1:0] Wgt_6_259,input [WEIGHT_SIZE-1:0] Wgt_6_260,input [WEIGHT_SIZE-1:0] Wgt_6_261,input [WEIGHT_SIZE-1:0] Wgt_6_262,input [WEIGHT_SIZE-1:0] Wgt_6_263,input [WEIGHT_SIZE-1:0] Wgt_6_264,input [WEIGHT_SIZE-1:0] Wgt_6_265,input [WEIGHT_SIZE-1:0] Wgt_6_266,input [WEIGHT_SIZE-1:0] Wgt_6_267,input [WEIGHT_SIZE-1:0] Wgt_6_268,input [WEIGHT_SIZE-1:0] Wgt_6_269,input [WEIGHT_SIZE-1:0] Wgt_6_270,input [WEIGHT_SIZE-1:0] Wgt_6_271,input [WEIGHT_SIZE-1:0] Wgt_6_272,input [WEIGHT_SIZE-1:0] Wgt_6_273,input [WEIGHT_SIZE-1:0] Wgt_6_274,input [WEIGHT_SIZE-1:0] Wgt_6_275,input [WEIGHT_SIZE-1:0] Wgt_6_276,input [WEIGHT_SIZE-1:0] Wgt_6_277,input [WEIGHT_SIZE-1:0] Wgt_6_278,input [WEIGHT_SIZE-1:0] Wgt_6_279,input [WEIGHT_SIZE-1:0] Wgt_6_280,input [WEIGHT_SIZE-1:0] Wgt_6_281,input [WEIGHT_SIZE-1:0] Wgt_6_282,input [WEIGHT_SIZE-1:0] Wgt_6_283,input [WEIGHT_SIZE-1:0] Wgt_6_284,input [WEIGHT_SIZE-1:0] Wgt_6_285,input [WEIGHT_SIZE-1:0] Wgt_6_286,input [WEIGHT_SIZE-1:0] Wgt_6_287,input [WEIGHT_SIZE-1:0] Wgt_6_288,input [WEIGHT_SIZE-1:0] Wgt_6_289,input [WEIGHT_SIZE-1:0] Wgt_6_290,input [WEIGHT_SIZE-1:0] Wgt_6_291,input [WEIGHT_SIZE-1:0] Wgt_6_292,input [WEIGHT_SIZE-1:0] Wgt_6_293,input [WEIGHT_SIZE-1:0] Wgt_6_294,input [WEIGHT_SIZE-1:0] Wgt_6_295,input [WEIGHT_SIZE-1:0] Wgt_6_296,input [WEIGHT_SIZE-1:0] Wgt_6_297,input [WEIGHT_SIZE-1:0] Wgt_6_298,input [WEIGHT_SIZE-1:0] Wgt_6_299,input [WEIGHT_SIZE-1:0] Wgt_6_300,input [WEIGHT_SIZE-1:0] Wgt_6_301,input [WEIGHT_SIZE-1:0] Wgt_6_302,input [WEIGHT_SIZE-1:0] Wgt_6_303,input [WEIGHT_SIZE-1:0] Wgt_6_304,input [WEIGHT_SIZE-1:0] Wgt_6_305,input [WEIGHT_SIZE-1:0] Wgt_6_306,input [WEIGHT_SIZE-1:0] Wgt_6_307,input [WEIGHT_SIZE-1:0] Wgt_6_308,input [WEIGHT_SIZE-1:0] Wgt_6_309,input [WEIGHT_SIZE-1:0] Wgt_6_310,input [WEIGHT_SIZE-1:0] Wgt_6_311,input [WEIGHT_SIZE-1:0] Wgt_6_312,input [WEIGHT_SIZE-1:0] Wgt_6_313,input [WEIGHT_SIZE-1:0] Wgt_6_314,input [WEIGHT_SIZE-1:0] Wgt_6_315,input [WEIGHT_SIZE-1:0] Wgt_6_316,input [WEIGHT_SIZE-1:0] Wgt_6_317,input [WEIGHT_SIZE-1:0] Wgt_6_318,input [WEIGHT_SIZE-1:0] Wgt_6_319,input [WEIGHT_SIZE-1:0] Wgt_6_320,input [WEIGHT_SIZE-1:0] Wgt_6_321,input [WEIGHT_SIZE-1:0] Wgt_6_322,input [WEIGHT_SIZE-1:0] Wgt_6_323,input [WEIGHT_SIZE-1:0] Wgt_6_324,input [WEIGHT_SIZE-1:0] Wgt_6_325,input [WEIGHT_SIZE-1:0] Wgt_6_326,input [WEIGHT_SIZE-1:0] Wgt_6_327,input [WEIGHT_SIZE-1:0] Wgt_6_328,input [WEIGHT_SIZE-1:0] Wgt_6_329,input [WEIGHT_SIZE-1:0] Wgt_6_330,input [WEIGHT_SIZE-1:0] Wgt_6_331,input [WEIGHT_SIZE-1:0] Wgt_6_332,input [WEIGHT_SIZE-1:0] Wgt_6_333,input [WEIGHT_SIZE-1:0] Wgt_6_334,input [WEIGHT_SIZE-1:0] Wgt_6_335,input [WEIGHT_SIZE-1:0] Wgt_6_336,input [WEIGHT_SIZE-1:0] Wgt_6_337,input [WEIGHT_SIZE-1:0] Wgt_6_338,input [WEIGHT_SIZE-1:0] Wgt_6_339,input [WEIGHT_SIZE-1:0] Wgt_6_340,input [WEIGHT_SIZE-1:0] Wgt_6_341,input [WEIGHT_SIZE-1:0] Wgt_6_342,input [WEIGHT_SIZE-1:0] Wgt_6_343,input [WEIGHT_SIZE-1:0] Wgt_6_344,input [WEIGHT_SIZE-1:0] Wgt_6_345,input [WEIGHT_SIZE-1:0] Wgt_6_346,input [WEIGHT_SIZE-1:0] Wgt_6_347,input [WEIGHT_SIZE-1:0] Wgt_6_348,input [WEIGHT_SIZE-1:0] Wgt_6_349,input [WEIGHT_SIZE-1:0] Wgt_6_350,input [WEIGHT_SIZE-1:0] Wgt_6_351,input [WEIGHT_SIZE-1:0] Wgt_6_352,input [WEIGHT_SIZE-1:0] Wgt_6_353,input [WEIGHT_SIZE-1:0] Wgt_6_354,input [WEIGHT_SIZE-1:0] Wgt_6_355,input [WEIGHT_SIZE-1:0] Wgt_6_356,input [WEIGHT_SIZE-1:0] Wgt_6_357,input [WEIGHT_SIZE-1:0] Wgt_6_358,input [WEIGHT_SIZE-1:0] Wgt_6_359,input [WEIGHT_SIZE-1:0] Wgt_6_360,input [WEIGHT_SIZE-1:0] Wgt_6_361,input [WEIGHT_SIZE-1:0] Wgt_6_362,input [WEIGHT_SIZE-1:0] Wgt_6_363,input [WEIGHT_SIZE-1:0] Wgt_6_364,input [WEIGHT_SIZE-1:0] Wgt_6_365,input [WEIGHT_SIZE-1:0] Wgt_6_366,input [WEIGHT_SIZE-1:0] Wgt_6_367,input [WEIGHT_SIZE-1:0] Wgt_6_368,input [WEIGHT_SIZE-1:0] Wgt_6_369,input [WEIGHT_SIZE-1:0] Wgt_6_370,input [WEIGHT_SIZE-1:0] Wgt_6_371,input [WEIGHT_SIZE-1:0] Wgt_6_372,input [WEIGHT_SIZE-1:0] Wgt_6_373,input [WEIGHT_SIZE-1:0] Wgt_6_374,input [WEIGHT_SIZE-1:0] Wgt_6_375,input [WEIGHT_SIZE-1:0] Wgt_6_376,input [WEIGHT_SIZE-1:0] Wgt_6_377,input [WEIGHT_SIZE-1:0] Wgt_6_378,input [WEIGHT_SIZE-1:0] Wgt_6_379,input [WEIGHT_SIZE-1:0] Wgt_6_380,input [WEIGHT_SIZE-1:0] Wgt_6_381,input [WEIGHT_SIZE-1:0] Wgt_6_382,input [WEIGHT_SIZE-1:0] Wgt_6_383,input [WEIGHT_SIZE-1:0] Wgt_6_384,input [WEIGHT_SIZE-1:0] Wgt_6_385,input [WEIGHT_SIZE-1:0] Wgt_6_386,input [WEIGHT_SIZE-1:0] Wgt_6_387,input [WEIGHT_SIZE-1:0] Wgt_6_388,input [WEIGHT_SIZE-1:0] Wgt_6_389,input [WEIGHT_SIZE-1:0] Wgt_6_390,input [WEIGHT_SIZE-1:0] Wgt_6_391,input [WEIGHT_SIZE-1:0] Wgt_6_392,input [WEIGHT_SIZE-1:0] Wgt_6_393,input [WEIGHT_SIZE-1:0] Wgt_6_394,input [WEIGHT_SIZE-1:0] Wgt_6_395,input [WEIGHT_SIZE-1:0] Wgt_6_396,input [WEIGHT_SIZE-1:0] Wgt_6_397,input [WEIGHT_SIZE-1:0] Wgt_6_398,input [WEIGHT_SIZE-1:0] Wgt_6_399,input [WEIGHT_SIZE-1:0] Wgt_6_400,input [WEIGHT_SIZE-1:0] Wgt_6_401,input [WEIGHT_SIZE-1:0] Wgt_6_402,input [WEIGHT_SIZE-1:0] Wgt_6_403,input [WEIGHT_SIZE-1:0] Wgt_6_404,input [WEIGHT_SIZE-1:0] Wgt_6_405,input [WEIGHT_SIZE-1:0] Wgt_6_406,input [WEIGHT_SIZE-1:0] Wgt_6_407,input [WEIGHT_SIZE-1:0] Wgt_6_408,input [WEIGHT_SIZE-1:0] Wgt_6_409,input [WEIGHT_SIZE-1:0] Wgt_6_410,input [WEIGHT_SIZE-1:0] Wgt_6_411,input [WEIGHT_SIZE-1:0] Wgt_6_412,input [WEIGHT_SIZE-1:0] Wgt_6_413,input [WEIGHT_SIZE-1:0] Wgt_6_414,input [WEIGHT_SIZE-1:0] Wgt_6_415,input [WEIGHT_SIZE-1:0] Wgt_6_416,input [WEIGHT_SIZE-1:0] Wgt_6_417,input [WEIGHT_SIZE-1:0] Wgt_6_418,input [WEIGHT_SIZE-1:0] Wgt_6_419,input [WEIGHT_SIZE-1:0] Wgt_6_420,input [WEIGHT_SIZE-1:0] Wgt_6_421,input [WEIGHT_SIZE-1:0] Wgt_6_422,input [WEIGHT_SIZE-1:0] Wgt_6_423,input [WEIGHT_SIZE-1:0] Wgt_6_424,input [WEIGHT_SIZE-1:0] Wgt_6_425,input [WEIGHT_SIZE-1:0] Wgt_6_426,input [WEIGHT_SIZE-1:0] Wgt_6_427,input [WEIGHT_SIZE-1:0] Wgt_6_428,input [WEIGHT_SIZE-1:0] Wgt_6_429,input [WEIGHT_SIZE-1:0] Wgt_6_430,input [WEIGHT_SIZE-1:0] Wgt_6_431,input [WEIGHT_SIZE-1:0] Wgt_6_432,input [WEIGHT_SIZE-1:0] Wgt_6_433,input [WEIGHT_SIZE-1:0] Wgt_6_434,input [WEIGHT_SIZE-1:0] Wgt_6_435,input [WEIGHT_SIZE-1:0] Wgt_6_436,input [WEIGHT_SIZE-1:0] Wgt_6_437,input [WEIGHT_SIZE-1:0] Wgt_6_438,input [WEIGHT_SIZE-1:0] Wgt_6_439,input [WEIGHT_SIZE-1:0] Wgt_6_440,input [WEIGHT_SIZE-1:0] Wgt_6_441,input [WEIGHT_SIZE-1:0] Wgt_6_442,input [WEIGHT_SIZE-1:0] Wgt_6_443,input [WEIGHT_SIZE-1:0] Wgt_6_444,input [WEIGHT_SIZE-1:0] Wgt_6_445,input [WEIGHT_SIZE-1:0] Wgt_6_446,input [WEIGHT_SIZE-1:0] Wgt_6_447,input [WEIGHT_SIZE-1:0] Wgt_6_448,input [WEIGHT_SIZE-1:0] Wgt_6_449,input [WEIGHT_SIZE-1:0] Wgt_6_450,input [WEIGHT_SIZE-1:0] Wgt_6_451,input [WEIGHT_SIZE-1:0] Wgt_6_452,input [WEIGHT_SIZE-1:0] Wgt_6_453,input [WEIGHT_SIZE-1:0] Wgt_6_454,input [WEIGHT_SIZE-1:0] Wgt_6_455,input [WEIGHT_SIZE-1:0] Wgt_6_456,input [WEIGHT_SIZE-1:0] Wgt_6_457,input [WEIGHT_SIZE-1:0] Wgt_6_458,input [WEIGHT_SIZE-1:0] Wgt_6_459,input [WEIGHT_SIZE-1:0] Wgt_6_460,input [WEIGHT_SIZE-1:0] Wgt_6_461,input [WEIGHT_SIZE-1:0] Wgt_6_462,input [WEIGHT_SIZE-1:0] Wgt_6_463,input [WEIGHT_SIZE-1:0] Wgt_6_464,input [WEIGHT_SIZE-1:0] Wgt_6_465,input [WEIGHT_SIZE-1:0] Wgt_6_466,input [WEIGHT_SIZE-1:0] Wgt_6_467,input [WEIGHT_SIZE-1:0] Wgt_6_468,input [WEIGHT_SIZE-1:0] Wgt_6_469,input [WEIGHT_SIZE-1:0] Wgt_6_470,input [WEIGHT_SIZE-1:0] Wgt_6_471,input [WEIGHT_SIZE-1:0] Wgt_6_472,input [WEIGHT_SIZE-1:0] Wgt_6_473,input [WEIGHT_SIZE-1:0] Wgt_6_474,input [WEIGHT_SIZE-1:0] Wgt_6_475,input [WEIGHT_SIZE-1:0] Wgt_6_476,input [WEIGHT_SIZE-1:0] Wgt_6_477,input [WEIGHT_SIZE-1:0] Wgt_6_478,input [WEIGHT_SIZE-1:0] Wgt_6_479,input [WEIGHT_SIZE-1:0] Wgt_6_480,input [WEIGHT_SIZE-1:0] Wgt_6_481,input [WEIGHT_SIZE-1:0] Wgt_6_482,input [WEIGHT_SIZE-1:0] Wgt_6_483,input [WEIGHT_SIZE-1:0] Wgt_6_484,input [WEIGHT_SIZE-1:0] Wgt_6_485,input [WEIGHT_SIZE-1:0] Wgt_6_486,input [WEIGHT_SIZE-1:0] Wgt_6_487,input [WEIGHT_SIZE-1:0] Wgt_6_488,input [WEIGHT_SIZE-1:0] Wgt_6_489,input [WEIGHT_SIZE-1:0] Wgt_6_490,input [WEIGHT_SIZE-1:0] Wgt_6_491,input [WEIGHT_SIZE-1:0] Wgt_6_492,input [WEIGHT_SIZE-1:0] Wgt_6_493,input [WEIGHT_SIZE-1:0] Wgt_6_494,input [WEIGHT_SIZE-1:0] Wgt_6_495,input [WEIGHT_SIZE-1:0] Wgt_6_496,input [WEIGHT_SIZE-1:0] Wgt_6_497,input [WEIGHT_SIZE-1:0] Wgt_6_498,input [WEIGHT_SIZE-1:0] Wgt_6_499,input [WEIGHT_SIZE-1:0] Wgt_6_500,input [WEIGHT_SIZE-1:0] Wgt_6_501,input [WEIGHT_SIZE-1:0] Wgt_6_502,input [WEIGHT_SIZE-1:0] Wgt_6_503,input [WEIGHT_SIZE-1:0] Wgt_6_504,input [WEIGHT_SIZE-1:0] Wgt_6_505,input [WEIGHT_SIZE-1:0] Wgt_6_506,input [WEIGHT_SIZE-1:0] Wgt_6_507,input [WEIGHT_SIZE-1:0] Wgt_6_508,input [WEIGHT_SIZE-1:0] Wgt_6_509,input [WEIGHT_SIZE-1:0] Wgt_6_510,input [WEIGHT_SIZE-1:0] Wgt_6_511,input [WEIGHT_SIZE-1:0] Wgt_6_512,input [WEIGHT_SIZE-1:0] Wgt_6_513,input [WEIGHT_SIZE-1:0] Wgt_6_514,input [WEIGHT_SIZE-1:0] Wgt_6_515,input [WEIGHT_SIZE-1:0] Wgt_6_516,input [WEIGHT_SIZE-1:0] Wgt_6_517,input [WEIGHT_SIZE-1:0] Wgt_6_518,input [WEIGHT_SIZE-1:0] Wgt_6_519,input [WEIGHT_SIZE-1:0] Wgt_6_520,input [WEIGHT_SIZE-1:0] Wgt_6_521,input [WEIGHT_SIZE-1:0] Wgt_6_522,input [WEIGHT_SIZE-1:0] Wgt_6_523,input [WEIGHT_SIZE-1:0] Wgt_6_524,input [WEIGHT_SIZE-1:0] Wgt_6_525,input [WEIGHT_SIZE-1:0] Wgt_6_526,input [WEIGHT_SIZE-1:0] Wgt_6_527,input [WEIGHT_SIZE-1:0] Wgt_6_528,input [WEIGHT_SIZE-1:0] Wgt_6_529,input [WEIGHT_SIZE-1:0] Wgt_6_530,input [WEIGHT_SIZE-1:0] Wgt_6_531,input [WEIGHT_SIZE-1:0] Wgt_6_532,input [WEIGHT_SIZE-1:0] Wgt_6_533,input [WEIGHT_SIZE-1:0] Wgt_6_534,input [WEIGHT_SIZE-1:0] Wgt_6_535,input [WEIGHT_SIZE-1:0] Wgt_6_536,input [WEIGHT_SIZE-1:0] Wgt_6_537,input [WEIGHT_SIZE-1:0] Wgt_6_538,input [WEIGHT_SIZE-1:0] Wgt_6_539,input [WEIGHT_SIZE-1:0] Wgt_6_540,input [WEIGHT_SIZE-1:0] Wgt_6_541,input [WEIGHT_SIZE-1:0] Wgt_6_542,input [WEIGHT_SIZE-1:0] Wgt_6_543,input [WEIGHT_SIZE-1:0] Wgt_6_544,input [WEIGHT_SIZE-1:0] Wgt_6_545,input [WEIGHT_SIZE-1:0] Wgt_6_546,input [WEIGHT_SIZE-1:0] Wgt_6_547,input [WEIGHT_SIZE-1:0] Wgt_6_548,input [WEIGHT_SIZE-1:0] Wgt_6_549,input [WEIGHT_SIZE-1:0] Wgt_6_550,input [WEIGHT_SIZE-1:0] Wgt_6_551,input [WEIGHT_SIZE-1:0] Wgt_6_552,input [WEIGHT_SIZE-1:0] Wgt_6_553,input [WEIGHT_SIZE-1:0] Wgt_6_554,input [WEIGHT_SIZE-1:0] Wgt_6_555,input [WEIGHT_SIZE-1:0] Wgt_6_556,input [WEIGHT_SIZE-1:0] Wgt_6_557,input [WEIGHT_SIZE-1:0] Wgt_6_558,input [WEIGHT_SIZE-1:0] Wgt_6_559,input [WEIGHT_SIZE-1:0] Wgt_6_560,input [WEIGHT_SIZE-1:0] Wgt_6_561,input [WEIGHT_SIZE-1:0] Wgt_6_562,input [WEIGHT_SIZE-1:0] Wgt_6_563,input [WEIGHT_SIZE-1:0] Wgt_6_564,input [WEIGHT_SIZE-1:0] Wgt_6_565,input [WEIGHT_SIZE-1:0] Wgt_6_566,input [WEIGHT_SIZE-1:0] Wgt_6_567,input [WEIGHT_SIZE-1:0] Wgt_6_568,input [WEIGHT_SIZE-1:0] Wgt_6_569,input [WEIGHT_SIZE-1:0] Wgt_6_570,input [WEIGHT_SIZE-1:0] Wgt_6_571,input [WEIGHT_SIZE-1:0] Wgt_6_572,input [WEIGHT_SIZE-1:0] Wgt_6_573,input [WEIGHT_SIZE-1:0] Wgt_6_574,input [WEIGHT_SIZE-1:0] Wgt_6_575,input [WEIGHT_SIZE-1:0] Wgt_6_576,input [WEIGHT_SIZE-1:0] Wgt_6_577,input [WEIGHT_SIZE-1:0] Wgt_6_578,input [WEIGHT_SIZE-1:0] Wgt_6_579,input [WEIGHT_SIZE-1:0] Wgt_6_580,input [WEIGHT_SIZE-1:0] Wgt_6_581,input [WEIGHT_SIZE-1:0] Wgt_6_582,input [WEIGHT_SIZE-1:0] Wgt_6_583,input [WEIGHT_SIZE-1:0] Wgt_6_584,input [WEIGHT_SIZE-1:0] Wgt_6_585,input [WEIGHT_SIZE-1:0] Wgt_6_586,input [WEIGHT_SIZE-1:0] Wgt_6_587,input [WEIGHT_SIZE-1:0] Wgt_6_588,input [WEIGHT_SIZE-1:0] Wgt_6_589,input [WEIGHT_SIZE-1:0] Wgt_6_590,input [WEIGHT_SIZE-1:0] Wgt_6_591,input [WEIGHT_SIZE-1:0] Wgt_6_592,input [WEIGHT_SIZE-1:0] Wgt_6_593,input [WEIGHT_SIZE-1:0] Wgt_6_594,input [WEIGHT_SIZE-1:0] Wgt_6_595,input [WEIGHT_SIZE-1:0] Wgt_6_596,input [WEIGHT_SIZE-1:0] Wgt_6_597,input [WEIGHT_SIZE-1:0] Wgt_6_598,input [WEIGHT_SIZE-1:0] Wgt_6_599,input [WEIGHT_SIZE-1:0] Wgt_6_600,input [WEIGHT_SIZE-1:0] Wgt_6_601,input [WEIGHT_SIZE-1:0] Wgt_6_602,input [WEIGHT_SIZE-1:0] Wgt_6_603,input [WEIGHT_SIZE-1:0] Wgt_6_604,input [WEIGHT_SIZE-1:0] Wgt_6_605,input [WEIGHT_SIZE-1:0] Wgt_6_606,input [WEIGHT_SIZE-1:0] Wgt_6_607,input [WEIGHT_SIZE-1:0] Wgt_6_608,input [WEIGHT_SIZE-1:0] Wgt_6_609,input [WEIGHT_SIZE-1:0] Wgt_6_610,input [WEIGHT_SIZE-1:0] Wgt_6_611,input [WEIGHT_SIZE-1:0] Wgt_6_612,input [WEIGHT_SIZE-1:0] Wgt_6_613,input [WEIGHT_SIZE-1:0] Wgt_6_614,input [WEIGHT_SIZE-1:0] Wgt_6_615,input [WEIGHT_SIZE-1:0] Wgt_6_616,input [WEIGHT_SIZE-1:0] Wgt_6_617,input [WEIGHT_SIZE-1:0] Wgt_6_618,input [WEIGHT_SIZE-1:0] Wgt_6_619,input [WEIGHT_SIZE-1:0] Wgt_6_620,input [WEIGHT_SIZE-1:0] Wgt_6_621,input [WEIGHT_SIZE-1:0] Wgt_6_622,input [WEIGHT_SIZE-1:0] Wgt_6_623,input [WEIGHT_SIZE-1:0] Wgt_6_624,input [WEIGHT_SIZE-1:0] Wgt_6_625,input [WEIGHT_SIZE-1:0] Wgt_6_626,input [WEIGHT_SIZE-1:0] Wgt_6_627,input [WEIGHT_SIZE-1:0] Wgt_6_628,input [WEIGHT_SIZE-1:0] Wgt_6_629,input [WEIGHT_SIZE-1:0] Wgt_6_630,input [WEIGHT_SIZE-1:0] Wgt_6_631,input [WEIGHT_SIZE-1:0] Wgt_6_632,input [WEIGHT_SIZE-1:0] Wgt_6_633,input [WEIGHT_SIZE-1:0] Wgt_6_634,input [WEIGHT_SIZE-1:0] Wgt_6_635,input [WEIGHT_SIZE-1:0] Wgt_6_636,input [WEIGHT_SIZE-1:0] Wgt_6_637,input [WEIGHT_SIZE-1:0] Wgt_6_638,input [WEIGHT_SIZE-1:0] Wgt_6_639,input [WEIGHT_SIZE-1:0] Wgt_6_640,input [WEIGHT_SIZE-1:0] Wgt_6_641,input [WEIGHT_SIZE-1:0] Wgt_6_642,input [WEIGHT_SIZE-1:0] Wgt_6_643,input [WEIGHT_SIZE-1:0] Wgt_6_644,input [WEIGHT_SIZE-1:0] Wgt_6_645,input [WEIGHT_SIZE-1:0] Wgt_6_646,input [WEIGHT_SIZE-1:0] Wgt_6_647,input [WEIGHT_SIZE-1:0] Wgt_6_648,input [WEIGHT_SIZE-1:0] Wgt_6_649,input [WEIGHT_SIZE-1:0] Wgt_6_650,input [WEIGHT_SIZE-1:0] Wgt_6_651,input [WEIGHT_SIZE-1:0] Wgt_6_652,input [WEIGHT_SIZE-1:0] Wgt_6_653,input [WEIGHT_SIZE-1:0] Wgt_6_654,input [WEIGHT_SIZE-1:0] Wgt_6_655,input [WEIGHT_SIZE-1:0] Wgt_6_656,input [WEIGHT_SIZE-1:0] Wgt_6_657,input [WEIGHT_SIZE-1:0] Wgt_6_658,input [WEIGHT_SIZE-1:0] Wgt_6_659,input [WEIGHT_SIZE-1:0] Wgt_6_660,input [WEIGHT_SIZE-1:0] Wgt_6_661,input [WEIGHT_SIZE-1:0] Wgt_6_662,input [WEIGHT_SIZE-1:0] Wgt_6_663,input [WEIGHT_SIZE-1:0] Wgt_6_664,input [WEIGHT_SIZE-1:0] Wgt_6_665,input [WEIGHT_SIZE-1:0] Wgt_6_666,input [WEIGHT_SIZE-1:0] Wgt_6_667,input [WEIGHT_SIZE-1:0] Wgt_6_668,input [WEIGHT_SIZE-1:0] Wgt_6_669,input [WEIGHT_SIZE-1:0] Wgt_6_670,input [WEIGHT_SIZE-1:0] Wgt_6_671,input [WEIGHT_SIZE-1:0] Wgt_6_672,input [WEIGHT_SIZE-1:0] Wgt_6_673,input [WEIGHT_SIZE-1:0] Wgt_6_674,input [WEIGHT_SIZE-1:0] Wgt_6_675,input [WEIGHT_SIZE-1:0] Wgt_6_676,input [WEIGHT_SIZE-1:0] Wgt_6_677,input [WEIGHT_SIZE-1:0] Wgt_6_678,input [WEIGHT_SIZE-1:0] Wgt_6_679,input [WEIGHT_SIZE-1:0] Wgt_6_680,input [WEIGHT_SIZE-1:0] Wgt_6_681,input [WEIGHT_SIZE-1:0] Wgt_6_682,input [WEIGHT_SIZE-1:0] Wgt_6_683,input [WEIGHT_SIZE-1:0] Wgt_6_684,input [WEIGHT_SIZE-1:0] Wgt_6_685,input [WEIGHT_SIZE-1:0] Wgt_6_686,input [WEIGHT_SIZE-1:0] Wgt_6_687,input [WEIGHT_SIZE-1:0] Wgt_6_688,input [WEIGHT_SIZE-1:0] Wgt_6_689,input [WEIGHT_SIZE-1:0] Wgt_6_690,input [WEIGHT_SIZE-1:0] Wgt_6_691,input [WEIGHT_SIZE-1:0] Wgt_6_692,input [WEIGHT_SIZE-1:0] Wgt_6_693,input [WEIGHT_SIZE-1:0] Wgt_6_694,input [WEIGHT_SIZE-1:0] Wgt_6_695,input [WEIGHT_SIZE-1:0] Wgt_6_696,input [WEIGHT_SIZE-1:0] Wgt_6_697,input [WEIGHT_SIZE-1:0] Wgt_6_698,input [WEIGHT_SIZE-1:0] Wgt_6_699,input [WEIGHT_SIZE-1:0] Wgt_6_700,input [WEIGHT_SIZE-1:0] Wgt_6_701,input [WEIGHT_SIZE-1:0] Wgt_6_702,input [WEIGHT_SIZE-1:0] Wgt_6_703,input [WEIGHT_SIZE-1:0] Wgt_6_704,input [WEIGHT_SIZE-1:0] Wgt_6_705,input [WEIGHT_SIZE-1:0] Wgt_6_706,input [WEIGHT_SIZE-1:0] Wgt_6_707,input [WEIGHT_SIZE-1:0] Wgt_6_708,input [WEIGHT_SIZE-1:0] Wgt_6_709,input [WEIGHT_SIZE-1:0] Wgt_6_710,input [WEIGHT_SIZE-1:0] Wgt_6_711,input [WEIGHT_SIZE-1:0] Wgt_6_712,input [WEIGHT_SIZE-1:0] Wgt_6_713,input [WEIGHT_SIZE-1:0] Wgt_6_714,input [WEIGHT_SIZE-1:0] Wgt_6_715,input [WEIGHT_SIZE-1:0] Wgt_6_716,input [WEIGHT_SIZE-1:0] Wgt_6_717,input [WEIGHT_SIZE-1:0] Wgt_6_718,input [WEIGHT_SIZE-1:0] Wgt_6_719,input [WEIGHT_SIZE-1:0] Wgt_6_720,input [WEIGHT_SIZE-1:0] Wgt_6_721,input [WEIGHT_SIZE-1:0] Wgt_6_722,input [WEIGHT_SIZE-1:0] Wgt_6_723,input [WEIGHT_SIZE-1:0] Wgt_6_724,input [WEIGHT_SIZE-1:0] Wgt_6_725,input [WEIGHT_SIZE-1:0] Wgt_6_726,input [WEIGHT_SIZE-1:0] Wgt_6_727,input [WEIGHT_SIZE-1:0] Wgt_6_728,input [WEIGHT_SIZE-1:0] Wgt_6_729,input [WEIGHT_SIZE-1:0] Wgt_6_730,input [WEIGHT_SIZE-1:0] Wgt_6_731,input [WEIGHT_SIZE-1:0] Wgt_6_732,input [WEIGHT_SIZE-1:0] Wgt_6_733,input [WEIGHT_SIZE-1:0] Wgt_6_734,input [WEIGHT_SIZE-1:0] Wgt_6_735,input [WEIGHT_SIZE-1:0] Wgt_6_736,input [WEIGHT_SIZE-1:0] Wgt_6_737,input [WEIGHT_SIZE-1:0] Wgt_6_738,input [WEIGHT_SIZE-1:0] Wgt_6_739,input [WEIGHT_SIZE-1:0] Wgt_6_740,input [WEIGHT_SIZE-1:0] Wgt_6_741,input [WEIGHT_SIZE-1:0] Wgt_6_742,input [WEIGHT_SIZE-1:0] Wgt_6_743,input [WEIGHT_SIZE-1:0] Wgt_6_744,input [WEIGHT_SIZE-1:0] Wgt_6_745,input [WEIGHT_SIZE-1:0] Wgt_6_746,input [WEIGHT_SIZE-1:0] Wgt_6_747,input [WEIGHT_SIZE-1:0] Wgt_6_748,input [WEIGHT_SIZE-1:0] Wgt_6_749,input [WEIGHT_SIZE-1:0] Wgt_6_750,input [WEIGHT_SIZE-1:0] Wgt_6_751,input [WEIGHT_SIZE-1:0] Wgt_6_752,input [WEIGHT_SIZE-1:0] Wgt_6_753,input [WEIGHT_SIZE-1:0] Wgt_6_754,input [WEIGHT_SIZE-1:0] Wgt_6_755,input [WEIGHT_SIZE-1:0] Wgt_6_756,input [WEIGHT_SIZE-1:0] Wgt_6_757,input [WEIGHT_SIZE-1:0] Wgt_6_758,input [WEIGHT_SIZE-1:0] Wgt_6_759,input [WEIGHT_SIZE-1:0] Wgt_6_760,input [WEIGHT_SIZE-1:0] Wgt_6_761,input [WEIGHT_SIZE-1:0] Wgt_6_762,input [WEIGHT_SIZE-1:0] Wgt_6_763,input [WEIGHT_SIZE-1:0] Wgt_6_764,input [WEIGHT_SIZE-1:0] Wgt_6_765,input [WEIGHT_SIZE-1:0] Wgt_6_766,input [WEIGHT_SIZE-1:0] Wgt_6_767,input [WEIGHT_SIZE-1:0] Wgt_6_768,input [WEIGHT_SIZE-1:0] Wgt_6_769,input [WEIGHT_SIZE-1:0] Wgt_6_770,input [WEIGHT_SIZE-1:0] Wgt_6_771,input [WEIGHT_SIZE-1:0] Wgt_6_772,input [WEIGHT_SIZE-1:0] Wgt_6_773,input [WEIGHT_SIZE-1:0] Wgt_6_774,input [WEIGHT_SIZE-1:0] Wgt_6_775,input [WEIGHT_SIZE-1:0] Wgt_6_776,input [WEIGHT_SIZE-1:0] Wgt_6_777,input [WEIGHT_SIZE-1:0] Wgt_6_778,input [WEIGHT_SIZE-1:0] Wgt_6_779,input [WEIGHT_SIZE-1:0] Wgt_6_780,input [WEIGHT_SIZE-1:0] Wgt_6_781,input [WEIGHT_SIZE-1:0] Wgt_6_782,input [WEIGHT_SIZE-1:0] Wgt_6_783,input [WEIGHT_SIZE-1:0] Wgt_6_784,input [WEIGHT_SIZE-1:0] Wgt_7_0,input [WEIGHT_SIZE-1:0] Wgt_7_1,input [WEIGHT_SIZE-1:0] Wgt_7_2,input [WEIGHT_SIZE-1:0] Wgt_7_3,input [WEIGHT_SIZE-1:0] Wgt_7_4,input [WEIGHT_SIZE-1:0] Wgt_7_5,input [WEIGHT_SIZE-1:0] Wgt_7_6,input [WEIGHT_SIZE-1:0] Wgt_7_7,input [WEIGHT_SIZE-1:0] Wgt_7_8,input [WEIGHT_SIZE-1:0] Wgt_7_9,input [WEIGHT_SIZE-1:0] Wgt_7_10,input [WEIGHT_SIZE-1:0] Wgt_7_11,input [WEIGHT_SIZE-1:0] Wgt_7_12,input [WEIGHT_SIZE-1:0] Wgt_7_13,input [WEIGHT_SIZE-1:0] Wgt_7_14,input [WEIGHT_SIZE-1:0] Wgt_7_15,input [WEIGHT_SIZE-1:0] Wgt_7_16,input [WEIGHT_SIZE-1:0] Wgt_7_17,input [WEIGHT_SIZE-1:0] Wgt_7_18,input [WEIGHT_SIZE-1:0] Wgt_7_19,input [WEIGHT_SIZE-1:0] Wgt_7_20,input [WEIGHT_SIZE-1:0] Wgt_7_21,input [WEIGHT_SIZE-1:0] Wgt_7_22,input [WEIGHT_SIZE-1:0] Wgt_7_23,input [WEIGHT_SIZE-1:0] Wgt_7_24,input [WEIGHT_SIZE-1:0] Wgt_7_25,input [WEIGHT_SIZE-1:0] Wgt_7_26,input [WEIGHT_SIZE-1:0] Wgt_7_27,input [WEIGHT_SIZE-1:0] Wgt_7_28,input [WEIGHT_SIZE-1:0] Wgt_7_29,input [WEIGHT_SIZE-1:0] Wgt_7_30,input [WEIGHT_SIZE-1:0] Wgt_7_31,input [WEIGHT_SIZE-1:0] Wgt_7_32,input [WEIGHT_SIZE-1:0] Wgt_7_33,input [WEIGHT_SIZE-1:0] Wgt_7_34,input [WEIGHT_SIZE-1:0] Wgt_7_35,input [WEIGHT_SIZE-1:0] Wgt_7_36,input [WEIGHT_SIZE-1:0] Wgt_7_37,input [WEIGHT_SIZE-1:0] Wgt_7_38,input [WEIGHT_SIZE-1:0] Wgt_7_39,input [WEIGHT_SIZE-1:0] Wgt_7_40,input [WEIGHT_SIZE-1:0] Wgt_7_41,input [WEIGHT_SIZE-1:0] Wgt_7_42,input [WEIGHT_SIZE-1:0] Wgt_7_43,input [WEIGHT_SIZE-1:0] Wgt_7_44,input [WEIGHT_SIZE-1:0] Wgt_7_45,input [WEIGHT_SIZE-1:0] Wgt_7_46,input [WEIGHT_SIZE-1:0] Wgt_7_47,input [WEIGHT_SIZE-1:0] Wgt_7_48,input [WEIGHT_SIZE-1:0] Wgt_7_49,input [WEIGHT_SIZE-1:0] Wgt_7_50,input [WEIGHT_SIZE-1:0] Wgt_7_51,input [WEIGHT_SIZE-1:0] Wgt_7_52,input [WEIGHT_SIZE-1:0] Wgt_7_53,input [WEIGHT_SIZE-1:0] Wgt_7_54,input [WEIGHT_SIZE-1:0] Wgt_7_55,input [WEIGHT_SIZE-1:0] Wgt_7_56,input [WEIGHT_SIZE-1:0] Wgt_7_57,input [WEIGHT_SIZE-1:0] Wgt_7_58,input [WEIGHT_SIZE-1:0] Wgt_7_59,input [WEIGHT_SIZE-1:0] Wgt_7_60,input [WEIGHT_SIZE-1:0] Wgt_7_61,input [WEIGHT_SIZE-1:0] Wgt_7_62,input [WEIGHT_SIZE-1:0] Wgt_7_63,input [WEIGHT_SIZE-1:0] Wgt_7_64,input [WEIGHT_SIZE-1:0] Wgt_7_65,input [WEIGHT_SIZE-1:0] Wgt_7_66,input [WEIGHT_SIZE-1:0] Wgt_7_67,input [WEIGHT_SIZE-1:0] Wgt_7_68,input [WEIGHT_SIZE-1:0] Wgt_7_69,input [WEIGHT_SIZE-1:0] Wgt_7_70,input [WEIGHT_SIZE-1:0] Wgt_7_71,input [WEIGHT_SIZE-1:0] Wgt_7_72,input [WEIGHT_SIZE-1:0] Wgt_7_73,input [WEIGHT_SIZE-1:0] Wgt_7_74,input [WEIGHT_SIZE-1:0] Wgt_7_75,input [WEIGHT_SIZE-1:0] Wgt_7_76,input [WEIGHT_SIZE-1:0] Wgt_7_77,input [WEIGHT_SIZE-1:0] Wgt_7_78,input [WEIGHT_SIZE-1:0] Wgt_7_79,input [WEIGHT_SIZE-1:0] Wgt_7_80,input [WEIGHT_SIZE-1:0] Wgt_7_81,input [WEIGHT_SIZE-1:0] Wgt_7_82,input [WEIGHT_SIZE-1:0] Wgt_7_83,input [WEIGHT_SIZE-1:0] Wgt_7_84,input [WEIGHT_SIZE-1:0] Wgt_7_85,input [WEIGHT_SIZE-1:0] Wgt_7_86,input [WEIGHT_SIZE-1:0] Wgt_7_87,input [WEIGHT_SIZE-1:0] Wgt_7_88,input [WEIGHT_SIZE-1:0] Wgt_7_89,input [WEIGHT_SIZE-1:0] Wgt_7_90,input [WEIGHT_SIZE-1:0] Wgt_7_91,input [WEIGHT_SIZE-1:0] Wgt_7_92,input [WEIGHT_SIZE-1:0] Wgt_7_93,input [WEIGHT_SIZE-1:0] Wgt_7_94,input [WEIGHT_SIZE-1:0] Wgt_7_95,input [WEIGHT_SIZE-1:0] Wgt_7_96,input [WEIGHT_SIZE-1:0] Wgt_7_97,input [WEIGHT_SIZE-1:0] Wgt_7_98,input [WEIGHT_SIZE-1:0] Wgt_7_99,input [WEIGHT_SIZE-1:0] Wgt_7_100,input [WEIGHT_SIZE-1:0] Wgt_7_101,input [WEIGHT_SIZE-1:0] Wgt_7_102,input [WEIGHT_SIZE-1:0] Wgt_7_103,input [WEIGHT_SIZE-1:0] Wgt_7_104,input [WEIGHT_SIZE-1:0] Wgt_7_105,input [WEIGHT_SIZE-1:0] Wgt_7_106,input [WEIGHT_SIZE-1:0] Wgt_7_107,input [WEIGHT_SIZE-1:0] Wgt_7_108,input [WEIGHT_SIZE-1:0] Wgt_7_109,input [WEIGHT_SIZE-1:0] Wgt_7_110,input [WEIGHT_SIZE-1:0] Wgt_7_111,input [WEIGHT_SIZE-1:0] Wgt_7_112,input [WEIGHT_SIZE-1:0] Wgt_7_113,input [WEIGHT_SIZE-1:0] Wgt_7_114,input [WEIGHT_SIZE-1:0] Wgt_7_115,input [WEIGHT_SIZE-1:0] Wgt_7_116,input [WEIGHT_SIZE-1:0] Wgt_7_117,input [WEIGHT_SIZE-1:0] Wgt_7_118,input [WEIGHT_SIZE-1:0] Wgt_7_119,input [WEIGHT_SIZE-1:0] Wgt_7_120,input [WEIGHT_SIZE-1:0] Wgt_7_121,input [WEIGHT_SIZE-1:0] Wgt_7_122,input [WEIGHT_SIZE-1:0] Wgt_7_123,input [WEIGHT_SIZE-1:0] Wgt_7_124,input [WEIGHT_SIZE-1:0] Wgt_7_125,input [WEIGHT_SIZE-1:0] Wgt_7_126,input [WEIGHT_SIZE-1:0] Wgt_7_127,input [WEIGHT_SIZE-1:0] Wgt_7_128,input [WEIGHT_SIZE-1:0] Wgt_7_129,input [WEIGHT_SIZE-1:0] Wgt_7_130,input [WEIGHT_SIZE-1:0] Wgt_7_131,input [WEIGHT_SIZE-1:0] Wgt_7_132,input [WEIGHT_SIZE-1:0] Wgt_7_133,input [WEIGHT_SIZE-1:0] Wgt_7_134,input [WEIGHT_SIZE-1:0] Wgt_7_135,input [WEIGHT_SIZE-1:0] Wgt_7_136,input [WEIGHT_SIZE-1:0] Wgt_7_137,input [WEIGHT_SIZE-1:0] Wgt_7_138,input [WEIGHT_SIZE-1:0] Wgt_7_139,input [WEIGHT_SIZE-1:0] Wgt_7_140,input [WEIGHT_SIZE-1:0] Wgt_7_141,input [WEIGHT_SIZE-1:0] Wgt_7_142,input [WEIGHT_SIZE-1:0] Wgt_7_143,input [WEIGHT_SIZE-1:0] Wgt_7_144,input [WEIGHT_SIZE-1:0] Wgt_7_145,input [WEIGHT_SIZE-1:0] Wgt_7_146,input [WEIGHT_SIZE-1:0] Wgt_7_147,input [WEIGHT_SIZE-1:0] Wgt_7_148,input [WEIGHT_SIZE-1:0] Wgt_7_149,input [WEIGHT_SIZE-1:0] Wgt_7_150,input [WEIGHT_SIZE-1:0] Wgt_7_151,input [WEIGHT_SIZE-1:0] Wgt_7_152,input [WEIGHT_SIZE-1:0] Wgt_7_153,input [WEIGHT_SIZE-1:0] Wgt_7_154,input [WEIGHT_SIZE-1:0] Wgt_7_155,input [WEIGHT_SIZE-1:0] Wgt_7_156,input [WEIGHT_SIZE-1:0] Wgt_7_157,input [WEIGHT_SIZE-1:0] Wgt_7_158,input [WEIGHT_SIZE-1:0] Wgt_7_159,input [WEIGHT_SIZE-1:0] Wgt_7_160,input [WEIGHT_SIZE-1:0] Wgt_7_161,input [WEIGHT_SIZE-1:0] Wgt_7_162,input [WEIGHT_SIZE-1:0] Wgt_7_163,input [WEIGHT_SIZE-1:0] Wgt_7_164,input [WEIGHT_SIZE-1:0] Wgt_7_165,input [WEIGHT_SIZE-1:0] Wgt_7_166,input [WEIGHT_SIZE-1:0] Wgt_7_167,input [WEIGHT_SIZE-1:0] Wgt_7_168,input [WEIGHT_SIZE-1:0] Wgt_7_169,input [WEIGHT_SIZE-1:0] Wgt_7_170,input [WEIGHT_SIZE-1:0] Wgt_7_171,input [WEIGHT_SIZE-1:0] Wgt_7_172,input [WEIGHT_SIZE-1:0] Wgt_7_173,input [WEIGHT_SIZE-1:0] Wgt_7_174,input [WEIGHT_SIZE-1:0] Wgt_7_175,input [WEIGHT_SIZE-1:0] Wgt_7_176,input [WEIGHT_SIZE-1:0] Wgt_7_177,input [WEIGHT_SIZE-1:0] Wgt_7_178,input [WEIGHT_SIZE-1:0] Wgt_7_179,input [WEIGHT_SIZE-1:0] Wgt_7_180,input [WEIGHT_SIZE-1:0] Wgt_7_181,input [WEIGHT_SIZE-1:0] Wgt_7_182,input [WEIGHT_SIZE-1:0] Wgt_7_183,input [WEIGHT_SIZE-1:0] Wgt_7_184,input [WEIGHT_SIZE-1:0] Wgt_7_185,input [WEIGHT_SIZE-1:0] Wgt_7_186,input [WEIGHT_SIZE-1:0] Wgt_7_187,input [WEIGHT_SIZE-1:0] Wgt_7_188,input [WEIGHT_SIZE-1:0] Wgt_7_189,input [WEIGHT_SIZE-1:0] Wgt_7_190,input [WEIGHT_SIZE-1:0] Wgt_7_191,input [WEIGHT_SIZE-1:0] Wgt_7_192,input [WEIGHT_SIZE-1:0] Wgt_7_193,input [WEIGHT_SIZE-1:0] Wgt_7_194,input [WEIGHT_SIZE-1:0] Wgt_7_195,input [WEIGHT_SIZE-1:0] Wgt_7_196,input [WEIGHT_SIZE-1:0] Wgt_7_197,input [WEIGHT_SIZE-1:0] Wgt_7_198,input [WEIGHT_SIZE-1:0] Wgt_7_199,input [WEIGHT_SIZE-1:0] Wgt_7_200,input [WEIGHT_SIZE-1:0] Wgt_7_201,input [WEIGHT_SIZE-1:0] Wgt_7_202,input [WEIGHT_SIZE-1:0] Wgt_7_203,input [WEIGHT_SIZE-1:0] Wgt_7_204,input [WEIGHT_SIZE-1:0] Wgt_7_205,input [WEIGHT_SIZE-1:0] Wgt_7_206,input [WEIGHT_SIZE-1:0] Wgt_7_207,input [WEIGHT_SIZE-1:0] Wgt_7_208,input [WEIGHT_SIZE-1:0] Wgt_7_209,input [WEIGHT_SIZE-1:0] Wgt_7_210,input [WEIGHT_SIZE-1:0] Wgt_7_211,input [WEIGHT_SIZE-1:0] Wgt_7_212,input [WEIGHT_SIZE-1:0] Wgt_7_213,input [WEIGHT_SIZE-1:0] Wgt_7_214,input [WEIGHT_SIZE-1:0] Wgt_7_215,input [WEIGHT_SIZE-1:0] Wgt_7_216,input [WEIGHT_SIZE-1:0] Wgt_7_217,input [WEIGHT_SIZE-1:0] Wgt_7_218,input [WEIGHT_SIZE-1:0] Wgt_7_219,input [WEIGHT_SIZE-1:0] Wgt_7_220,input [WEIGHT_SIZE-1:0] Wgt_7_221,input [WEIGHT_SIZE-1:0] Wgt_7_222,input [WEIGHT_SIZE-1:0] Wgt_7_223,input [WEIGHT_SIZE-1:0] Wgt_7_224,input [WEIGHT_SIZE-1:0] Wgt_7_225,input [WEIGHT_SIZE-1:0] Wgt_7_226,input [WEIGHT_SIZE-1:0] Wgt_7_227,input [WEIGHT_SIZE-1:0] Wgt_7_228,input [WEIGHT_SIZE-1:0] Wgt_7_229,input [WEIGHT_SIZE-1:0] Wgt_7_230,input [WEIGHT_SIZE-1:0] Wgt_7_231,input [WEIGHT_SIZE-1:0] Wgt_7_232,input [WEIGHT_SIZE-1:0] Wgt_7_233,input [WEIGHT_SIZE-1:0] Wgt_7_234,input [WEIGHT_SIZE-1:0] Wgt_7_235,input [WEIGHT_SIZE-1:0] Wgt_7_236,input [WEIGHT_SIZE-1:0] Wgt_7_237,input [WEIGHT_SIZE-1:0] Wgt_7_238,input [WEIGHT_SIZE-1:0] Wgt_7_239,input [WEIGHT_SIZE-1:0] Wgt_7_240,input [WEIGHT_SIZE-1:0] Wgt_7_241,input [WEIGHT_SIZE-1:0] Wgt_7_242,input [WEIGHT_SIZE-1:0] Wgt_7_243,input [WEIGHT_SIZE-1:0] Wgt_7_244,input [WEIGHT_SIZE-1:0] Wgt_7_245,input [WEIGHT_SIZE-1:0] Wgt_7_246,input [WEIGHT_SIZE-1:0] Wgt_7_247,input [WEIGHT_SIZE-1:0] Wgt_7_248,input [WEIGHT_SIZE-1:0] Wgt_7_249,input [WEIGHT_SIZE-1:0] Wgt_7_250,input [WEIGHT_SIZE-1:0] Wgt_7_251,input [WEIGHT_SIZE-1:0] Wgt_7_252,input [WEIGHT_SIZE-1:0] Wgt_7_253,input [WEIGHT_SIZE-1:0] Wgt_7_254,input [WEIGHT_SIZE-1:0] Wgt_7_255,input [WEIGHT_SIZE-1:0] Wgt_7_256,input [WEIGHT_SIZE-1:0] Wgt_7_257,input [WEIGHT_SIZE-1:0] Wgt_7_258,input [WEIGHT_SIZE-1:0] Wgt_7_259,input [WEIGHT_SIZE-1:0] Wgt_7_260,input [WEIGHT_SIZE-1:0] Wgt_7_261,input [WEIGHT_SIZE-1:0] Wgt_7_262,input [WEIGHT_SIZE-1:0] Wgt_7_263,input [WEIGHT_SIZE-1:0] Wgt_7_264,input [WEIGHT_SIZE-1:0] Wgt_7_265,input [WEIGHT_SIZE-1:0] Wgt_7_266,input [WEIGHT_SIZE-1:0] Wgt_7_267,input [WEIGHT_SIZE-1:0] Wgt_7_268,input [WEIGHT_SIZE-1:0] Wgt_7_269,input [WEIGHT_SIZE-1:0] Wgt_7_270,input [WEIGHT_SIZE-1:0] Wgt_7_271,input [WEIGHT_SIZE-1:0] Wgt_7_272,input [WEIGHT_SIZE-1:0] Wgt_7_273,input [WEIGHT_SIZE-1:0] Wgt_7_274,input [WEIGHT_SIZE-1:0] Wgt_7_275,input [WEIGHT_SIZE-1:0] Wgt_7_276,input [WEIGHT_SIZE-1:0] Wgt_7_277,input [WEIGHT_SIZE-1:0] Wgt_7_278,input [WEIGHT_SIZE-1:0] Wgt_7_279,input [WEIGHT_SIZE-1:0] Wgt_7_280,input [WEIGHT_SIZE-1:0] Wgt_7_281,input [WEIGHT_SIZE-1:0] Wgt_7_282,input [WEIGHT_SIZE-1:0] Wgt_7_283,input [WEIGHT_SIZE-1:0] Wgt_7_284,input [WEIGHT_SIZE-1:0] Wgt_7_285,input [WEIGHT_SIZE-1:0] Wgt_7_286,input [WEIGHT_SIZE-1:0] Wgt_7_287,input [WEIGHT_SIZE-1:0] Wgt_7_288,input [WEIGHT_SIZE-1:0] Wgt_7_289,input [WEIGHT_SIZE-1:0] Wgt_7_290,input [WEIGHT_SIZE-1:0] Wgt_7_291,input [WEIGHT_SIZE-1:0] Wgt_7_292,input [WEIGHT_SIZE-1:0] Wgt_7_293,input [WEIGHT_SIZE-1:0] Wgt_7_294,input [WEIGHT_SIZE-1:0] Wgt_7_295,input [WEIGHT_SIZE-1:0] Wgt_7_296,input [WEIGHT_SIZE-1:0] Wgt_7_297,input [WEIGHT_SIZE-1:0] Wgt_7_298,input [WEIGHT_SIZE-1:0] Wgt_7_299,input [WEIGHT_SIZE-1:0] Wgt_7_300,input [WEIGHT_SIZE-1:0] Wgt_7_301,input [WEIGHT_SIZE-1:0] Wgt_7_302,input [WEIGHT_SIZE-1:0] Wgt_7_303,input [WEIGHT_SIZE-1:0] Wgt_7_304,input [WEIGHT_SIZE-1:0] Wgt_7_305,input [WEIGHT_SIZE-1:0] Wgt_7_306,input [WEIGHT_SIZE-1:0] Wgt_7_307,input [WEIGHT_SIZE-1:0] Wgt_7_308,input [WEIGHT_SIZE-1:0] Wgt_7_309,input [WEIGHT_SIZE-1:0] Wgt_7_310,input [WEIGHT_SIZE-1:0] Wgt_7_311,input [WEIGHT_SIZE-1:0] Wgt_7_312,input [WEIGHT_SIZE-1:0] Wgt_7_313,input [WEIGHT_SIZE-1:0] Wgt_7_314,input [WEIGHT_SIZE-1:0] Wgt_7_315,input [WEIGHT_SIZE-1:0] Wgt_7_316,input [WEIGHT_SIZE-1:0] Wgt_7_317,input [WEIGHT_SIZE-1:0] Wgt_7_318,input [WEIGHT_SIZE-1:0] Wgt_7_319,input [WEIGHT_SIZE-1:0] Wgt_7_320,input [WEIGHT_SIZE-1:0] Wgt_7_321,input [WEIGHT_SIZE-1:0] Wgt_7_322,input [WEIGHT_SIZE-1:0] Wgt_7_323,input [WEIGHT_SIZE-1:0] Wgt_7_324,input [WEIGHT_SIZE-1:0] Wgt_7_325,input [WEIGHT_SIZE-1:0] Wgt_7_326,input [WEIGHT_SIZE-1:0] Wgt_7_327,input [WEIGHT_SIZE-1:0] Wgt_7_328,input [WEIGHT_SIZE-1:0] Wgt_7_329,input [WEIGHT_SIZE-1:0] Wgt_7_330,input [WEIGHT_SIZE-1:0] Wgt_7_331,input [WEIGHT_SIZE-1:0] Wgt_7_332,input [WEIGHT_SIZE-1:0] Wgt_7_333,input [WEIGHT_SIZE-1:0] Wgt_7_334,input [WEIGHT_SIZE-1:0] Wgt_7_335,input [WEIGHT_SIZE-1:0] Wgt_7_336,input [WEIGHT_SIZE-1:0] Wgt_7_337,input [WEIGHT_SIZE-1:0] Wgt_7_338,input [WEIGHT_SIZE-1:0] Wgt_7_339,input [WEIGHT_SIZE-1:0] Wgt_7_340,input [WEIGHT_SIZE-1:0] Wgt_7_341,input [WEIGHT_SIZE-1:0] Wgt_7_342,input [WEIGHT_SIZE-1:0] Wgt_7_343,input [WEIGHT_SIZE-1:0] Wgt_7_344,input [WEIGHT_SIZE-1:0] Wgt_7_345,input [WEIGHT_SIZE-1:0] Wgt_7_346,input [WEIGHT_SIZE-1:0] Wgt_7_347,input [WEIGHT_SIZE-1:0] Wgt_7_348,input [WEIGHT_SIZE-1:0] Wgt_7_349,input [WEIGHT_SIZE-1:0] Wgt_7_350,input [WEIGHT_SIZE-1:0] Wgt_7_351,input [WEIGHT_SIZE-1:0] Wgt_7_352,input [WEIGHT_SIZE-1:0] Wgt_7_353,input [WEIGHT_SIZE-1:0] Wgt_7_354,input [WEIGHT_SIZE-1:0] Wgt_7_355,input [WEIGHT_SIZE-1:0] Wgt_7_356,input [WEIGHT_SIZE-1:0] Wgt_7_357,input [WEIGHT_SIZE-1:0] Wgt_7_358,input [WEIGHT_SIZE-1:0] Wgt_7_359,input [WEIGHT_SIZE-1:0] Wgt_7_360,input [WEIGHT_SIZE-1:0] Wgt_7_361,input [WEIGHT_SIZE-1:0] Wgt_7_362,input [WEIGHT_SIZE-1:0] Wgt_7_363,input [WEIGHT_SIZE-1:0] Wgt_7_364,input [WEIGHT_SIZE-1:0] Wgt_7_365,input [WEIGHT_SIZE-1:0] Wgt_7_366,input [WEIGHT_SIZE-1:0] Wgt_7_367,input [WEIGHT_SIZE-1:0] Wgt_7_368,input [WEIGHT_SIZE-1:0] Wgt_7_369,input [WEIGHT_SIZE-1:0] Wgt_7_370,input [WEIGHT_SIZE-1:0] Wgt_7_371,input [WEIGHT_SIZE-1:0] Wgt_7_372,input [WEIGHT_SIZE-1:0] Wgt_7_373,input [WEIGHT_SIZE-1:0] Wgt_7_374,input [WEIGHT_SIZE-1:0] Wgt_7_375,input [WEIGHT_SIZE-1:0] Wgt_7_376,input [WEIGHT_SIZE-1:0] Wgt_7_377,input [WEIGHT_SIZE-1:0] Wgt_7_378,input [WEIGHT_SIZE-1:0] Wgt_7_379,input [WEIGHT_SIZE-1:0] Wgt_7_380,input [WEIGHT_SIZE-1:0] Wgt_7_381,input [WEIGHT_SIZE-1:0] Wgt_7_382,input [WEIGHT_SIZE-1:0] Wgt_7_383,input [WEIGHT_SIZE-1:0] Wgt_7_384,input [WEIGHT_SIZE-1:0] Wgt_7_385,input [WEIGHT_SIZE-1:0] Wgt_7_386,input [WEIGHT_SIZE-1:0] Wgt_7_387,input [WEIGHT_SIZE-1:0] Wgt_7_388,input [WEIGHT_SIZE-1:0] Wgt_7_389,input [WEIGHT_SIZE-1:0] Wgt_7_390,input [WEIGHT_SIZE-1:0] Wgt_7_391,input [WEIGHT_SIZE-1:0] Wgt_7_392,input [WEIGHT_SIZE-1:0] Wgt_7_393,input [WEIGHT_SIZE-1:0] Wgt_7_394,input [WEIGHT_SIZE-1:0] Wgt_7_395,input [WEIGHT_SIZE-1:0] Wgt_7_396,input [WEIGHT_SIZE-1:0] Wgt_7_397,input [WEIGHT_SIZE-1:0] Wgt_7_398,input [WEIGHT_SIZE-1:0] Wgt_7_399,input [WEIGHT_SIZE-1:0] Wgt_7_400,input [WEIGHT_SIZE-1:0] Wgt_7_401,input [WEIGHT_SIZE-1:0] Wgt_7_402,input [WEIGHT_SIZE-1:0] Wgt_7_403,input [WEIGHT_SIZE-1:0] Wgt_7_404,input [WEIGHT_SIZE-1:0] Wgt_7_405,input [WEIGHT_SIZE-1:0] Wgt_7_406,input [WEIGHT_SIZE-1:0] Wgt_7_407,input [WEIGHT_SIZE-1:0] Wgt_7_408,input [WEIGHT_SIZE-1:0] Wgt_7_409,input [WEIGHT_SIZE-1:0] Wgt_7_410,input [WEIGHT_SIZE-1:0] Wgt_7_411,input [WEIGHT_SIZE-1:0] Wgt_7_412,input [WEIGHT_SIZE-1:0] Wgt_7_413,input [WEIGHT_SIZE-1:0] Wgt_7_414,input [WEIGHT_SIZE-1:0] Wgt_7_415,input [WEIGHT_SIZE-1:0] Wgt_7_416,input [WEIGHT_SIZE-1:0] Wgt_7_417,input [WEIGHT_SIZE-1:0] Wgt_7_418,input [WEIGHT_SIZE-1:0] Wgt_7_419,input [WEIGHT_SIZE-1:0] Wgt_7_420,input [WEIGHT_SIZE-1:0] Wgt_7_421,input [WEIGHT_SIZE-1:0] Wgt_7_422,input [WEIGHT_SIZE-1:0] Wgt_7_423,input [WEIGHT_SIZE-1:0] Wgt_7_424,input [WEIGHT_SIZE-1:0] Wgt_7_425,input [WEIGHT_SIZE-1:0] Wgt_7_426,input [WEIGHT_SIZE-1:0] Wgt_7_427,input [WEIGHT_SIZE-1:0] Wgt_7_428,input [WEIGHT_SIZE-1:0] Wgt_7_429,input [WEIGHT_SIZE-1:0] Wgt_7_430,input [WEIGHT_SIZE-1:0] Wgt_7_431,input [WEIGHT_SIZE-1:0] Wgt_7_432,input [WEIGHT_SIZE-1:0] Wgt_7_433,input [WEIGHT_SIZE-1:0] Wgt_7_434,input [WEIGHT_SIZE-1:0] Wgt_7_435,input [WEIGHT_SIZE-1:0] Wgt_7_436,input [WEIGHT_SIZE-1:0] Wgt_7_437,input [WEIGHT_SIZE-1:0] Wgt_7_438,input [WEIGHT_SIZE-1:0] Wgt_7_439,input [WEIGHT_SIZE-1:0] Wgt_7_440,input [WEIGHT_SIZE-1:0] Wgt_7_441,input [WEIGHT_SIZE-1:0] Wgt_7_442,input [WEIGHT_SIZE-1:0] Wgt_7_443,input [WEIGHT_SIZE-1:0] Wgt_7_444,input [WEIGHT_SIZE-1:0] Wgt_7_445,input [WEIGHT_SIZE-1:0] Wgt_7_446,input [WEIGHT_SIZE-1:0] Wgt_7_447,input [WEIGHT_SIZE-1:0] Wgt_7_448,input [WEIGHT_SIZE-1:0] Wgt_7_449,input [WEIGHT_SIZE-1:0] Wgt_7_450,input [WEIGHT_SIZE-1:0] Wgt_7_451,input [WEIGHT_SIZE-1:0] Wgt_7_452,input [WEIGHT_SIZE-1:0] Wgt_7_453,input [WEIGHT_SIZE-1:0] Wgt_7_454,input [WEIGHT_SIZE-1:0] Wgt_7_455,input [WEIGHT_SIZE-1:0] Wgt_7_456,input [WEIGHT_SIZE-1:0] Wgt_7_457,input [WEIGHT_SIZE-1:0] Wgt_7_458,input [WEIGHT_SIZE-1:0] Wgt_7_459,input [WEIGHT_SIZE-1:0] Wgt_7_460,input [WEIGHT_SIZE-1:0] Wgt_7_461,input [WEIGHT_SIZE-1:0] Wgt_7_462,input [WEIGHT_SIZE-1:0] Wgt_7_463,input [WEIGHT_SIZE-1:0] Wgt_7_464,input [WEIGHT_SIZE-1:0] Wgt_7_465,input [WEIGHT_SIZE-1:0] Wgt_7_466,input [WEIGHT_SIZE-1:0] Wgt_7_467,input [WEIGHT_SIZE-1:0] Wgt_7_468,input [WEIGHT_SIZE-1:0] Wgt_7_469,input [WEIGHT_SIZE-1:0] Wgt_7_470,input [WEIGHT_SIZE-1:0] Wgt_7_471,input [WEIGHT_SIZE-1:0] Wgt_7_472,input [WEIGHT_SIZE-1:0] Wgt_7_473,input [WEIGHT_SIZE-1:0] Wgt_7_474,input [WEIGHT_SIZE-1:0] Wgt_7_475,input [WEIGHT_SIZE-1:0] Wgt_7_476,input [WEIGHT_SIZE-1:0] Wgt_7_477,input [WEIGHT_SIZE-1:0] Wgt_7_478,input [WEIGHT_SIZE-1:0] Wgt_7_479,input [WEIGHT_SIZE-1:0] Wgt_7_480,input [WEIGHT_SIZE-1:0] Wgt_7_481,input [WEIGHT_SIZE-1:0] Wgt_7_482,input [WEIGHT_SIZE-1:0] Wgt_7_483,input [WEIGHT_SIZE-1:0] Wgt_7_484,input [WEIGHT_SIZE-1:0] Wgt_7_485,input [WEIGHT_SIZE-1:0] Wgt_7_486,input [WEIGHT_SIZE-1:0] Wgt_7_487,input [WEIGHT_SIZE-1:0] Wgt_7_488,input [WEIGHT_SIZE-1:0] Wgt_7_489,input [WEIGHT_SIZE-1:0] Wgt_7_490,input [WEIGHT_SIZE-1:0] Wgt_7_491,input [WEIGHT_SIZE-1:0] Wgt_7_492,input [WEIGHT_SIZE-1:0] Wgt_7_493,input [WEIGHT_SIZE-1:0] Wgt_7_494,input [WEIGHT_SIZE-1:0] Wgt_7_495,input [WEIGHT_SIZE-1:0] Wgt_7_496,input [WEIGHT_SIZE-1:0] Wgt_7_497,input [WEIGHT_SIZE-1:0] Wgt_7_498,input [WEIGHT_SIZE-1:0] Wgt_7_499,input [WEIGHT_SIZE-1:0] Wgt_7_500,input [WEIGHT_SIZE-1:0] Wgt_7_501,input [WEIGHT_SIZE-1:0] Wgt_7_502,input [WEIGHT_SIZE-1:0] Wgt_7_503,input [WEIGHT_SIZE-1:0] Wgt_7_504,input [WEIGHT_SIZE-1:0] Wgt_7_505,input [WEIGHT_SIZE-1:0] Wgt_7_506,input [WEIGHT_SIZE-1:0] Wgt_7_507,input [WEIGHT_SIZE-1:0] Wgt_7_508,input [WEIGHT_SIZE-1:0] Wgt_7_509,input [WEIGHT_SIZE-1:0] Wgt_7_510,input [WEIGHT_SIZE-1:0] Wgt_7_511,input [WEIGHT_SIZE-1:0] Wgt_7_512,input [WEIGHT_SIZE-1:0] Wgt_7_513,input [WEIGHT_SIZE-1:0] Wgt_7_514,input [WEIGHT_SIZE-1:0] Wgt_7_515,input [WEIGHT_SIZE-1:0] Wgt_7_516,input [WEIGHT_SIZE-1:0] Wgt_7_517,input [WEIGHT_SIZE-1:0] Wgt_7_518,input [WEIGHT_SIZE-1:0] Wgt_7_519,input [WEIGHT_SIZE-1:0] Wgt_7_520,input [WEIGHT_SIZE-1:0] Wgt_7_521,input [WEIGHT_SIZE-1:0] Wgt_7_522,input [WEIGHT_SIZE-1:0] Wgt_7_523,input [WEIGHT_SIZE-1:0] Wgt_7_524,input [WEIGHT_SIZE-1:0] Wgt_7_525,input [WEIGHT_SIZE-1:0] Wgt_7_526,input [WEIGHT_SIZE-1:0] Wgt_7_527,input [WEIGHT_SIZE-1:0] Wgt_7_528,input [WEIGHT_SIZE-1:0] Wgt_7_529,input [WEIGHT_SIZE-1:0] Wgt_7_530,input [WEIGHT_SIZE-1:0] Wgt_7_531,input [WEIGHT_SIZE-1:0] Wgt_7_532,input [WEIGHT_SIZE-1:0] Wgt_7_533,input [WEIGHT_SIZE-1:0] Wgt_7_534,input [WEIGHT_SIZE-1:0] Wgt_7_535,input [WEIGHT_SIZE-1:0] Wgt_7_536,input [WEIGHT_SIZE-1:0] Wgt_7_537,input [WEIGHT_SIZE-1:0] Wgt_7_538,input [WEIGHT_SIZE-1:0] Wgt_7_539,input [WEIGHT_SIZE-1:0] Wgt_7_540,input [WEIGHT_SIZE-1:0] Wgt_7_541,input [WEIGHT_SIZE-1:0] Wgt_7_542,input [WEIGHT_SIZE-1:0] Wgt_7_543,input [WEIGHT_SIZE-1:0] Wgt_7_544,input [WEIGHT_SIZE-1:0] Wgt_7_545,input [WEIGHT_SIZE-1:0] Wgt_7_546,input [WEIGHT_SIZE-1:0] Wgt_7_547,input [WEIGHT_SIZE-1:0] Wgt_7_548,input [WEIGHT_SIZE-1:0] Wgt_7_549,input [WEIGHT_SIZE-1:0] Wgt_7_550,input [WEIGHT_SIZE-1:0] Wgt_7_551,input [WEIGHT_SIZE-1:0] Wgt_7_552,input [WEIGHT_SIZE-1:0] Wgt_7_553,input [WEIGHT_SIZE-1:0] Wgt_7_554,input [WEIGHT_SIZE-1:0] Wgt_7_555,input [WEIGHT_SIZE-1:0] Wgt_7_556,input [WEIGHT_SIZE-1:0] Wgt_7_557,input [WEIGHT_SIZE-1:0] Wgt_7_558,input [WEIGHT_SIZE-1:0] Wgt_7_559,input [WEIGHT_SIZE-1:0] Wgt_7_560,input [WEIGHT_SIZE-1:0] Wgt_7_561,input [WEIGHT_SIZE-1:0] Wgt_7_562,input [WEIGHT_SIZE-1:0] Wgt_7_563,input [WEIGHT_SIZE-1:0] Wgt_7_564,input [WEIGHT_SIZE-1:0] Wgt_7_565,input [WEIGHT_SIZE-1:0] Wgt_7_566,input [WEIGHT_SIZE-1:0] Wgt_7_567,input [WEIGHT_SIZE-1:0] Wgt_7_568,input [WEIGHT_SIZE-1:0] Wgt_7_569,input [WEIGHT_SIZE-1:0] Wgt_7_570,input [WEIGHT_SIZE-1:0] Wgt_7_571,input [WEIGHT_SIZE-1:0] Wgt_7_572,input [WEIGHT_SIZE-1:0] Wgt_7_573,input [WEIGHT_SIZE-1:0] Wgt_7_574,input [WEIGHT_SIZE-1:0] Wgt_7_575,input [WEIGHT_SIZE-1:0] Wgt_7_576,input [WEIGHT_SIZE-1:0] Wgt_7_577,input [WEIGHT_SIZE-1:0] Wgt_7_578,input [WEIGHT_SIZE-1:0] Wgt_7_579,input [WEIGHT_SIZE-1:0] Wgt_7_580,input [WEIGHT_SIZE-1:0] Wgt_7_581,input [WEIGHT_SIZE-1:0] Wgt_7_582,input [WEIGHT_SIZE-1:0] Wgt_7_583,input [WEIGHT_SIZE-1:0] Wgt_7_584,input [WEIGHT_SIZE-1:0] Wgt_7_585,input [WEIGHT_SIZE-1:0] Wgt_7_586,input [WEIGHT_SIZE-1:0] Wgt_7_587,input [WEIGHT_SIZE-1:0] Wgt_7_588,input [WEIGHT_SIZE-1:0] Wgt_7_589,input [WEIGHT_SIZE-1:0] Wgt_7_590,input [WEIGHT_SIZE-1:0] Wgt_7_591,input [WEIGHT_SIZE-1:0] Wgt_7_592,input [WEIGHT_SIZE-1:0] Wgt_7_593,input [WEIGHT_SIZE-1:0] Wgt_7_594,input [WEIGHT_SIZE-1:0] Wgt_7_595,input [WEIGHT_SIZE-1:0] Wgt_7_596,input [WEIGHT_SIZE-1:0] Wgt_7_597,input [WEIGHT_SIZE-1:0] Wgt_7_598,input [WEIGHT_SIZE-1:0] Wgt_7_599,input [WEIGHT_SIZE-1:0] Wgt_7_600,input [WEIGHT_SIZE-1:0] Wgt_7_601,input [WEIGHT_SIZE-1:0] Wgt_7_602,input [WEIGHT_SIZE-1:0] Wgt_7_603,input [WEIGHT_SIZE-1:0] Wgt_7_604,input [WEIGHT_SIZE-1:0] Wgt_7_605,input [WEIGHT_SIZE-1:0] Wgt_7_606,input [WEIGHT_SIZE-1:0] Wgt_7_607,input [WEIGHT_SIZE-1:0] Wgt_7_608,input [WEIGHT_SIZE-1:0] Wgt_7_609,input [WEIGHT_SIZE-1:0] Wgt_7_610,input [WEIGHT_SIZE-1:0] Wgt_7_611,input [WEIGHT_SIZE-1:0] Wgt_7_612,input [WEIGHT_SIZE-1:0] Wgt_7_613,input [WEIGHT_SIZE-1:0] Wgt_7_614,input [WEIGHT_SIZE-1:0] Wgt_7_615,input [WEIGHT_SIZE-1:0] Wgt_7_616,input [WEIGHT_SIZE-1:0] Wgt_7_617,input [WEIGHT_SIZE-1:0] Wgt_7_618,input [WEIGHT_SIZE-1:0] Wgt_7_619,input [WEIGHT_SIZE-1:0] Wgt_7_620,input [WEIGHT_SIZE-1:0] Wgt_7_621,input [WEIGHT_SIZE-1:0] Wgt_7_622,input [WEIGHT_SIZE-1:0] Wgt_7_623,input [WEIGHT_SIZE-1:0] Wgt_7_624,input [WEIGHT_SIZE-1:0] Wgt_7_625,input [WEIGHT_SIZE-1:0] Wgt_7_626,input [WEIGHT_SIZE-1:0] Wgt_7_627,input [WEIGHT_SIZE-1:0] Wgt_7_628,input [WEIGHT_SIZE-1:0] Wgt_7_629,input [WEIGHT_SIZE-1:0] Wgt_7_630,input [WEIGHT_SIZE-1:0] Wgt_7_631,input [WEIGHT_SIZE-1:0] Wgt_7_632,input [WEIGHT_SIZE-1:0] Wgt_7_633,input [WEIGHT_SIZE-1:0] Wgt_7_634,input [WEIGHT_SIZE-1:0] Wgt_7_635,input [WEIGHT_SIZE-1:0] Wgt_7_636,input [WEIGHT_SIZE-1:0] Wgt_7_637,input [WEIGHT_SIZE-1:0] Wgt_7_638,input [WEIGHT_SIZE-1:0] Wgt_7_639,input [WEIGHT_SIZE-1:0] Wgt_7_640,input [WEIGHT_SIZE-1:0] Wgt_7_641,input [WEIGHT_SIZE-1:0] Wgt_7_642,input [WEIGHT_SIZE-1:0] Wgt_7_643,input [WEIGHT_SIZE-1:0] Wgt_7_644,input [WEIGHT_SIZE-1:0] Wgt_7_645,input [WEIGHT_SIZE-1:0] Wgt_7_646,input [WEIGHT_SIZE-1:0] Wgt_7_647,input [WEIGHT_SIZE-1:0] Wgt_7_648,input [WEIGHT_SIZE-1:0] Wgt_7_649,input [WEIGHT_SIZE-1:0] Wgt_7_650,input [WEIGHT_SIZE-1:0] Wgt_7_651,input [WEIGHT_SIZE-1:0] Wgt_7_652,input [WEIGHT_SIZE-1:0] Wgt_7_653,input [WEIGHT_SIZE-1:0] Wgt_7_654,input [WEIGHT_SIZE-1:0] Wgt_7_655,input [WEIGHT_SIZE-1:0] Wgt_7_656,input [WEIGHT_SIZE-1:0] Wgt_7_657,input [WEIGHT_SIZE-1:0] Wgt_7_658,input [WEIGHT_SIZE-1:0] Wgt_7_659,input [WEIGHT_SIZE-1:0] Wgt_7_660,input [WEIGHT_SIZE-1:0] Wgt_7_661,input [WEIGHT_SIZE-1:0] Wgt_7_662,input [WEIGHT_SIZE-1:0] Wgt_7_663,input [WEIGHT_SIZE-1:0] Wgt_7_664,input [WEIGHT_SIZE-1:0] Wgt_7_665,input [WEIGHT_SIZE-1:0] Wgt_7_666,input [WEIGHT_SIZE-1:0] Wgt_7_667,input [WEIGHT_SIZE-1:0] Wgt_7_668,input [WEIGHT_SIZE-1:0] Wgt_7_669,input [WEIGHT_SIZE-1:0] Wgt_7_670,input [WEIGHT_SIZE-1:0] Wgt_7_671,input [WEIGHT_SIZE-1:0] Wgt_7_672,input [WEIGHT_SIZE-1:0] Wgt_7_673,input [WEIGHT_SIZE-1:0] Wgt_7_674,input [WEIGHT_SIZE-1:0] Wgt_7_675,input [WEIGHT_SIZE-1:0] Wgt_7_676,input [WEIGHT_SIZE-1:0] Wgt_7_677,input [WEIGHT_SIZE-1:0] Wgt_7_678,input [WEIGHT_SIZE-1:0] Wgt_7_679,input [WEIGHT_SIZE-1:0] Wgt_7_680,input [WEIGHT_SIZE-1:0] Wgt_7_681,input [WEIGHT_SIZE-1:0] Wgt_7_682,input [WEIGHT_SIZE-1:0] Wgt_7_683,input [WEIGHT_SIZE-1:0] Wgt_7_684,input [WEIGHT_SIZE-1:0] Wgt_7_685,input [WEIGHT_SIZE-1:0] Wgt_7_686,input [WEIGHT_SIZE-1:0] Wgt_7_687,input [WEIGHT_SIZE-1:0] Wgt_7_688,input [WEIGHT_SIZE-1:0] Wgt_7_689,input [WEIGHT_SIZE-1:0] Wgt_7_690,input [WEIGHT_SIZE-1:0] Wgt_7_691,input [WEIGHT_SIZE-1:0] Wgt_7_692,input [WEIGHT_SIZE-1:0] Wgt_7_693,input [WEIGHT_SIZE-1:0] Wgt_7_694,input [WEIGHT_SIZE-1:0] Wgt_7_695,input [WEIGHT_SIZE-1:0] Wgt_7_696,input [WEIGHT_SIZE-1:0] Wgt_7_697,input [WEIGHT_SIZE-1:0] Wgt_7_698,input [WEIGHT_SIZE-1:0] Wgt_7_699,input [WEIGHT_SIZE-1:0] Wgt_7_700,input [WEIGHT_SIZE-1:0] Wgt_7_701,input [WEIGHT_SIZE-1:0] Wgt_7_702,input [WEIGHT_SIZE-1:0] Wgt_7_703,input [WEIGHT_SIZE-1:0] Wgt_7_704,input [WEIGHT_SIZE-1:0] Wgt_7_705,input [WEIGHT_SIZE-1:0] Wgt_7_706,input [WEIGHT_SIZE-1:0] Wgt_7_707,input [WEIGHT_SIZE-1:0] Wgt_7_708,input [WEIGHT_SIZE-1:0] Wgt_7_709,input [WEIGHT_SIZE-1:0] Wgt_7_710,input [WEIGHT_SIZE-1:0] Wgt_7_711,input [WEIGHT_SIZE-1:0] Wgt_7_712,input [WEIGHT_SIZE-1:0] Wgt_7_713,input [WEIGHT_SIZE-1:0] Wgt_7_714,input [WEIGHT_SIZE-1:0] Wgt_7_715,input [WEIGHT_SIZE-1:0] Wgt_7_716,input [WEIGHT_SIZE-1:0] Wgt_7_717,input [WEIGHT_SIZE-1:0] Wgt_7_718,input [WEIGHT_SIZE-1:0] Wgt_7_719,input [WEIGHT_SIZE-1:0] Wgt_7_720,input [WEIGHT_SIZE-1:0] Wgt_7_721,input [WEIGHT_SIZE-1:0] Wgt_7_722,input [WEIGHT_SIZE-1:0] Wgt_7_723,input [WEIGHT_SIZE-1:0] Wgt_7_724,input [WEIGHT_SIZE-1:0] Wgt_7_725,input [WEIGHT_SIZE-1:0] Wgt_7_726,input [WEIGHT_SIZE-1:0] Wgt_7_727,input [WEIGHT_SIZE-1:0] Wgt_7_728,input [WEIGHT_SIZE-1:0] Wgt_7_729,input [WEIGHT_SIZE-1:0] Wgt_7_730,input [WEIGHT_SIZE-1:0] Wgt_7_731,input [WEIGHT_SIZE-1:0] Wgt_7_732,input [WEIGHT_SIZE-1:0] Wgt_7_733,input [WEIGHT_SIZE-1:0] Wgt_7_734,input [WEIGHT_SIZE-1:0] Wgt_7_735,input [WEIGHT_SIZE-1:0] Wgt_7_736,input [WEIGHT_SIZE-1:0] Wgt_7_737,input [WEIGHT_SIZE-1:0] Wgt_7_738,input [WEIGHT_SIZE-1:0] Wgt_7_739,input [WEIGHT_SIZE-1:0] Wgt_7_740,input [WEIGHT_SIZE-1:0] Wgt_7_741,input [WEIGHT_SIZE-1:0] Wgt_7_742,input [WEIGHT_SIZE-1:0] Wgt_7_743,input [WEIGHT_SIZE-1:0] Wgt_7_744,input [WEIGHT_SIZE-1:0] Wgt_7_745,input [WEIGHT_SIZE-1:0] Wgt_7_746,input [WEIGHT_SIZE-1:0] Wgt_7_747,input [WEIGHT_SIZE-1:0] Wgt_7_748,input [WEIGHT_SIZE-1:0] Wgt_7_749,input [WEIGHT_SIZE-1:0] Wgt_7_750,input [WEIGHT_SIZE-1:0] Wgt_7_751,input [WEIGHT_SIZE-1:0] Wgt_7_752,input [WEIGHT_SIZE-1:0] Wgt_7_753,input [WEIGHT_SIZE-1:0] Wgt_7_754,input [WEIGHT_SIZE-1:0] Wgt_7_755,input [WEIGHT_SIZE-1:0] Wgt_7_756,input [WEIGHT_SIZE-1:0] Wgt_7_757,input [WEIGHT_SIZE-1:0] Wgt_7_758,input [WEIGHT_SIZE-1:0] Wgt_7_759,input [WEIGHT_SIZE-1:0] Wgt_7_760,input [WEIGHT_SIZE-1:0] Wgt_7_761,input [WEIGHT_SIZE-1:0] Wgt_7_762,input [WEIGHT_SIZE-1:0] Wgt_7_763,input [WEIGHT_SIZE-1:0] Wgt_7_764,input [WEIGHT_SIZE-1:0] Wgt_7_765,input [WEIGHT_SIZE-1:0] Wgt_7_766,input [WEIGHT_SIZE-1:0] Wgt_7_767,input [WEIGHT_SIZE-1:0] Wgt_7_768,input [WEIGHT_SIZE-1:0] Wgt_7_769,input [WEIGHT_SIZE-1:0] Wgt_7_770,input [WEIGHT_SIZE-1:0] Wgt_7_771,input [WEIGHT_SIZE-1:0] Wgt_7_772,input [WEIGHT_SIZE-1:0] Wgt_7_773,input [WEIGHT_SIZE-1:0] Wgt_7_774,input [WEIGHT_SIZE-1:0] Wgt_7_775,input [WEIGHT_SIZE-1:0] Wgt_7_776,input [WEIGHT_SIZE-1:0] Wgt_7_777,input [WEIGHT_SIZE-1:0] Wgt_7_778,input [WEIGHT_SIZE-1:0] Wgt_7_779,input [WEIGHT_SIZE-1:0] Wgt_7_780,input [WEIGHT_SIZE-1:0] Wgt_7_781,input [WEIGHT_SIZE-1:0] Wgt_7_782,input [WEIGHT_SIZE-1:0] Wgt_7_783,input [WEIGHT_SIZE-1:0] Wgt_7_784,input [WEIGHT_SIZE-1:0] Wgt_8_0,input [WEIGHT_SIZE-1:0] Wgt_8_1,input [WEIGHT_SIZE-1:0] Wgt_8_2,input [WEIGHT_SIZE-1:0] Wgt_8_3,input [WEIGHT_SIZE-1:0] Wgt_8_4,input [WEIGHT_SIZE-1:0] Wgt_8_5,input [WEIGHT_SIZE-1:0] Wgt_8_6,input [WEIGHT_SIZE-1:0] Wgt_8_7,input [WEIGHT_SIZE-1:0] Wgt_8_8,input [WEIGHT_SIZE-1:0] Wgt_8_9,input [WEIGHT_SIZE-1:0] Wgt_8_10,input [WEIGHT_SIZE-1:0] Wgt_8_11,input [WEIGHT_SIZE-1:0] Wgt_8_12,input [WEIGHT_SIZE-1:0] Wgt_8_13,input [WEIGHT_SIZE-1:0] Wgt_8_14,input [WEIGHT_SIZE-1:0] Wgt_8_15,input [WEIGHT_SIZE-1:0] Wgt_8_16,input [WEIGHT_SIZE-1:0] Wgt_8_17,input [WEIGHT_SIZE-1:0] Wgt_8_18,input [WEIGHT_SIZE-1:0] Wgt_8_19,input [WEIGHT_SIZE-1:0] Wgt_8_20,input [WEIGHT_SIZE-1:0] Wgt_8_21,input [WEIGHT_SIZE-1:0] Wgt_8_22,input [WEIGHT_SIZE-1:0] Wgt_8_23,input [WEIGHT_SIZE-1:0] Wgt_8_24,input [WEIGHT_SIZE-1:0] Wgt_8_25,input [WEIGHT_SIZE-1:0] Wgt_8_26,input [WEIGHT_SIZE-1:0] Wgt_8_27,input [WEIGHT_SIZE-1:0] Wgt_8_28,input [WEIGHT_SIZE-1:0] Wgt_8_29,input [WEIGHT_SIZE-1:0] Wgt_8_30,input [WEIGHT_SIZE-1:0] Wgt_8_31,input [WEIGHT_SIZE-1:0] Wgt_8_32,input [WEIGHT_SIZE-1:0] Wgt_8_33,input [WEIGHT_SIZE-1:0] Wgt_8_34,input [WEIGHT_SIZE-1:0] Wgt_8_35,input [WEIGHT_SIZE-1:0] Wgt_8_36,input [WEIGHT_SIZE-1:0] Wgt_8_37,input [WEIGHT_SIZE-1:0] Wgt_8_38,input [WEIGHT_SIZE-1:0] Wgt_8_39,input [WEIGHT_SIZE-1:0] Wgt_8_40,input [WEIGHT_SIZE-1:0] Wgt_8_41,input [WEIGHT_SIZE-1:0] Wgt_8_42,input [WEIGHT_SIZE-1:0] Wgt_8_43,input [WEIGHT_SIZE-1:0] Wgt_8_44,input [WEIGHT_SIZE-1:0] Wgt_8_45,input [WEIGHT_SIZE-1:0] Wgt_8_46,input [WEIGHT_SIZE-1:0] Wgt_8_47,input [WEIGHT_SIZE-1:0] Wgt_8_48,input [WEIGHT_SIZE-1:0] Wgt_8_49,input [WEIGHT_SIZE-1:0] Wgt_8_50,input [WEIGHT_SIZE-1:0] Wgt_8_51,input [WEIGHT_SIZE-1:0] Wgt_8_52,input [WEIGHT_SIZE-1:0] Wgt_8_53,input [WEIGHT_SIZE-1:0] Wgt_8_54,input [WEIGHT_SIZE-1:0] Wgt_8_55,input [WEIGHT_SIZE-1:0] Wgt_8_56,input [WEIGHT_SIZE-1:0] Wgt_8_57,input [WEIGHT_SIZE-1:0] Wgt_8_58,input [WEIGHT_SIZE-1:0] Wgt_8_59,input [WEIGHT_SIZE-1:0] Wgt_8_60,input [WEIGHT_SIZE-1:0] Wgt_8_61,input [WEIGHT_SIZE-1:0] Wgt_8_62,input [WEIGHT_SIZE-1:0] Wgt_8_63,input [WEIGHT_SIZE-1:0] Wgt_8_64,input [WEIGHT_SIZE-1:0] Wgt_8_65,input [WEIGHT_SIZE-1:0] Wgt_8_66,input [WEIGHT_SIZE-1:0] Wgt_8_67,input [WEIGHT_SIZE-1:0] Wgt_8_68,input [WEIGHT_SIZE-1:0] Wgt_8_69,input [WEIGHT_SIZE-1:0] Wgt_8_70,input [WEIGHT_SIZE-1:0] Wgt_8_71,input [WEIGHT_SIZE-1:0] Wgt_8_72,input [WEIGHT_SIZE-1:0] Wgt_8_73,input [WEIGHT_SIZE-1:0] Wgt_8_74,input [WEIGHT_SIZE-1:0] Wgt_8_75,input [WEIGHT_SIZE-1:0] Wgt_8_76,input [WEIGHT_SIZE-1:0] Wgt_8_77,input [WEIGHT_SIZE-1:0] Wgt_8_78,input [WEIGHT_SIZE-1:0] Wgt_8_79,input [WEIGHT_SIZE-1:0] Wgt_8_80,input [WEIGHT_SIZE-1:0] Wgt_8_81,input [WEIGHT_SIZE-1:0] Wgt_8_82,input [WEIGHT_SIZE-1:0] Wgt_8_83,input [WEIGHT_SIZE-1:0] Wgt_8_84,input [WEIGHT_SIZE-1:0] Wgt_8_85,input [WEIGHT_SIZE-1:0] Wgt_8_86,input [WEIGHT_SIZE-1:0] Wgt_8_87,input [WEIGHT_SIZE-1:0] Wgt_8_88,input [WEIGHT_SIZE-1:0] Wgt_8_89,input [WEIGHT_SIZE-1:0] Wgt_8_90,input [WEIGHT_SIZE-1:0] Wgt_8_91,input [WEIGHT_SIZE-1:0] Wgt_8_92,input [WEIGHT_SIZE-1:0] Wgt_8_93,input [WEIGHT_SIZE-1:0] Wgt_8_94,input [WEIGHT_SIZE-1:0] Wgt_8_95,input [WEIGHT_SIZE-1:0] Wgt_8_96,input [WEIGHT_SIZE-1:0] Wgt_8_97,input [WEIGHT_SIZE-1:0] Wgt_8_98,input [WEIGHT_SIZE-1:0] Wgt_8_99,input [WEIGHT_SIZE-1:0] Wgt_8_100,input [WEIGHT_SIZE-1:0] Wgt_8_101,input [WEIGHT_SIZE-1:0] Wgt_8_102,input [WEIGHT_SIZE-1:0] Wgt_8_103,input [WEIGHT_SIZE-1:0] Wgt_8_104,input [WEIGHT_SIZE-1:0] Wgt_8_105,input [WEIGHT_SIZE-1:0] Wgt_8_106,input [WEIGHT_SIZE-1:0] Wgt_8_107,input [WEIGHT_SIZE-1:0] Wgt_8_108,input [WEIGHT_SIZE-1:0] Wgt_8_109,input [WEIGHT_SIZE-1:0] Wgt_8_110,input [WEIGHT_SIZE-1:0] Wgt_8_111,input [WEIGHT_SIZE-1:0] Wgt_8_112,input [WEIGHT_SIZE-1:0] Wgt_8_113,input [WEIGHT_SIZE-1:0] Wgt_8_114,input [WEIGHT_SIZE-1:0] Wgt_8_115,input [WEIGHT_SIZE-1:0] Wgt_8_116,input [WEIGHT_SIZE-1:0] Wgt_8_117,input [WEIGHT_SIZE-1:0] Wgt_8_118,input [WEIGHT_SIZE-1:0] Wgt_8_119,input [WEIGHT_SIZE-1:0] Wgt_8_120,input [WEIGHT_SIZE-1:0] Wgt_8_121,input [WEIGHT_SIZE-1:0] Wgt_8_122,input [WEIGHT_SIZE-1:0] Wgt_8_123,input [WEIGHT_SIZE-1:0] Wgt_8_124,input [WEIGHT_SIZE-1:0] Wgt_8_125,input [WEIGHT_SIZE-1:0] Wgt_8_126,input [WEIGHT_SIZE-1:0] Wgt_8_127,input [WEIGHT_SIZE-1:0] Wgt_8_128,input [WEIGHT_SIZE-1:0] Wgt_8_129,input [WEIGHT_SIZE-1:0] Wgt_8_130,input [WEIGHT_SIZE-1:0] Wgt_8_131,input [WEIGHT_SIZE-1:0] Wgt_8_132,input [WEIGHT_SIZE-1:0] Wgt_8_133,input [WEIGHT_SIZE-1:0] Wgt_8_134,input [WEIGHT_SIZE-1:0] Wgt_8_135,input [WEIGHT_SIZE-1:0] Wgt_8_136,input [WEIGHT_SIZE-1:0] Wgt_8_137,input [WEIGHT_SIZE-1:0] Wgt_8_138,input [WEIGHT_SIZE-1:0] Wgt_8_139,input [WEIGHT_SIZE-1:0] Wgt_8_140,input [WEIGHT_SIZE-1:0] Wgt_8_141,input [WEIGHT_SIZE-1:0] Wgt_8_142,input [WEIGHT_SIZE-1:0] Wgt_8_143,input [WEIGHT_SIZE-1:0] Wgt_8_144,input [WEIGHT_SIZE-1:0] Wgt_8_145,input [WEIGHT_SIZE-1:0] Wgt_8_146,input [WEIGHT_SIZE-1:0] Wgt_8_147,input [WEIGHT_SIZE-1:0] Wgt_8_148,input [WEIGHT_SIZE-1:0] Wgt_8_149,input [WEIGHT_SIZE-1:0] Wgt_8_150,input [WEIGHT_SIZE-1:0] Wgt_8_151,input [WEIGHT_SIZE-1:0] Wgt_8_152,input [WEIGHT_SIZE-1:0] Wgt_8_153,input [WEIGHT_SIZE-1:0] Wgt_8_154,input [WEIGHT_SIZE-1:0] Wgt_8_155,input [WEIGHT_SIZE-1:0] Wgt_8_156,input [WEIGHT_SIZE-1:0] Wgt_8_157,input [WEIGHT_SIZE-1:0] Wgt_8_158,input [WEIGHT_SIZE-1:0] Wgt_8_159,input [WEIGHT_SIZE-1:0] Wgt_8_160,input [WEIGHT_SIZE-1:0] Wgt_8_161,input [WEIGHT_SIZE-1:0] Wgt_8_162,input [WEIGHT_SIZE-1:0] Wgt_8_163,input [WEIGHT_SIZE-1:0] Wgt_8_164,input [WEIGHT_SIZE-1:0] Wgt_8_165,input [WEIGHT_SIZE-1:0] Wgt_8_166,input [WEIGHT_SIZE-1:0] Wgt_8_167,input [WEIGHT_SIZE-1:0] Wgt_8_168,input [WEIGHT_SIZE-1:0] Wgt_8_169,input [WEIGHT_SIZE-1:0] Wgt_8_170,input [WEIGHT_SIZE-1:0] Wgt_8_171,input [WEIGHT_SIZE-1:0] Wgt_8_172,input [WEIGHT_SIZE-1:0] Wgt_8_173,input [WEIGHT_SIZE-1:0] Wgt_8_174,input [WEIGHT_SIZE-1:0] Wgt_8_175,input [WEIGHT_SIZE-1:0] Wgt_8_176,input [WEIGHT_SIZE-1:0] Wgt_8_177,input [WEIGHT_SIZE-1:0] Wgt_8_178,input [WEIGHT_SIZE-1:0] Wgt_8_179,input [WEIGHT_SIZE-1:0] Wgt_8_180,input [WEIGHT_SIZE-1:0] Wgt_8_181,input [WEIGHT_SIZE-1:0] Wgt_8_182,input [WEIGHT_SIZE-1:0] Wgt_8_183,input [WEIGHT_SIZE-1:0] Wgt_8_184,input [WEIGHT_SIZE-1:0] Wgt_8_185,input [WEIGHT_SIZE-1:0] Wgt_8_186,input [WEIGHT_SIZE-1:0] Wgt_8_187,input [WEIGHT_SIZE-1:0] Wgt_8_188,input [WEIGHT_SIZE-1:0] Wgt_8_189,input [WEIGHT_SIZE-1:0] Wgt_8_190,input [WEIGHT_SIZE-1:0] Wgt_8_191,input [WEIGHT_SIZE-1:0] Wgt_8_192,input [WEIGHT_SIZE-1:0] Wgt_8_193,input [WEIGHT_SIZE-1:0] Wgt_8_194,input [WEIGHT_SIZE-1:0] Wgt_8_195,input [WEIGHT_SIZE-1:0] Wgt_8_196,input [WEIGHT_SIZE-1:0] Wgt_8_197,input [WEIGHT_SIZE-1:0] Wgt_8_198,input [WEIGHT_SIZE-1:0] Wgt_8_199,input [WEIGHT_SIZE-1:0] Wgt_8_200,input [WEIGHT_SIZE-1:0] Wgt_8_201,input [WEIGHT_SIZE-1:0] Wgt_8_202,input [WEIGHT_SIZE-1:0] Wgt_8_203,input [WEIGHT_SIZE-1:0] Wgt_8_204,input [WEIGHT_SIZE-1:0] Wgt_8_205,input [WEIGHT_SIZE-1:0] Wgt_8_206,input [WEIGHT_SIZE-1:0] Wgt_8_207,input [WEIGHT_SIZE-1:0] Wgt_8_208,input [WEIGHT_SIZE-1:0] Wgt_8_209,input [WEIGHT_SIZE-1:0] Wgt_8_210,input [WEIGHT_SIZE-1:0] Wgt_8_211,input [WEIGHT_SIZE-1:0] Wgt_8_212,input [WEIGHT_SIZE-1:0] Wgt_8_213,input [WEIGHT_SIZE-1:0] Wgt_8_214,input [WEIGHT_SIZE-1:0] Wgt_8_215,input [WEIGHT_SIZE-1:0] Wgt_8_216,input [WEIGHT_SIZE-1:0] Wgt_8_217,input [WEIGHT_SIZE-1:0] Wgt_8_218,input [WEIGHT_SIZE-1:0] Wgt_8_219,input [WEIGHT_SIZE-1:0] Wgt_8_220,input [WEIGHT_SIZE-1:0] Wgt_8_221,input [WEIGHT_SIZE-1:0] Wgt_8_222,input [WEIGHT_SIZE-1:0] Wgt_8_223,input [WEIGHT_SIZE-1:0] Wgt_8_224,input [WEIGHT_SIZE-1:0] Wgt_8_225,input [WEIGHT_SIZE-1:0] Wgt_8_226,input [WEIGHT_SIZE-1:0] Wgt_8_227,input [WEIGHT_SIZE-1:0] Wgt_8_228,input [WEIGHT_SIZE-1:0] Wgt_8_229,input [WEIGHT_SIZE-1:0] Wgt_8_230,input [WEIGHT_SIZE-1:0] Wgt_8_231,input [WEIGHT_SIZE-1:0] Wgt_8_232,input [WEIGHT_SIZE-1:0] Wgt_8_233,input [WEIGHT_SIZE-1:0] Wgt_8_234,input [WEIGHT_SIZE-1:0] Wgt_8_235,input [WEIGHT_SIZE-1:0] Wgt_8_236,input [WEIGHT_SIZE-1:0] Wgt_8_237,input [WEIGHT_SIZE-1:0] Wgt_8_238,input [WEIGHT_SIZE-1:0] Wgt_8_239,input [WEIGHT_SIZE-1:0] Wgt_8_240,input [WEIGHT_SIZE-1:0] Wgt_8_241,input [WEIGHT_SIZE-1:0] Wgt_8_242,input [WEIGHT_SIZE-1:0] Wgt_8_243,input [WEIGHT_SIZE-1:0] Wgt_8_244,input [WEIGHT_SIZE-1:0] Wgt_8_245,input [WEIGHT_SIZE-1:0] Wgt_8_246,input [WEIGHT_SIZE-1:0] Wgt_8_247,input [WEIGHT_SIZE-1:0] Wgt_8_248,input [WEIGHT_SIZE-1:0] Wgt_8_249,input [WEIGHT_SIZE-1:0] Wgt_8_250,input [WEIGHT_SIZE-1:0] Wgt_8_251,input [WEIGHT_SIZE-1:0] Wgt_8_252,input [WEIGHT_SIZE-1:0] Wgt_8_253,input [WEIGHT_SIZE-1:0] Wgt_8_254,input [WEIGHT_SIZE-1:0] Wgt_8_255,input [WEIGHT_SIZE-1:0] Wgt_8_256,input [WEIGHT_SIZE-1:0] Wgt_8_257,input [WEIGHT_SIZE-1:0] Wgt_8_258,input [WEIGHT_SIZE-1:0] Wgt_8_259,input [WEIGHT_SIZE-1:0] Wgt_8_260,input [WEIGHT_SIZE-1:0] Wgt_8_261,input [WEIGHT_SIZE-1:0] Wgt_8_262,input [WEIGHT_SIZE-1:0] Wgt_8_263,input [WEIGHT_SIZE-1:0] Wgt_8_264,input [WEIGHT_SIZE-1:0] Wgt_8_265,input [WEIGHT_SIZE-1:0] Wgt_8_266,input [WEIGHT_SIZE-1:0] Wgt_8_267,input [WEIGHT_SIZE-1:0] Wgt_8_268,input [WEIGHT_SIZE-1:0] Wgt_8_269,input [WEIGHT_SIZE-1:0] Wgt_8_270,input [WEIGHT_SIZE-1:0] Wgt_8_271,input [WEIGHT_SIZE-1:0] Wgt_8_272,input [WEIGHT_SIZE-1:0] Wgt_8_273,input [WEIGHT_SIZE-1:0] Wgt_8_274,input [WEIGHT_SIZE-1:0] Wgt_8_275,input [WEIGHT_SIZE-1:0] Wgt_8_276,input [WEIGHT_SIZE-1:0] Wgt_8_277,input [WEIGHT_SIZE-1:0] Wgt_8_278,input [WEIGHT_SIZE-1:0] Wgt_8_279,input [WEIGHT_SIZE-1:0] Wgt_8_280,input [WEIGHT_SIZE-1:0] Wgt_8_281,input [WEIGHT_SIZE-1:0] Wgt_8_282,input [WEIGHT_SIZE-1:0] Wgt_8_283,input [WEIGHT_SIZE-1:0] Wgt_8_284,input [WEIGHT_SIZE-1:0] Wgt_8_285,input [WEIGHT_SIZE-1:0] Wgt_8_286,input [WEIGHT_SIZE-1:0] Wgt_8_287,input [WEIGHT_SIZE-1:0] Wgt_8_288,input [WEIGHT_SIZE-1:0] Wgt_8_289,input [WEIGHT_SIZE-1:0] Wgt_8_290,input [WEIGHT_SIZE-1:0] Wgt_8_291,input [WEIGHT_SIZE-1:0] Wgt_8_292,input [WEIGHT_SIZE-1:0] Wgt_8_293,input [WEIGHT_SIZE-1:0] Wgt_8_294,input [WEIGHT_SIZE-1:0] Wgt_8_295,input [WEIGHT_SIZE-1:0] Wgt_8_296,input [WEIGHT_SIZE-1:0] Wgt_8_297,input [WEIGHT_SIZE-1:0] Wgt_8_298,input [WEIGHT_SIZE-1:0] Wgt_8_299,input [WEIGHT_SIZE-1:0] Wgt_8_300,input [WEIGHT_SIZE-1:0] Wgt_8_301,input [WEIGHT_SIZE-1:0] Wgt_8_302,input [WEIGHT_SIZE-1:0] Wgt_8_303,input [WEIGHT_SIZE-1:0] Wgt_8_304,input [WEIGHT_SIZE-1:0] Wgt_8_305,input [WEIGHT_SIZE-1:0] Wgt_8_306,input [WEIGHT_SIZE-1:0] Wgt_8_307,input [WEIGHT_SIZE-1:0] Wgt_8_308,input [WEIGHT_SIZE-1:0] Wgt_8_309,input [WEIGHT_SIZE-1:0] Wgt_8_310,input [WEIGHT_SIZE-1:0] Wgt_8_311,input [WEIGHT_SIZE-1:0] Wgt_8_312,input [WEIGHT_SIZE-1:0] Wgt_8_313,input [WEIGHT_SIZE-1:0] Wgt_8_314,input [WEIGHT_SIZE-1:0] Wgt_8_315,input [WEIGHT_SIZE-1:0] Wgt_8_316,input [WEIGHT_SIZE-1:0] Wgt_8_317,input [WEIGHT_SIZE-1:0] Wgt_8_318,input [WEIGHT_SIZE-1:0] Wgt_8_319,input [WEIGHT_SIZE-1:0] Wgt_8_320,input [WEIGHT_SIZE-1:0] Wgt_8_321,input [WEIGHT_SIZE-1:0] Wgt_8_322,input [WEIGHT_SIZE-1:0] Wgt_8_323,input [WEIGHT_SIZE-1:0] Wgt_8_324,input [WEIGHT_SIZE-1:0] Wgt_8_325,input [WEIGHT_SIZE-1:0] Wgt_8_326,input [WEIGHT_SIZE-1:0] Wgt_8_327,input [WEIGHT_SIZE-1:0] Wgt_8_328,input [WEIGHT_SIZE-1:0] Wgt_8_329,input [WEIGHT_SIZE-1:0] Wgt_8_330,input [WEIGHT_SIZE-1:0] Wgt_8_331,input [WEIGHT_SIZE-1:0] Wgt_8_332,input [WEIGHT_SIZE-1:0] Wgt_8_333,input [WEIGHT_SIZE-1:0] Wgt_8_334,input [WEIGHT_SIZE-1:0] Wgt_8_335,input [WEIGHT_SIZE-1:0] Wgt_8_336,input [WEIGHT_SIZE-1:0] Wgt_8_337,input [WEIGHT_SIZE-1:0] Wgt_8_338,input [WEIGHT_SIZE-1:0] Wgt_8_339,input [WEIGHT_SIZE-1:0] Wgt_8_340,input [WEIGHT_SIZE-1:0] Wgt_8_341,input [WEIGHT_SIZE-1:0] Wgt_8_342,input [WEIGHT_SIZE-1:0] Wgt_8_343,input [WEIGHT_SIZE-1:0] Wgt_8_344,input [WEIGHT_SIZE-1:0] Wgt_8_345,input [WEIGHT_SIZE-1:0] Wgt_8_346,input [WEIGHT_SIZE-1:0] Wgt_8_347,input [WEIGHT_SIZE-1:0] Wgt_8_348,input [WEIGHT_SIZE-1:0] Wgt_8_349,input [WEIGHT_SIZE-1:0] Wgt_8_350,input [WEIGHT_SIZE-1:0] Wgt_8_351,input [WEIGHT_SIZE-1:0] Wgt_8_352,input [WEIGHT_SIZE-1:0] Wgt_8_353,input [WEIGHT_SIZE-1:0] Wgt_8_354,input [WEIGHT_SIZE-1:0] Wgt_8_355,input [WEIGHT_SIZE-1:0] Wgt_8_356,input [WEIGHT_SIZE-1:0] Wgt_8_357,input [WEIGHT_SIZE-1:0] Wgt_8_358,input [WEIGHT_SIZE-1:0] Wgt_8_359,input [WEIGHT_SIZE-1:0] Wgt_8_360,input [WEIGHT_SIZE-1:0] Wgt_8_361,input [WEIGHT_SIZE-1:0] Wgt_8_362,input [WEIGHT_SIZE-1:0] Wgt_8_363,input [WEIGHT_SIZE-1:0] Wgt_8_364,input [WEIGHT_SIZE-1:0] Wgt_8_365,input [WEIGHT_SIZE-1:0] Wgt_8_366,input [WEIGHT_SIZE-1:0] Wgt_8_367,input [WEIGHT_SIZE-1:0] Wgt_8_368,input [WEIGHT_SIZE-1:0] Wgt_8_369,input [WEIGHT_SIZE-1:0] Wgt_8_370,input [WEIGHT_SIZE-1:0] Wgt_8_371,input [WEIGHT_SIZE-1:0] Wgt_8_372,input [WEIGHT_SIZE-1:0] Wgt_8_373,input [WEIGHT_SIZE-1:0] Wgt_8_374,input [WEIGHT_SIZE-1:0] Wgt_8_375,input [WEIGHT_SIZE-1:0] Wgt_8_376,input [WEIGHT_SIZE-1:0] Wgt_8_377,input [WEIGHT_SIZE-1:0] Wgt_8_378,input [WEIGHT_SIZE-1:0] Wgt_8_379,input [WEIGHT_SIZE-1:0] Wgt_8_380,input [WEIGHT_SIZE-1:0] Wgt_8_381,input [WEIGHT_SIZE-1:0] Wgt_8_382,input [WEIGHT_SIZE-1:0] Wgt_8_383,input [WEIGHT_SIZE-1:0] Wgt_8_384,input [WEIGHT_SIZE-1:0] Wgt_8_385,input [WEIGHT_SIZE-1:0] Wgt_8_386,input [WEIGHT_SIZE-1:0] Wgt_8_387,input [WEIGHT_SIZE-1:0] Wgt_8_388,input [WEIGHT_SIZE-1:0] Wgt_8_389,input [WEIGHT_SIZE-1:0] Wgt_8_390,input [WEIGHT_SIZE-1:0] Wgt_8_391,input [WEIGHT_SIZE-1:0] Wgt_8_392,input [WEIGHT_SIZE-1:0] Wgt_8_393,input [WEIGHT_SIZE-1:0] Wgt_8_394,input [WEIGHT_SIZE-1:0] Wgt_8_395,input [WEIGHT_SIZE-1:0] Wgt_8_396,input [WEIGHT_SIZE-1:0] Wgt_8_397,input [WEIGHT_SIZE-1:0] Wgt_8_398,input [WEIGHT_SIZE-1:0] Wgt_8_399,input [WEIGHT_SIZE-1:0] Wgt_8_400,input [WEIGHT_SIZE-1:0] Wgt_8_401,input [WEIGHT_SIZE-1:0] Wgt_8_402,input [WEIGHT_SIZE-1:0] Wgt_8_403,input [WEIGHT_SIZE-1:0] Wgt_8_404,input [WEIGHT_SIZE-1:0] Wgt_8_405,input [WEIGHT_SIZE-1:0] Wgt_8_406,input [WEIGHT_SIZE-1:0] Wgt_8_407,input [WEIGHT_SIZE-1:0] Wgt_8_408,input [WEIGHT_SIZE-1:0] Wgt_8_409,input [WEIGHT_SIZE-1:0] Wgt_8_410,input [WEIGHT_SIZE-1:0] Wgt_8_411,input [WEIGHT_SIZE-1:0] Wgt_8_412,input [WEIGHT_SIZE-1:0] Wgt_8_413,input [WEIGHT_SIZE-1:0] Wgt_8_414,input [WEIGHT_SIZE-1:0] Wgt_8_415,input [WEIGHT_SIZE-1:0] Wgt_8_416,input [WEIGHT_SIZE-1:0] Wgt_8_417,input [WEIGHT_SIZE-1:0] Wgt_8_418,input [WEIGHT_SIZE-1:0] Wgt_8_419,input [WEIGHT_SIZE-1:0] Wgt_8_420,input [WEIGHT_SIZE-1:0] Wgt_8_421,input [WEIGHT_SIZE-1:0] Wgt_8_422,input [WEIGHT_SIZE-1:0] Wgt_8_423,input [WEIGHT_SIZE-1:0] Wgt_8_424,input [WEIGHT_SIZE-1:0] Wgt_8_425,input [WEIGHT_SIZE-1:0] Wgt_8_426,input [WEIGHT_SIZE-1:0] Wgt_8_427,input [WEIGHT_SIZE-1:0] Wgt_8_428,input [WEIGHT_SIZE-1:0] Wgt_8_429,input [WEIGHT_SIZE-1:0] Wgt_8_430,input [WEIGHT_SIZE-1:0] Wgt_8_431,input [WEIGHT_SIZE-1:0] Wgt_8_432,input [WEIGHT_SIZE-1:0] Wgt_8_433,input [WEIGHT_SIZE-1:0] Wgt_8_434,input [WEIGHT_SIZE-1:0] Wgt_8_435,input [WEIGHT_SIZE-1:0] Wgt_8_436,input [WEIGHT_SIZE-1:0] Wgt_8_437,input [WEIGHT_SIZE-1:0] Wgt_8_438,input [WEIGHT_SIZE-1:0] Wgt_8_439,input [WEIGHT_SIZE-1:0] Wgt_8_440,input [WEIGHT_SIZE-1:0] Wgt_8_441,input [WEIGHT_SIZE-1:0] Wgt_8_442,input [WEIGHT_SIZE-1:0] Wgt_8_443,input [WEIGHT_SIZE-1:0] Wgt_8_444,input [WEIGHT_SIZE-1:0] Wgt_8_445,input [WEIGHT_SIZE-1:0] Wgt_8_446,input [WEIGHT_SIZE-1:0] Wgt_8_447,input [WEIGHT_SIZE-1:0] Wgt_8_448,input [WEIGHT_SIZE-1:0] Wgt_8_449,input [WEIGHT_SIZE-1:0] Wgt_8_450,input [WEIGHT_SIZE-1:0] Wgt_8_451,input [WEIGHT_SIZE-1:0] Wgt_8_452,input [WEIGHT_SIZE-1:0] Wgt_8_453,input [WEIGHT_SIZE-1:0] Wgt_8_454,input [WEIGHT_SIZE-1:0] Wgt_8_455,input [WEIGHT_SIZE-1:0] Wgt_8_456,input [WEIGHT_SIZE-1:0] Wgt_8_457,input [WEIGHT_SIZE-1:0] Wgt_8_458,input [WEIGHT_SIZE-1:0] Wgt_8_459,input [WEIGHT_SIZE-1:0] Wgt_8_460,input [WEIGHT_SIZE-1:0] Wgt_8_461,input [WEIGHT_SIZE-1:0] Wgt_8_462,input [WEIGHT_SIZE-1:0] Wgt_8_463,input [WEIGHT_SIZE-1:0] Wgt_8_464,input [WEIGHT_SIZE-1:0] Wgt_8_465,input [WEIGHT_SIZE-1:0] Wgt_8_466,input [WEIGHT_SIZE-1:0] Wgt_8_467,input [WEIGHT_SIZE-1:0] Wgt_8_468,input [WEIGHT_SIZE-1:0] Wgt_8_469,input [WEIGHT_SIZE-1:0] Wgt_8_470,input [WEIGHT_SIZE-1:0] Wgt_8_471,input [WEIGHT_SIZE-1:0] Wgt_8_472,input [WEIGHT_SIZE-1:0] Wgt_8_473,input [WEIGHT_SIZE-1:0] Wgt_8_474,input [WEIGHT_SIZE-1:0] Wgt_8_475,input [WEIGHT_SIZE-1:0] Wgt_8_476,input [WEIGHT_SIZE-1:0] Wgt_8_477,input [WEIGHT_SIZE-1:0] Wgt_8_478,input [WEIGHT_SIZE-1:0] Wgt_8_479,input [WEIGHT_SIZE-1:0] Wgt_8_480,input [WEIGHT_SIZE-1:0] Wgt_8_481,input [WEIGHT_SIZE-1:0] Wgt_8_482,input [WEIGHT_SIZE-1:0] Wgt_8_483,input [WEIGHT_SIZE-1:0] Wgt_8_484,input [WEIGHT_SIZE-1:0] Wgt_8_485,input [WEIGHT_SIZE-1:0] Wgt_8_486,input [WEIGHT_SIZE-1:0] Wgt_8_487,input [WEIGHT_SIZE-1:0] Wgt_8_488,input [WEIGHT_SIZE-1:0] Wgt_8_489,input [WEIGHT_SIZE-1:0] Wgt_8_490,input [WEIGHT_SIZE-1:0] Wgt_8_491,input [WEIGHT_SIZE-1:0] Wgt_8_492,input [WEIGHT_SIZE-1:0] Wgt_8_493,input [WEIGHT_SIZE-1:0] Wgt_8_494,input [WEIGHT_SIZE-1:0] Wgt_8_495,input [WEIGHT_SIZE-1:0] Wgt_8_496,input [WEIGHT_SIZE-1:0] Wgt_8_497,input [WEIGHT_SIZE-1:0] Wgt_8_498,input [WEIGHT_SIZE-1:0] Wgt_8_499,input [WEIGHT_SIZE-1:0] Wgt_8_500,input [WEIGHT_SIZE-1:0] Wgt_8_501,input [WEIGHT_SIZE-1:0] Wgt_8_502,input [WEIGHT_SIZE-1:0] Wgt_8_503,input [WEIGHT_SIZE-1:0] Wgt_8_504,input [WEIGHT_SIZE-1:0] Wgt_8_505,input [WEIGHT_SIZE-1:0] Wgt_8_506,input [WEIGHT_SIZE-1:0] Wgt_8_507,input [WEIGHT_SIZE-1:0] Wgt_8_508,input [WEIGHT_SIZE-1:0] Wgt_8_509,input [WEIGHT_SIZE-1:0] Wgt_8_510,input [WEIGHT_SIZE-1:0] Wgt_8_511,input [WEIGHT_SIZE-1:0] Wgt_8_512,input [WEIGHT_SIZE-1:0] Wgt_8_513,input [WEIGHT_SIZE-1:0] Wgt_8_514,input [WEIGHT_SIZE-1:0] Wgt_8_515,input [WEIGHT_SIZE-1:0] Wgt_8_516,input [WEIGHT_SIZE-1:0] Wgt_8_517,input [WEIGHT_SIZE-1:0] Wgt_8_518,input [WEIGHT_SIZE-1:0] Wgt_8_519,input [WEIGHT_SIZE-1:0] Wgt_8_520,input [WEIGHT_SIZE-1:0] Wgt_8_521,input [WEIGHT_SIZE-1:0] Wgt_8_522,input [WEIGHT_SIZE-1:0] Wgt_8_523,input [WEIGHT_SIZE-1:0] Wgt_8_524,input [WEIGHT_SIZE-1:0] Wgt_8_525,input [WEIGHT_SIZE-1:0] Wgt_8_526,input [WEIGHT_SIZE-1:0] Wgt_8_527,input [WEIGHT_SIZE-1:0] Wgt_8_528,input [WEIGHT_SIZE-1:0] Wgt_8_529,input [WEIGHT_SIZE-1:0] Wgt_8_530,input [WEIGHT_SIZE-1:0] Wgt_8_531,input [WEIGHT_SIZE-1:0] Wgt_8_532,input [WEIGHT_SIZE-1:0] Wgt_8_533,input [WEIGHT_SIZE-1:0] Wgt_8_534,input [WEIGHT_SIZE-1:0] Wgt_8_535,input [WEIGHT_SIZE-1:0] Wgt_8_536,input [WEIGHT_SIZE-1:0] Wgt_8_537,input [WEIGHT_SIZE-1:0] Wgt_8_538,input [WEIGHT_SIZE-1:0] Wgt_8_539,input [WEIGHT_SIZE-1:0] Wgt_8_540,input [WEIGHT_SIZE-1:0] Wgt_8_541,input [WEIGHT_SIZE-1:0] Wgt_8_542,input [WEIGHT_SIZE-1:0] Wgt_8_543,input [WEIGHT_SIZE-1:0] Wgt_8_544,input [WEIGHT_SIZE-1:0] Wgt_8_545,input [WEIGHT_SIZE-1:0] Wgt_8_546,input [WEIGHT_SIZE-1:0] Wgt_8_547,input [WEIGHT_SIZE-1:0] Wgt_8_548,input [WEIGHT_SIZE-1:0] Wgt_8_549,input [WEIGHT_SIZE-1:0] Wgt_8_550,input [WEIGHT_SIZE-1:0] Wgt_8_551,input [WEIGHT_SIZE-1:0] Wgt_8_552,input [WEIGHT_SIZE-1:0] Wgt_8_553,input [WEIGHT_SIZE-1:0] Wgt_8_554,input [WEIGHT_SIZE-1:0] Wgt_8_555,input [WEIGHT_SIZE-1:0] Wgt_8_556,input [WEIGHT_SIZE-1:0] Wgt_8_557,input [WEIGHT_SIZE-1:0] Wgt_8_558,input [WEIGHT_SIZE-1:0] Wgt_8_559,input [WEIGHT_SIZE-1:0] Wgt_8_560,input [WEIGHT_SIZE-1:0] Wgt_8_561,input [WEIGHT_SIZE-1:0] Wgt_8_562,input [WEIGHT_SIZE-1:0] Wgt_8_563,input [WEIGHT_SIZE-1:0] Wgt_8_564,input [WEIGHT_SIZE-1:0] Wgt_8_565,input [WEIGHT_SIZE-1:0] Wgt_8_566,input [WEIGHT_SIZE-1:0] Wgt_8_567,input [WEIGHT_SIZE-1:0] Wgt_8_568,input [WEIGHT_SIZE-1:0] Wgt_8_569,input [WEIGHT_SIZE-1:0] Wgt_8_570,input [WEIGHT_SIZE-1:0] Wgt_8_571,input [WEIGHT_SIZE-1:0] Wgt_8_572,input [WEIGHT_SIZE-1:0] Wgt_8_573,input [WEIGHT_SIZE-1:0] Wgt_8_574,input [WEIGHT_SIZE-1:0] Wgt_8_575,input [WEIGHT_SIZE-1:0] Wgt_8_576,input [WEIGHT_SIZE-1:0] Wgt_8_577,input [WEIGHT_SIZE-1:0] Wgt_8_578,input [WEIGHT_SIZE-1:0] Wgt_8_579,input [WEIGHT_SIZE-1:0] Wgt_8_580,input [WEIGHT_SIZE-1:0] Wgt_8_581,input [WEIGHT_SIZE-1:0] Wgt_8_582,input [WEIGHT_SIZE-1:0] Wgt_8_583,input [WEIGHT_SIZE-1:0] Wgt_8_584,input [WEIGHT_SIZE-1:0] Wgt_8_585,input [WEIGHT_SIZE-1:0] Wgt_8_586,input [WEIGHT_SIZE-1:0] Wgt_8_587,input [WEIGHT_SIZE-1:0] Wgt_8_588,input [WEIGHT_SIZE-1:0] Wgt_8_589,input [WEIGHT_SIZE-1:0] Wgt_8_590,input [WEIGHT_SIZE-1:0] Wgt_8_591,input [WEIGHT_SIZE-1:0] Wgt_8_592,input [WEIGHT_SIZE-1:0] Wgt_8_593,input [WEIGHT_SIZE-1:0] Wgt_8_594,input [WEIGHT_SIZE-1:0] Wgt_8_595,input [WEIGHT_SIZE-1:0] Wgt_8_596,input [WEIGHT_SIZE-1:0] Wgt_8_597,input [WEIGHT_SIZE-1:0] Wgt_8_598,input [WEIGHT_SIZE-1:0] Wgt_8_599,input [WEIGHT_SIZE-1:0] Wgt_8_600,input [WEIGHT_SIZE-1:0] Wgt_8_601,input [WEIGHT_SIZE-1:0] Wgt_8_602,input [WEIGHT_SIZE-1:0] Wgt_8_603,input [WEIGHT_SIZE-1:0] Wgt_8_604,input [WEIGHT_SIZE-1:0] Wgt_8_605,input [WEIGHT_SIZE-1:0] Wgt_8_606,input [WEIGHT_SIZE-1:0] Wgt_8_607,input [WEIGHT_SIZE-1:0] Wgt_8_608,input [WEIGHT_SIZE-1:0] Wgt_8_609,input [WEIGHT_SIZE-1:0] Wgt_8_610,input [WEIGHT_SIZE-1:0] Wgt_8_611,input [WEIGHT_SIZE-1:0] Wgt_8_612,input [WEIGHT_SIZE-1:0] Wgt_8_613,input [WEIGHT_SIZE-1:0] Wgt_8_614,input [WEIGHT_SIZE-1:0] Wgt_8_615,input [WEIGHT_SIZE-1:0] Wgt_8_616,input [WEIGHT_SIZE-1:0] Wgt_8_617,input [WEIGHT_SIZE-1:0] Wgt_8_618,input [WEIGHT_SIZE-1:0] Wgt_8_619,input [WEIGHT_SIZE-1:0] Wgt_8_620,input [WEIGHT_SIZE-1:0] Wgt_8_621,input [WEIGHT_SIZE-1:0] Wgt_8_622,input [WEIGHT_SIZE-1:0] Wgt_8_623,input [WEIGHT_SIZE-1:0] Wgt_8_624,input [WEIGHT_SIZE-1:0] Wgt_8_625,input [WEIGHT_SIZE-1:0] Wgt_8_626,input [WEIGHT_SIZE-1:0] Wgt_8_627,input [WEIGHT_SIZE-1:0] Wgt_8_628,input [WEIGHT_SIZE-1:0] Wgt_8_629,input [WEIGHT_SIZE-1:0] Wgt_8_630,input [WEIGHT_SIZE-1:0] Wgt_8_631,input [WEIGHT_SIZE-1:0] Wgt_8_632,input [WEIGHT_SIZE-1:0] Wgt_8_633,input [WEIGHT_SIZE-1:0] Wgt_8_634,input [WEIGHT_SIZE-1:0] Wgt_8_635,input [WEIGHT_SIZE-1:0] Wgt_8_636,input [WEIGHT_SIZE-1:0] Wgt_8_637,input [WEIGHT_SIZE-1:0] Wgt_8_638,input [WEIGHT_SIZE-1:0] Wgt_8_639,input [WEIGHT_SIZE-1:0] Wgt_8_640,input [WEIGHT_SIZE-1:0] Wgt_8_641,input [WEIGHT_SIZE-1:0] Wgt_8_642,input [WEIGHT_SIZE-1:0] Wgt_8_643,input [WEIGHT_SIZE-1:0] Wgt_8_644,input [WEIGHT_SIZE-1:0] Wgt_8_645,input [WEIGHT_SIZE-1:0] Wgt_8_646,input [WEIGHT_SIZE-1:0] Wgt_8_647,input [WEIGHT_SIZE-1:0] Wgt_8_648,input [WEIGHT_SIZE-1:0] Wgt_8_649,input [WEIGHT_SIZE-1:0] Wgt_8_650,input [WEIGHT_SIZE-1:0] Wgt_8_651,input [WEIGHT_SIZE-1:0] Wgt_8_652,input [WEIGHT_SIZE-1:0] Wgt_8_653,input [WEIGHT_SIZE-1:0] Wgt_8_654,input [WEIGHT_SIZE-1:0] Wgt_8_655,input [WEIGHT_SIZE-1:0] Wgt_8_656,input [WEIGHT_SIZE-1:0] Wgt_8_657,input [WEIGHT_SIZE-1:0] Wgt_8_658,input [WEIGHT_SIZE-1:0] Wgt_8_659,input [WEIGHT_SIZE-1:0] Wgt_8_660,input [WEIGHT_SIZE-1:0] Wgt_8_661,input [WEIGHT_SIZE-1:0] Wgt_8_662,input [WEIGHT_SIZE-1:0] Wgt_8_663,input [WEIGHT_SIZE-1:0] Wgt_8_664,input [WEIGHT_SIZE-1:0] Wgt_8_665,input [WEIGHT_SIZE-1:0] Wgt_8_666,input [WEIGHT_SIZE-1:0] Wgt_8_667,input [WEIGHT_SIZE-1:0] Wgt_8_668,input [WEIGHT_SIZE-1:0] Wgt_8_669,input [WEIGHT_SIZE-1:0] Wgt_8_670,input [WEIGHT_SIZE-1:0] Wgt_8_671,input [WEIGHT_SIZE-1:0] Wgt_8_672,input [WEIGHT_SIZE-1:0] Wgt_8_673,input [WEIGHT_SIZE-1:0] Wgt_8_674,input [WEIGHT_SIZE-1:0] Wgt_8_675,input [WEIGHT_SIZE-1:0] Wgt_8_676,input [WEIGHT_SIZE-1:0] Wgt_8_677,input [WEIGHT_SIZE-1:0] Wgt_8_678,input [WEIGHT_SIZE-1:0] Wgt_8_679,input [WEIGHT_SIZE-1:0] Wgt_8_680,input [WEIGHT_SIZE-1:0] Wgt_8_681,input [WEIGHT_SIZE-1:0] Wgt_8_682,input [WEIGHT_SIZE-1:0] Wgt_8_683,input [WEIGHT_SIZE-1:0] Wgt_8_684,input [WEIGHT_SIZE-1:0] Wgt_8_685,input [WEIGHT_SIZE-1:0] Wgt_8_686,input [WEIGHT_SIZE-1:0] Wgt_8_687,input [WEIGHT_SIZE-1:0] Wgt_8_688,input [WEIGHT_SIZE-1:0] Wgt_8_689,input [WEIGHT_SIZE-1:0] Wgt_8_690,input [WEIGHT_SIZE-1:0] Wgt_8_691,input [WEIGHT_SIZE-1:0] Wgt_8_692,input [WEIGHT_SIZE-1:0] Wgt_8_693,input [WEIGHT_SIZE-1:0] Wgt_8_694,input [WEIGHT_SIZE-1:0] Wgt_8_695,input [WEIGHT_SIZE-1:0] Wgt_8_696,input [WEIGHT_SIZE-1:0] Wgt_8_697,input [WEIGHT_SIZE-1:0] Wgt_8_698,input [WEIGHT_SIZE-1:0] Wgt_8_699,input [WEIGHT_SIZE-1:0] Wgt_8_700,input [WEIGHT_SIZE-1:0] Wgt_8_701,input [WEIGHT_SIZE-1:0] Wgt_8_702,input [WEIGHT_SIZE-1:0] Wgt_8_703,input [WEIGHT_SIZE-1:0] Wgt_8_704,input [WEIGHT_SIZE-1:0] Wgt_8_705,input [WEIGHT_SIZE-1:0] Wgt_8_706,input [WEIGHT_SIZE-1:0] Wgt_8_707,input [WEIGHT_SIZE-1:0] Wgt_8_708,input [WEIGHT_SIZE-1:0] Wgt_8_709,input [WEIGHT_SIZE-1:0] Wgt_8_710,input [WEIGHT_SIZE-1:0] Wgt_8_711,input [WEIGHT_SIZE-1:0] Wgt_8_712,input [WEIGHT_SIZE-1:0] Wgt_8_713,input [WEIGHT_SIZE-1:0] Wgt_8_714,input [WEIGHT_SIZE-1:0] Wgt_8_715,input [WEIGHT_SIZE-1:0] Wgt_8_716,input [WEIGHT_SIZE-1:0] Wgt_8_717,input [WEIGHT_SIZE-1:0] Wgt_8_718,input [WEIGHT_SIZE-1:0] Wgt_8_719,input [WEIGHT_SIZE-1:0] Wgt_8_720,input [WEIGHT_SIZE-1:0] Wgt_8_721,input [WEIGHT_SIZE-1:0] Wgt_8_722,input [WEIGHT_SIZE-1:0] Wgt_8_723,input [WEIGHT_SIZE-1:0] Wgt_8_724,input [WEIGHT_SIZE-1:0] Wgt_8_725,input [WEIGHT_SIZE-1:0] Wgt_8_726,input [WEIGHT_SIZE-1:0] Wgt_8_727,input [WEIGHT_SIZE-1:0] Wgt_8_728,input [WEIGHT_SIZE-1:0] Wgt_8_729,input [WEIGHT_SIZE-1:0] Wgt_8_730,input [WEIGHT_SIZE-1:0] Wgt_8_731,input [WEIGHT_SIZE-1:0] Wgt_8_732,input [WEIGHT_SIZE-1:0] Wgt_8_733,input [WEIGHT_SIZE-1:0] Wgt_8_734,input [WEIGHT_SIZE-1:0] Wgt_8_735,input [WEIGHT_SIZE-1:0] Wgt_8_736,input [WEIGHT_SIZE-1:0] Wgt_8_737,input [WEIGHT_SIZE-1:0] Wgt_8_738,input [WEIGHT_SIZE-1:0] Wgt_8_739,input [WEIGHT_SIZE-1:0] Wgt_8_740,input [WEIGHT_SIZE-1:0] Wgt_8_741,input [WEIGHT_SIZE-1:0] Wgt_8_742,input [WEIGHT_SIZE-1:0] Wgt_8_743,input [WEIGHT_SIZE-1:0] Wgt_8_744,input [WEIGHT_SIZE-1:0] Wgt_8_745,input [WEIGHT_SIZE-1:0] Wgt_8_746,input [WEIGHT_SIZE-1:0] Wgt_8_747,input [WEIGHT_SIZE-1:0] Wgt_8_748,input [WEIGHT_SIZE-1:0] Wgt_8_749,input [WEIGHT_SIZE-1:0] Wgt_8_750,input [WEIGHT_SIZE-1:0] Wgt_8_751,input [WEIGHT_SIZE-1:0] Wgt_8_752,input [WEIGHT_SIZE-1:0] Wgt_8_753,input [WEIGHT_SIZE-1:0] Wgt_8_754,input [WEIGHT_SIZE-1:0] Wgt_8_755,input [WEIGHT_SIZE-1:0] Wgt_8_756,input [WEIGHT_SIZE-1:0] Wgt_8_757,input [WEIGHT_SIZE-1:0] Wgt_8_758,input [WEIGHT_SIZE-1:0] Wgt_8_759,input [WEIGHT_SIZE-1:0] Wgt_8_760,input [WEIGHT_SIZE-1:0] Wgt_8_761,input [WEIGHT_SIZE-1:0] Wgt_8_762,input [WEIGHT_SIZE-1:0] Wgt_8_763,input [WEIGHT_SIZE-1:0] Wgt_8_764,input [WEIGHT_SIZE-1:0] Wgt_8_765,input [WEIGHT_SIZE-1:0] Wgt_8_766,input [WEIGHT_SIZE-1:0] Wgt_8_767,input [WEIGHT_SIZE-1:0] Wgt_8_768,input [WEIGHT_SIZE-1:0] Wgt_8_769,input [WEIGHT_SIZE-1:0] Wgt_8_770,input [WEIGHT_SIZE-1:0] Wgt_8_771,input [WEIGHT_SIZE-1:0] Wgt_8_772,input [WEIGHT_SIZE-1:0] Wgt_8_773,input [WEIGHT_SIZE-1:0] Wgt_8_774,input [WEIGHT_SIZE-1:0] Wgt_8_775,input [WEIGHT_SIZE-1:0] Wgt_8_776,input [WEIGHT_SIZE-1:0] Wgt_8_777,input [WEIGHT_SIZE-1:0] Wgt_8_778,input [WEIGHT_SIZE-1:0] Wgt_8_779,input [WEIGHT_SIZE-1:0] Wgt_8_780,input [WEIGHT_SIZE-1:0] Wgt_8_781,input [WEIGHT_SIZE-1:0] Wgt_8_782,input [WEIGHT_SIZE-1:0] Wgt_8_783,input [WEIGHT_SIZE-1:0] Wgt_8_784,input [WEIGHT_SIZE-1:0] Wgt_9_0,input [WEIGHT_SIZE-1:0] Wgt_9_1,input [WEIGHT_SIZE-1:0] Wgt_9_2,input [WEIGHT_SIZE-1:0] Wgt_9_3,input [WEIGHT_SIZE-1:0] Wgt_9_4,input [WEIGHT_SIZE-1:0] Wgt_9_5,input [WEIGHT_SIZE-1:0] Wgt_9_6,input [WEIGHT_SIZE-1:0] Wgt_9_7,input [WEIGHT_SIZE-1:0] Wgt_9_8,input [WEIGHT_SIZE-1:0] Wgt_9_9,input [WEIGHT_SIZE-1:0] Wgt_9_10,input [WEIGHT_SIZE-1:0] Wgt_9_11,input [WEIGHT_SIZE-1:0] Wgt_9_12,input [WEIGHT_SIZE-1:0] Wgt_9_13,input [WEIGHT_SIZE-1:0] Wgt_9_14,input [WEIGHT_SIZE-1:0] Wgt_9_15,input [WEIGHT_SIZE-1:0] Wgt_9_16,input [WEIGHT_SIZE-1:0] Wgt_9_17,input [WEIGHT_SIZE-1:0] Wgt_9_18,input [WEIGHT_SIZE-1:0] Wgt_9_19,input [WEIGHT_SIZE-1:0] Wgt_9_20,input [WEIGHT_SIZE-1:0] Wgt_9_21,input [WEIGHT_SIZE-1:0] Wgt_9_22,input [WEIGHT_SIZE-1:0] Wgt_9_23,input [WEIGHT_SIZE-1:0] Wgt_9_24,input [WEIGHT_SIZE-1:0] Wgt_9_25,input [WEIGHT_SIZE-1:0] Wgt_9_26,input [WEIGHT_SIZE-1:0] Wgt_9_27,input [WEIGHT_SIZE-1:0] Wgt_9_28,input [WEIGHT_SIZE-1:0] Wgt_9_29,input [WEIGHT_SIZE-1:0] Wgt_9_30,input [WEIGHT_SIZE-1:0] Wgt_9_31,input [WEIGHT_SIZE-1:0] Wgt_9_32,input [WEIGHT_SIZE-1:0] Wgt_9_33,input [WEIGHT_SIZE-1:0] Wgt_9_34,input [WEIGHT_SIZE-1:0] Wgt_9_35,input [WEIGHT_SIZE-1:0] Wgt_9_36,input [WEIGHT_SIZE-1:0] Wgt_9_37,input [WEIGHT_SIZE-1:0] Wgt_9_38,input [WEIGHT_SIZE-1:0] Wgt_9_39,input [WEIGHT_SIZE-1:0] Wgt_9_40,input [WEIGHT_SIZE-1:0] Wgt_9_41,input [WEIGHT_SIZE-1:0] Wgt_9_42,input [WEIGHT_SIZE-1:0] Wgt_9_43,input [WEIGHT_SIZE-1:0] Wgt_9_44,input [WEIGHT_SIZE-1:0] Wgt_9_45,input [WEIGHT_SIZE-1:0] Wgt_9_46,input [WEIGHT_SIZE-1:0] Wgt_9_47,input [WEIGHT_SIZE-1:0] Wgt_9_48,input [WEIGHT_SIZE-1:0] Wgt_9_49,input [WEIGHT_SIZE-1:0] Wgt_9_50,input [WEIGHT_SIZE-1:0] Wgt_9_51,input [WEIGHT_SIZE-1:0] Wgt_9_52,input [WEIGHT_SIZE-1:0] Wgt_9_53,input [WEIGHT_SIZE-1:0] Wgt_9_54,input [WEIGHT_SIZE-1:0] Wgt_9_55,input [WEIGHT_SIZE-1:0] Wgt_9_56,input [WEIGHT_SIZE-1:0] Wgt_9_57,input [WEIGHT_SIZE-1:0] Wgt_9_58,input [WEIGHT_SIZE-1:0] Wgt_9_59,input [WEIGHT_SIZE-1:0] Wgt_9_60,input [WEIGHT_SIZE-1:0] Wgt_9_61,input [WEIGHT_SIZE-1:0] Wgt_9_62,input [WEIGHT_SIZE-1:0] Wgt_9_63,input [WEIGHT_SIZE-1:0] Wgt_9_64,input [WEIGHT_SIZE-1:0] Wgt_9_65,input [WEIGHT_SIZE-1:0] Wgt_9_66,input [WEIGHT_SIZE-1:0] Wgt_9_67,input [WEIGHT_SIZE-1:0] Wgt_9_68,input [WEIGHT_SIZE-1:0] Wgt_9_69,input [WEIGHT_SIZE-1:0] Wgt_9_70,input [WEIGHT_SIZE-1:0] Wgt_9_71,input [WEIGHT_SIZE-1:0] Wgt_9_72,input [WEIGHT_SIZE-1:0] Wgt_9_73,input [WEIGHT_SIZE-1:0] Wgt_9_74,input [WEIGHT_SIZE-1:0] Wgt_9_75,input [WEIGHT_SIZE-1:0] Wgt_9_76,input [WEIGHT_SIZE-1:0] Wgt_9_77,input [WEIGHT_SIZE-1:0] Wgt_9_78,input [WEIGHT_SIZE-1:0] Wgt_9_79,input [WEIGHT_SIZE-1:0] Wgt_9_80,input [WEIGHT_SIZE-1:0] Wgt_9_81,input [WEIGHT_SIZE-1:0] Wgt_9_82,input [WEIGHT_SIZE-1:0] Wgt_9_83,input [WEIGHT_SIZE-1:0] Wgt_9_84,input [WEIGHT_SIZE-1:0] Wgt_9_85,input [WEIGHT_SIZE-1:0] Wgt_9_86,input [WEIGHT_SIZE-1:0] Wgt_9_87,input [WEIGHT_SIZE-1:0] Wgt_9_88,input [WEIGHT_SIZE-1:0] Wgt_9_89,input [WEIGHT_SIZE-1:0] Wgt_9_90,input [WEIGHT_SIZE-1:0] Wgt_9_91,input [WEIGHT_SIZE-1:0] Wgt_9_92,input [WEIGHT_SIZE-1:0] Wgt_9_93,input [WEIGHT_SIZE-1:0] Wgt_9_94,input [WEIGHT_SIZE-1:0] Wgt_9_95,input [WEIGHT_SIZE-1:0] Wgt_9_96,input [WEIGHT_SIZE-1:0] Wgt_9_97,input [WEIGHT_SIZE-1:0] Wgt_9_98,input [WEIGHT_SIZE-1:0] Wgt_9_99,input [WEIGHT_SIZE-1:0] Wgt_9_100,input [WEIGHT_SIZE-1:0] Wgt_9_101,input [WEIGHT_SIZE-1:0] Wgt_9_102,input [WEIGHT_SIZE-1:0] Wgt_9_103,input [WEIGHT_SIZE-1:0] Wgt_9_104,input [WEIGHT_SIZE-1:0] Wgt_9_105,input [WEIGHT_SIZE-1:0] Wgt_9_106,input [WEIGHT_SIZE-1:0] Wgt_9_107,input [WEIGHT_SIZE-1:0] Wgt_9_108,input [WEIGHT_SIZE-1:0] Wgt_9_109,input [WEIGHT_SIZE-1:0] Wgt_9_110,input [WEIGHT_SIZE-1:0] Wgt_9_111,input [WEIGHT_SIZE-1:0] Wgt_9_112,input [WEIGHT_SIZE-1:0] Wgt_9_113,input [WEIGHT_SIZE-1:0] Wgt_9_114,input [WEIGHT_SIZE-1:0] Wgt_9_115,input [WEIGHT_SIZE-1:0] Wgt_9_116,input [WEIGHT_SIZE-1:0] Wgt_9_117,input [WEIGHT_SIZE-1:0] Wgt_9_118,input [WEIGHT_SIZE-1:0] Wgt_9_119,input [WEIGHT_SIZE-1:0] Wgt_9_120,input [WEIGHT_SIZE-1:0] Wgt_9_121,input [WEIGHT_SIZE-1:0] Wgt_9_122,input [WEIGHT_SIZE-1:0] Wgt_9_123,input [WEIGHT_SIZE-1:0] Wgt_9_124,input [WEIGHT_SIZE-1:0] Wgt_9_125,input [WEIGHT_SIZE-1:0] Wgt_9_126,input [WEIGHT_SIZE-1:0] Wgt_9_127,input [WEIGHT_SIZE-1:0] Wgt_9_128,input [WEIGHT_SIZE-1:0] Wgt_9_129,input [WEIGHT_SIZE-1:0] Wgt_9_130,input [WEIGHT_SIZE-1:0] Wgt_9_131,input [WEIGHT_SIZE-1:0] Wgt_9_132,input [WEIGHT_SIZE-1:0] Wgt_9_133,input [WEIGHT_SIZE-1:0] Wgt_9_134,input [WEIGHT_SIZE-1:0] Wgt_9_135,input [WEIGHT_SIZE-1:0] Wgt_9_136,input [WEIGHT_SIZE-1:0] Wgt_9_137,input [WEIGHT_SIZE-1:0] Wgt_9_138,input [WEIGHT_SIZE-1:0] Wgt_9_139,input [WEIGHT_SIZE-1:0] Wgt_9_140,input [WEIGHT_SIZE-1:0] Wgt_9_141,input [WEIGHT_SIZE-1:0] Wgt_9_142,input [WEIGHT_SIZE-1:0] Wgt_9_143,input [WEIGHT_SIZE-1:0] Wgt_9_144,input [WEIGHT_SIZE-1:0] Wgt_9_145,input [WEIGHT_SIZE-1:0] Wgt_9_146,input [WEIGHT_SIZE-1:0] Wgt_9_147,input [WEIGHT_SIZE-1:0] Wgt_9_148,input [WEIGHT_SIZE-1:0] Wgt_9_149,input [WEIGHT_SIZE-1:0] Wgt_9_150,input [WEIGHT_SIZE-1:0] Wgt_9_151,input [WEIGHT_SIZE-1:0] Wgt_9_152,input [WEIGHT_SIZE-1:0] Wgt_9_153,input [WEIGHT_SIZE-1:0] Wgt_9_154,input [WEIGHT_SIZE-1:0] Wgt_9_155,input [WEIGHT_SIZE-1:0] Wgt_9_156,input [WEIGHT_SIZE-1:0] Wgt_9_157,input [WEIGHT_SIZE-1:0] Wgt_9_158,input [WEIGHT_SIZE-1:0] Wgt_9_159,input [WEIGHT_SIZE-1:0] Wgt_9_160,input [WEIGHT_SIZE-1:0] Wgt_9_161,input [WEIGHT_SIZE-1:0] Wgt_9_162,input [WEIGHT_SIZE-1:0] Wgt_9_163,input [WEIGHT_SIZE-1:0] Wgt_9_164,input [WEIGHT_SIZE-1:0] Wgt_9_165,input [WEIGHT_SIZE-1:0] Wgt_9_166,input [WEIGHT_SIZE-1:0] Wgt_9_167,input [WEIGHT_SIZE-1:0] Wgt_9_168,input [WEIGHT_SIZE-1:0] Wgt_9_169,input [WEIGHT_SIZE-1:0] Wgt_9_170,input [WEIGHT_SIZE-1:0] Wgt_9_171,input [WEIGHT_SIZE-1:0] Wgt_9_172,input [WEIGHT_SIZE-1:0] Wgt_9_173,input [WEIGHT_SIZE-1:0] Wgt_9_174,input [WEIGHT_SIZE-1:0] Wgt_9_175,input [WEIGHT_SIZE-1:0] Wgt_9_176,input [WEIGHT_SIZE-1:0] Wgt_9_177,input [WEIGHT_SIZE-1:0] Wgt_9_178,input [WEIGHT_SIZE-1:0] Wgt_9_179,input [WEIGHT_SIZE-1:0] Wgt_9_180,input [WEIGHT_SIZE-1:0] Wgt_9_181,input [WEIGHT_SIZE-1:0] Wgt_9_182,input [WEIGHT_SIZE-1:0] Wgt_9_183,input [WEIGHT_SIZE-1:0] Wgt_9_184,input [WEIGHT_SIZE-1:0] Wgt_9_185,input [WEIGHT_SIZE-1:0] Wgt_9_186,input [WEIGHT_SIZE-1:0] Wgt_9_187,input [WEIGHT_SIZE-1:0] Wgt_9_188,input [WEIGHT_SIZE-1:0] Wgt_9_189,input [WEIGHT_SIZE-1:0] Wgt_9_190,input [WEIGHT_SIZE-1:0] Wgt_9_191,input [WEIGHT_SIZE-1:0] Wgt_9_192,input [WEIGHT_SIZE-1:0] Wgt_9_193,input [WEIGHT_SIZE-1:0] Wgt_9_194,input [WEIGHT_SIZE-1:0] Wgt_9_195,input [WEIGHT_SIZE-1:0] Wgt_9_196,input [WEIGHT_SIZE-1:0] Wgt_9_197,input [WEIGHT_SIZE-1:0] Wgt_9_198,input [WEIGHT_SIZE-1:0] Wgt_9_199,input [WEIGHT_SIZE-1:0] Wgt_9_200,input [WEIGHT_SIZE-1:0] Wgt_9_201,input [WEIGHT_SIZE-1:0] Wgt_9_202,input [WEIGHT_SIZE-1:0] Wgt_9_203,input [WEIGHT_SIZE-1:0] Wgt_9_204,input [WEIGHT_SIZE-1:0] Wgt_9_205,input [WEIGHT_SIZE-1:0] Wgt_9_206,input [WEIGHT_SIZE-1:0] Wgt_9_207,input [WEIGHT_SIZE-1:0] Wgt_9_208,input [WEIGHT_SIZE-1:0] Wgt_9_209,input [WEIGHT_SIZE-1:0] Wgt_9_210,input [WEIGHT_SIZE-1:0] Wgt_9_211,input [WEIGHT_SIZE-1:0] Wgt_9_212,input [WEIGHT_SIZE-1:0] Wgt_9_213,input [WEIGHT_SIZE-1:0] Wgt_9_214,input [WEIGHT_SIZE-1:0] Wgt_9_215,input [WEIGHT_SIZE-1:0] Wgt_9_216,input [WEIGHT_SIZE-1:0] Wgt_9_217,input [WEIGHT_SIZE-1:0] Wgt_9_218,input [WEIGHT_SIZE-1:0] Wgt_9_219,input [WEIGHT_SIZE-1:0] Wgt_9_220,input [WEIGHT_SIZE-1:0] Wgt_9_221,input [WEIGHT_SIZE-1:0] Wgt_9_222,input [WEIGHT_SIZE-1:0] Wgt_9_223,input [WEIGHT_SIZE-1:0] Wgt_9_224,input [WEIGHT_SIZE-1:0] Wgt_9_225,input [WEIGHT_SIZE-1:0] Wgt_9_226,input [WEIGHT_SIZE-1:0] Wgt_9_227,input [WEIGHT_SIZE-1:0] Wgt_9_228,input [WEIGHT_SIZE-1:0] Wgt_9_229,input [WEIGHT_SIZE-1:0] Wgt_9_230,input [WEIGHT_SIZE-1:0] Wgt_9_231,input [WEIGHT_SIZE-1:0] Wgt_9_232,input [WEIGHT_SIZE-1:0] Wgt_9_233,input [WEIGHT_SIZE-1:0] Wgt_9_234,input [WEIGHT_SIZE-1:0] Wgt_9_235,input [WEIGHT_SIZE-1:0] Wgt_9_236,input [WEIGHT_SIZE-1:0] Wgt_9_237,input [WEIGHT_SIZE-1:0] Wgt_9_238,input [WEIGHT_SIZE-1:0] Wgt_9_239,input [WEIGHT_SIZE-1:0] Wgt_9_240,input [WEIGHT_SIZE-1:0] Wgt_9_241,input [WEIGHT_SIZE-1:0] Wgt_9_242,input [WEIGHT_SIZE-1:0] Wgt_9_243,input [WEIGHT_SIZE-1:0] Wgt_9_244,input [WEIGHT_SIZE-1:0] Wgt_9_245,input [WEIGHT_SIZE-1:0] Wgt_9_246,input [WEIGHT_SIZE-1:0] Wgt_9_247,input [WEIGHT_SIZE-1:0] Wgt_9_248,input [WEIGHT_SIZE-1:0] Wgt_9_249,input [WEIGHT_SIZE-1:0] Wgt_9_250,input [WEIGHT_SIZE-1:0] Wgt_9_251,input [WEIGHT_SIZE-1:0] Wgt_9_252,input [WEIGHT_SIZE-1:0] Wgt_9_253,input [WEIGHT_SIZE-1:0] Wgt_9_254,input [WEIGHT_SIZE-1:0] Wgt_9_255,input [WEIGHT_SIZE-1:0] Wgt_9_256,input [WEIGHT_SIZE-1:0] Wgt_9_257,input [WEIGHT_SIZE-1:0] Wgt_9_258,input [WEIGHT_SIZE-1:0] Wgt_9_259,input [WEIGHT_SIZE-1:0] Wgt_9_260,input [WEIGHT_SIZE-1:0] Wgt_9_261,input [WEIGHT_SIZE-1:0] Wgt_9_262,input [WEIGHT_SIZE-1:0] Wgt_9_263,input [WEIGHT_SIZE-1:0] Wgt_9_264,input [WEIGHT_SIZE-1:0] Wgt_9_265,input [WEIGHT_SIZE-1:0] Wgt_9_266,input [WEIGHT_SIZE-1:0] Wgt_9_267,input [WEIGHT_SIZE-1:0] Wgt_9_268,input [WEIGHT_SIZE-1:0] Wgt_9_269,input [WEIGHT_SIZE-1:0] Wgt_9_270,input [WEIGHT_SIZE-1:0] Wgt_9_271,input [WEIGHT_SIZE-1:0] Wgt_9_272,input [WEIGHT_SIZE-1:0] Wgt_9_273,input [WEIGHT_SIZE-1:0] Wgt_9_274,input [WEIGHT_SIZE-1:0] Wgt_9_275,input [WEIGHT_SIZE-1:0] Wgt_9_276,input [WEIGHT_SIZE-1:0] Wgt_9_277,input [WEIGHT_SIZE-1:0] Wgt_9_278,input [WEIGHT_SIZE-1:0] Wgt_9_279,input [WEIGHT_SIZE-1:0] Wgt_9_280,input [WEIGHT_SIZE-1:0] Wgt_9_281,input [WEIGHT_SIZE-1:0] Wgt_9_282,input [WEIGHT_SIZE-1:0] Wgt_9_283,input [WEIGHT_SIZE-1:0] Wgt_9_284,input [WEIGHT_SIZE-1:0] Wgt_9_285,input [WEIGHT_SIZE-1:0] Wgt_9_286,input [WEIGHT_SIZE-1:0] Wgt_9_287,input [WEIGHT_SIZE-1:0] Wgt_9_288,input [WEIGHT_SIZE-1:0] Wgt_9_289,input [WEIGHT_SIZE-1:0] Wgt_9_290,input [WEIGHT_SIZE-1:0] Wgt_9_291,input [WEIGHT_SIZE-1:0] Wgt_9_292,input [WEIGHT_SIZE-1:0] Wgt_9_293,input [WEIGHT_SIZE-1:0] Wgt_9_294,input [WEIGHT_SIZE-1:0] Wgt_9_295,input [WEIGHT_SIZE-1:0] Wgt_9_296,input [WEIGHT_SIZE-1:0] Wgt_9_297,input [WEIGHT_SIZE-1:0] Wgt_9_298,input [WEIGHT_SIZE-1:0] Wgt_9_299,input [WEIGHT_SIZE-1:0] Wgt_9_300,input [WEIGHT_SIZE-1:0] Wgt_9_301,input [WEIGHT_SIZE-1:0] Wgt_9_302,input [WEIGHT_SIZE-1:0] Wgt_9_303,input [WEIGHT_SIZE-1:0] Wgt_9_304,input [WEIGHT_SIZE-1:0] Wgt_9_305,input [WEIGHT_SIZE-1:0] Wgt_9_306,input [WEIGHT_SIZE-1:0] Wgt_9_307,input [WEIGHT_SIZE-1:0] Wgt_9_308,input [WEIGHT_SIZE-1:0] Wgt_9_309,input [WEIGHT_SIZE-1:0] Wgt_9_310,input [WEIGHT_SIZE-1:0] Wgt_9_311,input [WEIGHT_SIZE-1:0] Wgt_9_312,input [WEIGHT_SIZE-1:0] Wgt_9_313,input [WEIGHT_SIZE-1:0] Wgt_9_314,input [WEIGHT_SIZE-1:0] Wgt_9_315,input [WEIGHT_SIZE-1:0] Wgt_9_316,input [WEIGHT_SIZE-1:0] Wgt_9_317,input [WEIGHT_SIZE-1:0] Wgt_9_318,input [WEIGHT_SIZE-1:0] Wgt_9_319,input [WEIGHT_SIZE-1:0] Wgt_9_320,input [WEIGHT_SIZE-1:0] Wgt_9_321,input [WEIGHT_SIZE-1:0] Wgt_9_322,input [WEIGHT_SIZE-1:0] Wgt_9_323,input [WEIGHT_SIZE-1:0] Wgt_9_324,input [WEIGHT_SIZE-1:0] Wgt_9_325,input [WEIGHT_SIZE-1:0] Wgt_9_326,input [WEIGHT_SIZE-1:0] Wgt_9_327,input [WEIGHT_SIZE-1:0] Wgt_9_328,input [WEIGHT_SIZE-1:0] Wgt_9_329,input [WEIGHT_SIZE-1:0] Wgt_9_330,input [WEIGHT_SIZE-1:0] Wgt_9_331,input [WEIGHT_SIZE-1:0] Wgt_9_332,input [WEIGHT_SIZE-1:0] Wgt_9_333,input [WEIGHT_SIZE-1:0] Wgt_9_334,input [WEIGHT_SIZE-1:0] Wgt_9_335,input [WEIGHT_SIZE-1:0] Wgt_9_336,input [WEIGHT_SIZE-1:0] Wgt_9_337,input [WEIGHT_SIZE-1:0] Wgt_9_338,input [WEIGHT_SIZE-1:0] Wgt_9_339,input [WEIGHT_SIZE-1:0] Wgt_9_340,input [WEIGHT_SIZE-1:0] Wgt_9_341,input [WEIGHT_SIZE-1:0] Wgt_9_342,input [WEIGHT_SIZE-1:0] Wgt_9_343,input [WEIGHT_SIZE-1:0] Wgt_9_344,input [WEIGHT_SIZE-1:0] Wgt_9_345,input [WEIGHT_SIZE-1:0] Wgt_9_346,input [WEIGHT_SIZE-1:0] Wgt_9_347,input [WEIGHT_SIZE-1:0] Wgt_9_348,input [WEIGHT_SIZE-1:0] Wgt_9_349,input [WEIGHT_SIZE-1:0] Wgt_9_350,input [WEIGHT_SIZE-1:0] Wgt_9_351,input [WEIGHT_SIZE-1:0] Wgt_9_352,input [WEIGHT_SIZE-1:0] Wgt_9_353,input [WEIGHT_SIZE-1:0] Wgt_9_354,input [WEIGHT_SIZE-1:0] Wgt_9_355,input [WEIGHT_SIZE-1:0] Wgt_9_356,input [WEIGHT_SIZE-1:0] Wgt_9_357,input [WEIGHT_SIZE-1:0] Wgt_9_358,input [WEIGHT_SIZE-1:0] Wgt_9_359,input [WEIGHT_SIZE-1:0] Wgt_9_360,input [WEIGHT_SIZE-1:0] Wgt_9_361,input [WEIGHT_SIZE-1:0] Wgt_9_362,input [WEIGHT_SIZE-1:0] Wgt_9_363,input [WEIGHT_SIZE-1:0] Wgt_9_364,input [WEIGHT_SIZE-1:0] Wgt_9_365,input [WEIGHT_SIZE-1:0] Wgt_9_366,input [WEIGHT_SIZE-1:0] Wgt_9_367,input [WEIGHT_SIZE-1:0] Wgt_9_368,input [WEIGHT_SIZE-1:0] Wgt_9_369,input [WEIGHT_SIZE-1:0] Wgt_9_370,input [WEIGHT_SIZE-1:0] Wgt_9_371,input [WEIGHT_SIZE-1:0] Wgt_9_372,input [WEIGHT_SIZE-1:0] Wgt_9_373,input [WEIGHT_SIZE-1:0] Wgt_9_374,input [WEIGHT_SIZE-1:0] Wgt_9_375,input [WEIGHT_SIZE-1:0] Wgt_9_376,input [WEIGHT_SIZE-1:0] Wgt_9_377,input [WEIGHT_SIZE-1:0] Wgt_9_378,input [WEIGHT_SIZE-1:0] Wgt_9_379,input [WEIGHT_SIZE-1:0] Wgt_9_380,input [WEIGHT_SIZE-1:0] Wgt_9_381,input [WEIGHT_SIZE-1:0] Wgt_9_382,input [WEIGHT_SIZE-1:0] Wgt_9_383,input [WEIGHT_SIZE-1:0] Wgt_9_384,input [WEIGHT_SIZE-1:0] Wgt_9_385,input [WEIGHT_SIZE-1:0] Wgt_9_386,input [WEIGHT_SIZE-1:0] Wgt_9_387,input [WEIGHT_SIZE-1:0] Wgt_9_388,input [WEIGHT_SIZE-1:0] Wgt_9_389,input [WEIGHT_SIZE-1:0] Wgt_9_390,input [WEIGHT_SIZE-1:0] Wgt_9_391,input [WEIGHT_SIZE-1:0] Wgt_9_392,input [WEIGHT_SIZE-1:0] Wgt_9_393,input [WEIGHT_SIZE-1:0] Wgt_9_394,input [WEIGHT_SIZE-1:0] Wgt_9_395,input [WEIGHT_SIZE-1:0] Wgt_9_396,input [WEIGHT_SIZE-1:0] Wgt_9_397,input [WEIGHT_SIZE-1:0] Wgt_9_398,input [WEIGHT_SIZE-1:0] Wgt_9_399,input [WEIGHT_SIZE-1:0] Wgt_9_400,input [WEIGHT_SIZE-1:0] Wgt_9_401,input [WEIGHT_SIZE-1:0] Wgt_9_402,input [WEIGHT_SIZE-1:0] Wgt_9_403,input [WEIGHT_SIZE-1:0] Wgt_9_404,input [WEIGHT_SIZE-1:0] Wgt_9_405,input [WEIGHT_SIZE-1:0] Wgt_9_406,input [WEIGHT_SIZE-1:0] Wgt_9_407,input [WEIGHT_SIZE-1:0] Wgt_9_408,input [WEIGHT_SIZE-1:0] Wgt_9_409,input [WEIGHT_SIZE-1:0] Wgt_9_410,input [WEIGHT_SIZE-1:0] Wgt_9_411,input [WEIGHT_SIZE-1:0] Wgt_9_412,input [WEIGHT_SIZE-1:0] Wgt_9_413,input [WEIGHT_SIZE-1:0] Wgt_9_414,input [WEIGHT_SIZE-1:0] Wgt_9_415,input [WEIGHT_SIZE-1:0] Wgt_9_416,input [WEIGHT_SIZE-1:0] Wgt_9_417,input [WEIGHT_SIZE-1:0] Wgt_9_418,input [WEIGHT_SIZE-1:0] Wgt_9_419,input [WEIGHT_SIZE-1:0] Wgt_9_420,input [WEIGHT_SIZE-1:0] Wgt_9_421,input [WEIGHT_SIZE-1:0] Wgt_9_422,input [WEIGHT_SIZE-1:0] Wgt_9_423,input [WEIGHT_SIZE-1:0] Wgt_9_424,input [WEIGHT_SIZE-1:0] Wgt_9_425,input [WEIGHT_SIZE-1:0] Wgt_9_426,input [WEIGHT_SIZE-1:0] Wgt_9_427,input [WEIGHT_SIZE-1:0] Wgt_9_428,input [WEIGHT_SIZE-1:0] Wgt_9_429,input [WEIGHT_SIZE-1:0] Wgt_9_430,input [WEIGHT_SIZE-1:0] Wgt_9_431,input [WEIGHT_SIZE-1:0] Wgt_9_432,input [WEIGHT_SIZE-1:0] Wgt_9_433,input [WEIGHT_SIZE-1:0] Wgt_9_434,input [WEIGHT_SIZE-1:0] Wgt_9_435,input [WEIGHT_SIZE-1:0] Wgt_9_436,input [WEIGHT_SIZE-1:0] Wgt_9_437,input [WEIGHT_SIZE-1:0] Wgt_9_438,input [WEIGHT_SIZE-1:0] Wgt_9_439,input [WEIGHT_SIZE-1:0] Wgt_9_440,input [WEIGHT_SIZE-1:0] Wgt_9_441,input [WEIGHT_SIZE-1:0] Wgt_9_442,input [WEIGHT_SIZE-1:0] Wgt_9_443,input [WEIGHT_SIZE-1:0] Wgt_9_444,input [WEIGHT_SIZE-1:0] Wgt_9_445,input [WEIGHT_SIZE-1:0] Wgt_9_446,input [WEIGHT_SIZE-1:0] Wgt_9_447,input [WEIGHT_SIZE-1:0] Wgt_9_448,input [WEIGHT_SIZE-1:0] Wgt_9_449,input [WEIGHT_SIZE-1:0] Wgt_9_450,input [WEIGHT_SIZE-1:0] Wgt_9_451,input [WEIGHT_SIZE-1:0] Wgt_9_452,input [WEIGHT_SIZE-1:0] Wgt_9_453,input [WEIGHT_SIZE-1:0] Wgt_9_454,input [WEIGHT_SIZE-1:0] Wgt_9_455,input [WEIGHT_SIZE-1:0] Wgt_9_456,input [WEIGHT_SIZE-1:0] Wgt_9_457,input [WEIGHT_SIZE-1:0] Wgt_9_458,input [WEIGHT_SIZE-1:0] Wgt_9_459,input [WEIGHT_SIZE-1:0] Wgt_9_460,input [WEIGHT_SIZE-1:0] Wgt_9_461,input [WEIGHT_SIZE-1:0] Wgt_9_462,input [WEIGHT_SIZE-1:0] Wgt_9_463,input [WEIGHT_SIZE-1:0] Wgt_9_464,input [WEIGHT_SIZE-1:0] Wgt_9_465,input [WEIGHT_SIZE-1:0] Wgt_9_466,input [WEIGHT_SIZE-1:0] Wgt_9_467,input [WEIGHT_SIZE-1:0] Wgt_9_468,input [WEIGHT_SIZE-1:0] Wgt_9_469,input [WEIGHT_SIZE-1:0] Wgt_9_470,input [WEIGHT_SIZE-1:0] Wgt_9_471,input [WEIGHT_SIZE-1:0] Wgt_9_472,input [WEIGHT_SIZE-1:0] Wgt_9_473,input [WEIGHT_SIZE-1:0] Wgt_9_474,input [WEIGHT_SIZE-1:0] Wgt_9_475,input [WEIGHT_SIZE-1:0] Wgt_9_476,input [WEIGHT_SIZE-1:0] Wgt_9_477,input [WEIGHT_SIZE-1:0] Wgt_9_478,input [WEIGHT_SIZE-1:0] Wgt_9_479,input [WEIGHT_SIZE-1:0] Wgt_9_480,input [WEIGHT_SIZE-1:0] Wgt_9_481,input [WEIGHT_SIZE-1:0] Wgt_9_482,input [WEIGHT_SIZE-1:0] Wgt_9_483,input [WEIGHT_SIZE-1:0] Wgt_9_484,input [WEIGHT_SIZE-1:0] Wgt_9_485,input [WEIGHT_SIZE-1:0] Wgt_9_486,input [WEIGHT_SIZE-1:0] Wgt_9_487,input [WEIGHT_SIZE-1:0] Wgt_9_488,input [WEIGHT_SIZE-1:0] Wgt_9_489,input [WEIGHT_SIZE-1:0] Wgt_9_490,input [WEIGHT_SIZE-1:0] Wgt_9_491,input [WEIGHT_SIZE-1:0] Wgt_9_492,input [WEIGHT_SIZE-1:0] Wgt_9_493,input [WEIGHT_SIZE-1:0] Wgt_9_494,input [WEIGHT_SIZE-1:0] Wgt_9_495,input [WEIGHT_SIZE-1:0] Wgt_9_496,input [WEIGHT_SIZE-1:0] Wgt_9_497,input [WEIGHT_SIZE-1:0] Wgt_9_498,input [WEIGHT_SIZE-1:0] Wgt_9_499,input [WEIGHT_SIZE-1:0] Wgt_9_500,input [WEIGHT_SIZE-1:0] Wgt_9_501,input [WEIGHT_SIZE-1:0] Wgt_9_502,input [WEIGHT_SIZE-1:0] Wgt_9_503,input [WEIGHT_SIZE-1:0] Wgt_9_504,input [WEIGHT_SIZE-1:0] Wgt_9_505,input [WEIGHT_SIZE-1:0] Wgt_9_506,input [WEIGHT_SIZE-1:0] Wgt_9_507,input [WEIGHT_SIZE-1:0] Wgt_9_508,input [WEIGHT_SIZE-1:0] Wgt_9_509,input [WEIGHT_SIZE-1:0] Wgt_9_510,input [WEIGHT_SIZE-1:0] Wgt_9_511,input [WEIGHT_SIZE-1:0] Wgt_9_512,input [WEIGHT_SIZE-1:0] Wgt_9_513,input [WEIGHT_SIZE-1:0] Wgt_9_514,input [WEIGHT_SIZE-1:0] Wgt_9_515,input [WEIGHT_SIZE-1:0] Wgt_9_516,input [WEIGHT_SIZE-1:0] Wgt_9_517,input [WEIGHT_SIZE-1:0] Wgt_9_518,input [WEIGHT_SIZE-1:0] Wgt_9_519,input [WEIGHT_SIZE-1:0] Wgt_9_520,input [WEIGHT_SIZE-1:0] Wgt_9_521,input [WEIGHT_SIZE-1:0] Wgt_9_522,input [WEIGHT_SIZE-1:0] Wgt_9_523,input [WEIGHT_SIZE-1:0] Wgt_9_524,input [WEIGHT_SIZE-1:0] Wgt_9_525,input [WEIGHT_SIZE-1:0] Wgt_9_526,input [WEIGHT_SIZE-1:0] Wgt_9_527,input [WEIGHT_SIZE-1:0] Wgt_9_528,input [WEIGHT_SIZE-1:0] Wgt_9_529,input [WEIGHT_SIZE-1:0] Wgt_9_530,input [WEIGHT_SIZE-1:0] Wgt_9_531,input [WEIGHT_SIZE-1:0] Wgt_9_532,input [WEIGHT_SIZE-1:0] Wgt_9_533,input [WEIGHT_SIZE-1:0] Wgt_9_534,input [WEIGHT_SIZE-1:0] Wgt_9_535,input [WEIGHT_SIZE-1:0] Wgt_9_536,input [WEIGHT_SIZE-1:0] Wgt_9_537,input [WEIGHT_SIZE-1:0] Wgt_9_538,input [WEIGHT_SIZE-1:0] Wgt_9_539,input [WEIGHT_SIZE-1:0] Wgt_9_540,input [WEIGHT_SIZE-1:0] Wgt_9_541,input [WEIGHT_SIZE-1:0] Wgt_9_542,input [WEIGHT_SIZE-1:0] Wgt_9_543,input [WEIGHT_SIZE-1:0] Wgt_9_544,input [WEIGHT_SIZE-1:0] Wgt_9_545,input [WEIGHT_SIZE-1:0] Wgt_9_546,input [WEIGHT_SIZE-1:0] Wgt_9_547,input [WEIGHT_SIZE-1:0] Wgt_9_548,input [WEIGHT_SIZE-1:0] Wgt_9_549,input [WEIGHT_SIZE-1:0] Wgt_9_550,input [WEIGHT_SIZE-1:0] Wgt_9_551,input [WEIGHT_SIZE-1:0] Wgt_9_552,input [WEIGHT_SIZE-1:0] Wgt_9_553,input [WEIGHT_SIZE-1:0] Wgt_9_554,input [WEIGHT_SIZE-1:0] Wgt_9_555,input [WEIGHT_SIZE-1:0] Wgt_9_556,input [WEIGHT_SIZE-1:0] Wgt_9_557,input [WEIGHT_SIZE-1:0] Wgt_9_558,input [WEIGHT_SIZE-1:0] Wgt_9_559,input [WEIGHT_SIZE-1:0] Wgt_9_560,input [WEIGHT_SIZE-1:0] Wgt_9_561,input [WEIGHT_SIZE-1:0] Wgt_9_562,input [WEIGHT_SIZE-1:0] Wgt_9_563,input [WEIGHT_SIZE-1:0] Wgt_9_564,input [WEIGHT_SIZE-1:0] Wgt_9_565,input [WEIGHT_SIZE-1:0] Wgt_9_566,input [WEIGHT_SIZE-1:0] Wgt_9_567,input [WEIGHT_SIZE-1:0] Wgt_9_568,input [WEIGHT_SIZE-1:0] Wgt_9_569,input [WEIGHT_SIZE-1:0] Wgt_9_570,input [WEIGHT_SIZE-1:0] Wgt_9_571,input [WEIGHT_SIZE-1:0] Wgt_9_572,input [WEIGHT_SIZE-1:0] Wgt_9_573,input [WEIGHT_SIZE-1:0] Wgt_9_574,input [WEIGHT_SIZE-1:0] Wgt_9_575,input [WEIGHT_SIZE-1:0] Wgt_9_576,input [WEIGHT_SIZE-1:0] Wgt_9_577,input [WEIGHT_SIZE-1:0] Wgt_9_578,input [WEIGHT_SIZE-1:0] Wgt_9_579,input [WEIGHT_SIZE-1:0] Wgt_9_580,input [WEIGHT_SIZE-1:0] Wgt_9_581,input [WEIGHT_SIZE-1:0] Wgt_9_582,input [WEIGHT_SIZE-1:0] Wgt_9_583,input [WEIGHT_SIZE-1:0] Wgt_9_584,input [WEIGHT_SIZE-1:0] Wgt_9_585,input [WEIGHT_SIZE-1:0] Wgt_9_586,input [WEIGHT_SIZE-1:0] Wgt_9_587,input [WEIGHT_SIZE-1:0] Wgt_9_588,input [WEIGHT_SIZE-1:0] Wgt_9_589,input [WEIGHT_SIZE-1:0] Wgt_9_590,input [WEIGHT_SIZE-1:0] Wgt_9_591,input [WEIGHT_SIZE-1:0] Wgt_9_592,input [WEIGHT_SIZE-1:0] Wgt_9_593,input [WEIGHT_SIZE-1:0] Wgt_9_594,input [WEIGHT_SIZE-1:0] Wgt_9_595,input [WEIGHT_SIZE-1:0] Wgt_9_596,input [WEIGHT_SIZE-1:0] Wgt_9_597,input [WEIGHT_SIZE-1:0] Wgt_9_598,input [WEIGHT_SIZE-1:0] Wgt_9_599,input [WEIGHT_SIZE-1:0] Wgt_9_600,input [WEIGHT_SIZE-1:0] Wgt_9_601,input [WEIGHT_SIZE-1:0] Wgt_9_602,input [WEIGHT_SIZE-1:0] Wgt_9_603,input [WEIGHT_SIZE-1:0] Wgt_9_604,input [WEIGHT_SIZE-1:0] Wgt_9_605,input [WEIGHT_SIZE-1:0] Wgt_9_606,input [WEIGHT_SIZE-1:0] Wgt_9_607,input [WEIGHT_SIZE-1:0] Wgt_9_608,input [WEIGHT_SIZE-1:0] Wgt_9_609,input [WEIGHT_SIZE-1:0] Wgt_9_610,input [WEIGHT_SIZE-1:0] Wgt_9_611,input [WEIGHT_SIZE-1:0] Wgt_9_612,input [WEIGHT_SIZE-1:0] Wgt_9_613,input [WEIGHT_SIZE-1:0] Wgt_9_614,input [WEIGHT_SIZE-1:0] Wgt_9_615,input [WEIGHT_SIZE-1:0] Wgt_9_616,input [WEIGHT_SIZE-1:0] Wgt_9_617,input [WEIGHT_SIZE-1:0] Wgt_9_618,input [WEIGHT_SIZE-1:0] Wgt_9_619,input [WEIGHT_SIZE-1:0] Wgt_9_620,input [WEIGHT_SIZE-1:0] Wgt_9_621,input [WEIGHT_SIZE-1:0] Wgt_9_622,input [WEIGHT_SIZE-1:0] Wgt_9_623,input [WEIGHT_SIZE-1:0] Wgt_9_624,input [WEIGHT_SIZE-1:0] Wgt_9_625,input [WEIGHT_SIZE-1:0] Wgt_9_626,input [WEIGHT_SIZE-1:0] Wgt_9_627,input [WEIGHT_SIZE-1:0] Wgt_9_628,input [WEIGHT_SIZE-1:0] Wgt_9_629,input [WEIGHT_SIZE-1:0] Wgt_9_630,input [WEIGHT_SIZE-1:0] Wgt_9_631,input [WEIGHT_SIZE-1:0] Wgt_9_632,input [WEIGHT_SIZE-1:0] Wgt_9_633,input [WEIGHT_SIZE-1:0] Wgt_9_634,input [WEIGHT_SIZE-1:0] Wgt_9_635,input [WEIGHT_SIZE-1:0] Wgt_9_636,input [WEIGHT_SIZE-1:0] Wgt_9_637,input [WEIGHT_SIZE-1:0] Wgt_9_638,input [WEIGHT_SIZE-1:0] Wgt_9_639,input [WEIGHT_SIZE-1:0] Wgt_9_640,input [WEIGHT_SIZE-1:0] Wgt_9_641,input [WEIGHT_SIZE-1:0] Wgt_9_642,input [WEIGHT_SIZE-1:0] Wgt_9_643,input [WEIGHT_SIZE-1:0] Wgt_9_644,input [WEIGHT_SIZE-1:0] Wgt_9_645,input [WEIGHT_SIZE-1:0] Wgt_9_646,input [WEIGHT_SIZE-1:0] Wgt_9_647,input [WEIGHT_SIZE-1:0] Wgt_9_648,input [WEIGHT_SIZE-1:0] Wgt_9_649,input [WEIGHT_SIZE-1:0] Wgt_9_650,input [WEIGHT_SIZE-1:0] Wgt_9_651,input [WEIGHT_SIZE-1:0] Wgt_9_652,input [WEIGHT_SIZE-1:0] Wgt_9_653,input [WEIGHT_SIZE-1:0] Wgt_9_654,input [WEIGHT_SIZE-1:0] Wgt_9_655,input [WEIGHT_SIZE-1:0] Wgt_9_656,input [WEIGHT_SIZE-1:0] Wgt_9_657,input [WEIGHT_SIZE-1:0] Wgt_9_658,input [WEIGHT_SIZE-1:0] Wgt_9_659,input [WEIGHT_SIZE-1:0] Wgt_9_660,input [WEIGHT_SIZE-1:0] Wgt_9_661,input [WEIGHT_SIZE-1:0] Wgt_9_662,input [WEIGHT_SIZE-1:0] Wgt_9_663,input [WEIGHT_SIZE-1:0] Wgt_9_664,input [WEIGHT_SIZE-1:0] Wgt_9_665,input [WEIGHT_SIZE-1:0] Wgt_9_666,input [WEIGHT_SIZE-1:0] Wgt_9_667,input [WEIGHT_SIZE-1:0] Wgt_9_668,input [WEIGHT_SIZE-1:0] Wgt_9_669,input [WEIGHT_SIZE-1:0] Wgt_9_670,input [WEIGHT_SIZE-1:0] Wgt_9_671,input [WEIGHT_SIZE-1:0] Wgt_9_672,input [WEIGHT_SIZE-1:0] Wgt_9_673,input [WEIGHT_SIZE-1:0] Wgt_9_674,input [WEIGHT_SIZE-1:0] Wgt_9_675,input [WEIGHT_SIZE-1:0] Wgt_9_676,input [WEIGHT_SIZE-1:0] Wgt_9_677,input [WEIGHT_SIZE-1:0] Wgt_9_678,input [WEIGHT_SIZE-1:0] Wgt_9_679,input [WEIGHT_SIZE-1:0] Wgt_9_680,input [WEIGHT_SIZE-1:0] Wgt_9_681,input [WEIGHT_SIZE-1:0] Wgt_9_682,input [WEIGHT_SIZE-1:0] Wgt_9_683,input [WEIGHT_SIZE-1:0] Wgt_9_684,input [WEIGHT_SIZE-1:0] Wgt_9_685,input [WEIGHT_SIZE-1:0] Wgt_9_686,input [WEIGHT_SIZE-1:0] Wgt_9_687,input [WEIGHT_SIZE-1:0] Wgt_9_688,input [WEIGHT_SIZE-1:0] Wgt_9_689,input [WEIGHT_SIZE-1:0] Wgt_9_690,input [WEIGHT_SIZE-1:0] Wgt_9_691,input [WEIGHT_SIZE-1:0] Wgt_9_692,input [WEIGHT_SIZE-1:0] Wgt_9_693,input [WEIGHT_SIZE-1:0] Wgt_9_694,input [WEIGHT_SIZE-1:0] Wgt_9_695,input [WEIGHT_SIZE-1:0] Wgt_9_696,input [WEIGHT_SIZE-1:0] Wgt_9_697,input [WEIGHT_SIZE-1:0] Wgt_9_698,input [WEIGHT_SIZE-1:0] Wgt_9_699,input [WEIGHT_SIZE-1:0] Wgt_9_700,input [WEIGHT_SIZE-1:0] Wgt_9_701,input [WEIGHT_SIZE-1:0] Wgt_9_702,input [WEIGHT_SIZE-1:0] Wgt_9_703,input [WEIGHT_SIZE-1:0] Wgt_9_704,input [WEIGHT_SIZE-1:0] Wgt_9_705,input [WEIGHT_SIZE-1:0] Wgt_9_706,input [WEIGHT_SIZE-1:0] Wgt_9_707,input [WEIGHT_SIZE-1:0] Wgt_9_708,input [WEIGHT_SIZE-1:0] Wgt_9_709,input [WEIGHT_SIZE-1:0] Wgt_9_710,input [WEIGHT_SIZE-1:0] Wgt_9_711,input [WEIGHT_SIZE-1:0] Wgt_9_712,input [WEIGHT_SIZE-1:0] Wgt_9_713,input [WEIGHT_SIZE-1:0] Wgt_9_714,input [WEIGHT_SIZE-1:0] Wgt_9_715,input [WEIGHT_SIZE-1:0] Wgt_9_716,input [WEIGHT_SIZE-1:0] Wgt_9_717,input [WEIGHT_SIZE-1:0] Wgt_9_718,input [WEIGHT_SIZE-1:0] Wgt_9_719,input [WEIGHT_SIZE-1:0] Wgt_9_720,input [WEIGHT_SIZE-1:0] Wgt_9_721,input [WEIGHT_SIZE-1:0] Wgt_9_722,input [WEIGHT_SIZE-1:0] Wgt_9_723,input [WEIGHT_SIZE-1:0] Wgt_9_724,input [WEIGHT_SIZE-1:0] Wgt_9_725,input [WEIGHT_SIZE-1:0] Wgt_9_726,input [WEIGHT_SIZE-1:0] Wgt_9_727,input [WEIGHT_SIZE-1:0] Wgt_9_728,input [WEIGHT_SIZE-1:0] Wgt_9_729,input [WEIGHT_SIZE-1:0] Wgt_9_730,input [WEIGHT_SIZE-1:0] Wgt_9_731,input [WEIGHT_SIZE-1:0] Wgt_9_732,input [WEIGHT_SIZE-1:0] Wgt_9_733,input [WEIGHT_SIZE-1:0] Wgt_9_734,input [WEIGHT_SIZE-1:0] Wgt_9_735,input [WEIGHT_SIZE-1:0] Wgt_9_736,input [WEIGHT_SIZE-1:0] Wgt_9_737,input [WEIGHT_SIZE-1:0] Wgt_9_738,input [WEIGHT_SIZE-1:0] Wgt_9_739,input [WEIGHT_SIZE-1:0] Wgt_9_740,input [WEIGHT_SIZE-1:0] Wgt_9_741,input [WEIGHT_SIZE-1:0] Wgt_9_742,input [WEIGHT_SIZE-1:0] Wgt_9_743,input [WEIGHT_SIZE-1:0] Wgt_9_744,input [WEIGHT_SIZE-1:0] Wgt_9_745,input [WEIGHT_SIZE-1:0] Wgt_9_746,input [WEIGHT_SIZE-1:0] Wgt_9_747,input [WEIGHT_SIZE-1:0] Wgt_9_748,input [WEIGHT_SIZE-1:0] Wgt_9_749,input [WEIGHT_SIZE-1:0] Wgt_9_750,input [WEIGHT_SIZE-1:0] Wgt_9_751,input [WEIGHT_SIZE-1:0] Wgt_9_752,input [WEIGHT_SIZE-1:0] Wgt_9_753,input [WEIGHT_SIZE-1:0] Wgt_9_754,input [WEIGHT_SIZE-1:0] Wgt_9_755,input [WEIGHT_SIZE-1:0] Wgt_9_756,input [WEIGHT_SIZE-1:0] Wgt_9_757,input [WEIGHT_SIZE-1:0] Wgt_9_758,input [WEIGHT_SIZE-1:0] Wgt_9_759,input [WEIGHT_SIZE-1:0] Wgt_9_760,input [WEIGHT_SIZE-1:0] Wgt_9_761,input [WEIGHT_SIZE-1:0] Wgt_9_762,input [WEIGHT_SIZE-1:0] Wgt_9_763,input [WEIGHT_SIZE-1:0] Wgt_9_764,input [WEIGHT_SIZE-1:0] Wgt_9_765,input [WEIGHT_SIZE-1:0] Wgt_9_766,input [WEIGHT_SIZE-1:0] Wgt_9_767,input [WEIGHT_SIZE-1:0] Wgt_9_768,input [WEIGHT_SIZE-1:0] Wgt_9_769,input [WEIGHT_SIZE-1:0] Wgt_9_770,input [WEIGHT_SIZE-1:0] Wgt_9_771,input [WEIGHT_SIZE-1:0] Wgt_9_772,input [WEIGHT_SIZE-1:0] Wgt_9_773,input [WEIGHT_SIZE-1:0] Wgt_9_774,input [WEIGHT_SIZE-1:0] Wgt_9_775,input [WEIGHT_SIZE-1:0] Wgt_9_776,input [WEIGHT_SIZE-1:0] Wgt_9_777,input [WEIGHT_SIZE-1:0] Wgt_9_778,input [WEIGHT_SIZE-1:0] Wgt_9_779,input [WEIGHT_SIZE-1:0] Wgt_9_780,input [WEIGHT_SIZE-1:0] Wgt_9_781,input [WEIGHT_SIZE-1:0] Wgt_9_782,input [WEIGHT_SIZE-1:0] Wgt_9_783,input [WEIGHT_SIZE-1:0] Wgt_9_784,
input [PIXEL_SIZE-1:0] Pix_0,input [PIXEL_SIZE-1:0] Pix_1,input [PIXEL_SIZE-1:0] Pix_2,input [PIXEL_SIZE-1:0] Pix_3,input [PIXEL_SIZE-1:0] Pix_4,input [PIXEL_SIZE-1:0] Pix_5,input [PIXEL_SIZE-1:0] Pix_6,input [PIXEL_SIZE-1:0] Pix_7,input [PIXEL_SIZE-1:0] Pix_8,input [PIXEL_SIZE-1:0] Pix_9,input [PIXEL_SIZE-1:0] Pix_10,input [PIXEL_SIZE-1:0] Pix_11,input [PIXEL_SIZE-1:0] Pix_12,input [PIXEL_SIZE-1:0] Pix_13,input [PIXEL_SIZE-1:0] Pix_14,input [PIXEL_SIZE-1:0] Pix_15,input [PIXEL_SIZE-1:0] Pix_16,input [PIXEL_SIZE-1:0] Pix_17,input [PIXEL_SIZE-1:0] Pix_18,input [PIXEL_SIZE-1:0] Pix_19,input [PIXEL_SIZE-1:0] Pix_20,input [PIXEL_SIZE-1:0] Pix_21,input [PIXEL_SIZE-1:0] Pix_22,input [PIXEL_SIZE-1:0] Pix_23,input [PIXEL_SIZE-1:0] Pix_24,input [PIXEL_SIZE-1:0] Pix_25,input [PIXEL_SIZE-1:0] Pix_26,input [PIXEL_SIZE-1:0] Pix_27,input [PIXEL_SIZE-1:0] Pix_28,input [PIXEL_SIZE-1:0] Pix_29,input [PIXEL_SIZE-1:0] Pix_30,input [PIXEL_SIZE-1:0] Pix_31,input [PIXEL_SIZE-1:0] Pix_32,input [PIXEL_SIZE-1:0] Pix_33,input [PIXEL_SIZE-1:0] Pix_34,input [PIXEL_SIZE-1:0] Pix_35,input [PIXEL_SIZE-1:0] Pix_36,input [PIXEL_SIZE-1:0] Pix_37,input [PIXEL_SIZE-1:0] Pix_38,input [PIXEL_SIZE-1:0] Pix_39,input [PIXEL_SIZE-1:0] Pix_40,input [PIXEL_SIZE-1:0] Pix_41,input [PIXEL_SIZE-1:0] Pix_42,input [PIXEL_SIZE-1:0] Pix_43,input [PIXEL_SIZE-1:0] Pix_44,input [PIXEL_SIZE-1:0] Pix_45,input [PIXEL_SIZE-1:0] Pix_46,input [PIXEL_SIZE-1:0] Pix_47,input [PIXEL_SIZE-1:0] Pix_48,input [PIXEL_SIZE-1:0] Pix_49,input [PIXEL_SIZE-1:0] Pix_50,input [PIXEL_SIZE-1:0] Pix_51,input [PIXEL_SIZE-1:0] Pix_52,input [PIXEL_SIZE-1:0] Pix_53,input [PIXEL_SIZE-1:0] Pix_54,input [PIXEL_SIZE-1:0] Pix_55,input [PIXEL_SIZE-1:0] Pix_56,input [PIXEL_SIZE-1:0] Pix_57,input [PIXEL_SIZE-1:0] Pix_58,input [PIXEL_SIZE-1:0] Pix_59,input [PIXEL_SIZE-1:0] Pix_60,input [PIXEL_SIZE-1:0] Pix_61,input [PIXEL_SIZE-1:0] Pix_62,input [PIXEL_SIZE-1:0] Pix_63,input [PIXEL_SIZE-1:0] Pix_64,input [PIXEL_SIZE-1:0] Pix_65,input [PIXEL_SIZE-1:0] Pix_66,input [PIXEL_SIZE-1:0] Pix_67,input [PIXEL_SIZE-1:0] Pix_68,input [PIXEL_SIZE-1:0] Pix_69,input [PIXEL_SIZE-1:0] Pix_70,input [PIXEL_SIZE-1:0] Pix_71,input [PIXEL_SIZE-1:0] Pix_72,input [PIXEL_SIZE-1:0] Pix_73,input [PIXEL_SIZE-1:0] Pix_74,input [PIXEL_SIZE-1:0] Pix_75,input [PIXEL_SIZE-1:0] Pix_76,input [PIXEL_SIZE-1:0] Pix_77,input [PIXEL_SIZE-1:0] Pix_78,input [PIXEL_SIZE-1:0] Pix_79,input [PIXEL_SIZE-1:0] Pix_80,input [PIXEL_SIZE-1:0] Pix_81,input [PIXEL_SIZE-1:0] Pix_82,input [PIXEL_SIZE-1:0] Pix_83,input [PIXEL_SIZE-1:0] Pix_84,input [PIXEL_SIZE-1:0] Pix_85,input [PIXEL_SIZE-1:0] Pix_86,input [PIXEL_SIZE-1:0] Pix_87,input [PIXEL_SIZE-1:0] Pix_88,input [PIXEL_SIZE-1:0] Pix_89,input [PIXEL_SIZE-1:0] Pix_90,input [PIXEL_SIZE-1:0] Pix_91,input [PIXEL_SIZE-1:0] Pix_92,input [PIXEL_SIZE-1:0] Pix_93,input [PIXEL_SIZE-1:0] Pix_94,input [PIXEL_SIZE-1:0] Pix_95,input [PIXEL_SIZE-1:0] Pix_96,input [PIXEL_SIZE-1:0] Pix_97,input [PIXEL_SIZE-1:0] Pix_98,input [PIXEL_SIZE-1:0] Pix_99,input [PIXEL_SIZE-1:0] Pix_100,input [PIXEL_SIZE-1:0] Pix_101,input [PIXEL_SIZE-1:0] Pix_102,input [PIXEL_SIZE-1:0] Pix_103,input [PIXEL_SIZE-1:0] Pix_104,input [PIXEL_SIZE-1:0] Pix_105,input [PIXEL_SIZE-1:0] Pix_106,input [PIXEL_SIZE-1:0] Pix_107,input [PIXEL_SIZE-1:0] Pix_108,input [PIXEL_SIZE-1:0] Pix_109,input [PIXEL_SIZE-1:0] Pix_110,input [PIXEL_SIZE-1:0] Pix_111,input [PIXEL_SIZE-1:0] Pix_112,input [PIXEL_SIZE-1:0] Pix_113,input [PIXEL_SIZE-1:0] Pix_114,input [PIXEL_SIZE-1:0] Pix_115,input [PIXEL_SIZE-1:0] Pix_116,input [PIXEL_SIZE-1:0] Pix_117,input [PIXEL_SIZE-1:0] Pix_118,input [PIXEL_SIZE-1:0] Pix_119,input [PIXEL_SIZE-1:0] Pix_120,input [PIXEL_SIZE-1:0] Pix_121,input [PIXEL_SIZE-1:0] Pix_122,input [PIXEL_SIZE-1:0] Pix_123,input [PIXEL_SIZE-1:0] Pix_124,input [PIXEL_SIZE-1:0] Pix_125,input [PIXEL_SIZE-1:0] Pix_126,input [PIXEL_SIZE-1:0] Pix_127,input [PIXEL_SIZE-1:0] Pix_128,input [PIXEL_SIZE-1:0] Pix_129,input [PIXEL_SIZE-1:0] Pix_130,input [PIXEL_SIZE-1:0] Pix_131,input [PIXEL_SIZE-1:0] Pix_132,input [PIXEL_SIZE-1:0] Pix_133,input [PIXEL_SIZE-1:0] Pix_134,input [PIXEL_SIZE-1:0] Pix_135,input [PIXEL_SIZE-1:0] Pix_136,input [PIXEL_SIZE-1:0] Pix_137,input [PIXEL_SIZE-1:0] Pix_138,input [PIXEL_SIZE-1:0] Pix_139,input [PIXEL_SIZE-1:0] Pix_140,input [PIXEL_SIZE-1:0] Pix_141,input [PIXEL_SIZE-1:0] Pix_142,input [PIXEL_SIZE-1:0] Pix_143,input [PIXEL_SIZE-1:0] Pix_144,input [PIXEL_SIZE-1:0] Pix_145,input [PIXEL_SIZE-1:0] Pix_146,input [PIXEL_SIZE-1:0] Pix_147,input [PIXEL_SIZE-1:0] Pix_148,input [PIXEL_SIZE-1:0] Pix_149,input [PIXEL_SIZE-1:0] Pix_150,input [PIXEL_SIZE-1:0] Pix_151,input [PIXEL_SIZE-1:0] Pix_152,input [PIXEL_SIZE-1:0] Pix_153,input [PIXEL_SIZE-1:0] Pix_154,input [PIXEL_SIZE-1:0] Pix_155,input [PIXEL_SIZE-1:0] Pix_156,input [PIXEL_SIZE-1:0] Pix_157,input [PIXEL_SIZE-1:0] Pix_158,input [PIXEL_SIZE-1:0] Pix_159,input [PIXEL_SIZE-1:0] Pix_160,input [PIXEL_SIZE-1:0] Pix_161,input [PIXEL_SIZE-1:0] Pix_162,input [PIXEL_SIZE-1:0] Pix_163,input [PIXEL_SIZE-1:0] Pix_164,input [PIXEL_SIZE-1:0] Pix_165,input [PIXEL_SIZE-1:0] Pix_166,input [PIXEL_SIZE-1:0] Pix_167,input [PIXEL_SIZE-1:0] Pix_168,input [PIXEL_SIZE-1:0] Pix_169,input [PIXEL_SIZE-1:0] Pix_170,input [PIXEL_SIZE-1:0] Pix_171,input [PIXEL_SIZE-1:0] Pix_172,input [PIXEL_SIZE-1:0] Pix_173,input [PIXEL_SIZE-1:0] Pix_174,input [PIXEL_SIZE-1:0] Pix_175,input [PIXEL_SIZE-1:0] Pix_176,input [PIXEL_SIZE-1:0] Pix_177,input [PIXEL_SIZE-1:0] Pix_178,input [PIXEL_SIZE-1:0] Pix_179,input [PIXEL_SIZE-1:0] Pix_180,input [PIXEL_SIZE-1:0] Pix_181,input [PIXEL_SIZE-1:0] Pix_182,input [PIXEL_SIZE-1:0] Pix_183,input [PIXEL_SIZE-1:0] Pix_184,input [PIXEL_SIZE-1:0] Pix_185,input [PIXEL_SIZE-1:0] Pix_186,input [PIXEL_SIZE-1:0] Pix_187,input [PIXEL_SIZE-1:0] Pix_188,input [PIXEL_SIZE-1:0] Pix_189,input [PIXEL_SIZE-1:0] Pix_190,input [PIXEL_SIZE-1:0] Pix_191,input [PIXEL_SIZE-1:0] Pix_192,input [PIXEL_SIZE-1:0] Pix_193,input [PIXEL_SIZE-1:0] Pix_194,input [PIXEL_SIZE-1:0] Pix_195,input [PIXEL_SIZE-1:0] Pix_196,input [PIXEL_SIZE-1:0] Pix_197,input [PIXEL_SIZE-1:0] Pix_198,input [PIXEL_SIZE-1:0] Pix_199,input [PIXEL_SIZE-1:0] Pix_200,input [PIXEL_SIZE-1:0] Pix_201,input [PIXEL_SIZE-1:0] Pix_202,input [PIXEL_SIZE-1:0] Pix_203,input [PIXEL_SIZE-1:0] Pix_204,input [PIXEL_SIZE-1:0] Pix_205,input [PIXEL_SIZE-1:0] Pix_206,input [PIXEL_SIZE-1:0] Pix_207,input [PIXEL_SIZE-1:0] Pix_208,input [PIXEL_SIZE-1:0] Pix_209,input [PIXEL_SIZE-1:0] Pix_210,input [PIXEL_SIZE-1:0] Pix_211,input [PIXEL_SIZE-1:0] Pix_212,input [PIXEL_SIZE-1:0] Pix_213,input [PIXEL_SIZE-1:0] Pix_214,input [PIXEL_SIZE-1:0] Pix_215,input [PIXEL_SIZE-1:0] Pix_216,input [PIXEL_SIZE-1:0] Pix_217,input [PIXEL_SIZE-1:0] Pix_218,input [PIXEL_SIZE-1:0] Pix_219,input [PIXEL_SIZE-1:0] Pix_220,input [PIXEL_SIZE-1:0] Pix_221,input [PIXEL_SIZE-1:0] Pix_222,input [PIXEL_SIZE-1:0] Pix_223,input [PIXEL_SIZE-1:0] Pix_224,input [PIXEL_SIZE-1:0] Pix_225,input [PIXEL_SIZE-1:0] Pix_226,input [PIXEL_SIZE-1:0] Pix_227,input [PIXEL_SIZE-1:0] Pix_228,input [PIXEL_SIZE-1:0] Pix_229,input [PIXEL_SIZE-1:0] Pix_230,input [PIXEL_SIZE-1:0] Pix_231,input [PIXEL_SIZE-1:0] Pix_232,input [PIXEL_SIZE-1:0] Pix_233,input [PIXEL_SIZE-1:0] Pix_234,input [PIXEL_SIZE-1:0] Pix_235,input [PIXEL_SIZE-1:0] Pix_236,input [PIXEL_SIZE-1:0] Pix_237,input [PIXEL_SIZE-1:0] Pix_238,input [PIXEL_SIZE-1:0] Pix_239,input [PIXEL_SIZE-1:0] Pix_240,input [PIXEL_SIZE-1:0] Pix_241,input [PIXEL_SIZE-1:0] Pix_242,input [PIXEL_SIZE-1:0] Pix_243,input [PIXEL_SIZE-1:0] Pix_244,input [PIXEL_SIZE-1:0] Pix_245,input [PIXEL_SIZE-1:0] Pix_246,input [PIXEL_SIZE-1:0] Pix_247,input [PIXEL_SIZE-1:0] Pix_248,input [PIXEL_SIZE-1:0] Pix_249,input [PIXEL_SIZE-1:0] Pix_250,input [PIXEL_SIZE-1:0] Pix_251,input [PIXEL_SIZE-1:0] Pix_252,input [PIXEL_SIZE-1:0] Pix_253,input [PIXEL_SIZE-1:0] Pix_254,input [PIXEL_SIZE-1:0] Pix_255,input [PIXEL_SIZE-1:0] Pix_256,input [PIXEL_SIZE-1:0] Pix_257,input [PIXEL_SIZE-1:0] Pix_258,input [PIXEL_SIZE-1:0] Pix_259,input [PIXEL_SIZE-1:0] Pix_260,input [PIXEL_SIZE-1:0] Pix_261,input [PIXEL_SIZE-1:0] Pix_262,input [PIXEL_SIZE-1:0] Pix_263,input [PIXEL_SIZE-1:0] Pix_264,input [PIXEL_SIZE-1:0] Pix_265,input [PIXEL_SIZE-1:0] Pix_266,input [PIXEL_SIZE-1:0] Pix_267,input [PIXEL_SIZE-1:0] Pix_268,input [PIXEL_SIZE-1:0] Pix_269,input [PIXEL_SIZE-1:0] Pix_270,input [PIXEL_SIZE-1:0] Pix_271,input [PIXEL_SIZE-1:0] Pix_272,input [PIXEL_SIZE-1:0] Pix_273,input [PIXEL_SIZE-1:0] Pix_274,input [PIXEL_SIZE-1:0] Pix_275,input [PIXEL_SIZE-1:0] Pix_276,input [PIXEL_SIZE-1:0] Pix_277,input [PIXEL_SIZE-1:0] Pix_278,input [PIXEL_SIZE-1:0] Pix_279,input [PIXEL_SIZE-1:0] Pix_280,input [PIXEL_SIZE-1:0] Pix_281,input [PIXEL_SIZE-1:0] Pix_282,input [PIXEL_SIZE-1:0] Pix_283,input [PIXEL_SIZE-1:0] Pix_284,input [PIXEL_SIZE-1:0] Pix_285,input [PIXEL_SIZE-1:0] Pix_286,input [PIXEL_SIZE-1:0] Pix_287,input [PIXEL_SIZE-1:0] Pix_288,input [PIXEL_SIZE-1:0] Pix_289,input [PIXEL_SIZE-1:0] Pix_290,input [PIXEL_SIZE-1:0] Pix_291,input [PIXEL_SIZE-1:0] Pix_292,input [PIXEL_SIZE-1:0] Pix_293,input [PIXEL_SIZE-1:0] Pix_294,input [PIXEL_SIZE-1:0] Pix_295,input [PIXEL_SIZE-1:0] Pix_296,input [PIXEL_SIZE-1:0] Pix_297,input [PIXEL_SIZE-1:0] Pix_298,input [PIXEL_SIZE-1:0] Pix_299,input [PIXEL_SIZE-1:0] Pix_300,input [PIXEL_SIZE-1:0] Pix_301,input [PIXEL_SIZE-1:0] Pix_302,input [PIXEL_SIZE-1:0] Pix_303,input [PIXEL_SIZE-1:0] Pix_304,input [PIXEL_SIZE-1:0] Pix_305,input [PIXEL_SIZE-1:0] Pix_306,input [PIXEL_SIZE-1:0] Pix_307,input [PIXEL_SIZE-1:0] Pix_308,input [PIXEL_SIZE-1:0] Pix_309,input [PIXEL_SIZE-1:0] Pix_310,input [PIXEL_SIZE-1:0] Pix_311,input [PIXEL_SIZE-1:0] Pix_312,input [PIXEL_SIZE-1:0] Pix_313,input [PIXEL_SIZE-1:0] Pix_314,input [PIXEL_SIZE-1:0] Pix_315,input [PIXEL_SIZE-1:0] Pix_316,input [PIXEL_SIZE-1:0] Pix_317,input [PIXEL_SIZE-1:0] Pix_318,input [PIXEL_SIZE-1:0] Pix_319,input [PIXEL_SIZE-1:0] Pix_320,input [PIXEL_SIZE-1:0] Pix_321,input [PIXEL_SIZE-1:0] Pix_322,input [PIXEL_SIZE-1:0] Pix_323,input [PIXEL_SIZE-1:0] Pix_324,input [PIXEL_SIZE-1:0] Pix_325,input [PIXEL_SIZE-1:0] Pix_326,input [PIXEL_SIZE-1:0] Pix_327,input [PIXEL_SIZE-1:0] Pix_328,input [PIXEL_SIZE-1:0] Pix_329,input [PIXEL_SIZE-1:0] Pix_330,input [PIXEL_SIZE-1:0] Pix_331,input [PIXEL_SIZE-1:0] Pix_332,input [PIXEL_SIZE-1:0] Pix_333,input [PIXEL_SIZE-1:0] Pix_334,input [PIXEL_SIZE-1:0] Pix_335,input [PIXEL_SIZE-1:0] Pix_336,input [PIXEL_SIZE-1:0] Pix_337,input [PIXEL_SIZE-1:0] Pix_338,input [PIXEL_SIZE-1:0] Pix_339,input [PIXEL_SIZE-1:0] Pix_340,input [PIXEL_SIZE-1:0] Pix_341,input [PIXEL_SIZE-1:0] Pix_342,input [PIXEL_SIZE-1:0] Pix_343,input [PIXEL_SIZE-1:0] Pix_344,input [PIXEL_SIZE-1:0] Pix_345,input [PIXEL_SIZE-1:0] Pix_346,input [PIXEL_SIZE-1:0] Pix_347,input [PIXEL_SIZE-1:0] Pix_348,input [PIXEL_SIZE-1:0] Pix_349,input [PIXEL_SIZE-1:0] Pix_350,input [PIXEL_SIZE-1:0] Pix_351,input [PIXEL_SIZE-1:0] Pix_352,input [PIXEL_SIZE-1:0] Pix_353,input [PIXEL_SIZE-1:0] Pix_354,input [PIXEL_SIZE-1:0] Pix_355,input [PIXEL_SIZE-1:0] Pix_356,input [PIXEL_SIZE-1:0] Pix_357,input [PIXEL_SIZE-1:0] Pix_358,input [PIXEL_SIZE-1:0] Pix_359,input [PIXEL_SIZE-1:0] Pix_360,input [PIXEL_SIZE-1:0] Pix_361,input [PIXEL_SIZE-1:0] Pix_362,input [PIXEL_SIZE-1:0] Pix_363,input [PIXEL_SIZE-1:0] Pix_364,input [PIXEL_SIZE-1:0] Pix_365,input [PIXEL_SIZE-1:0] Pix_366,input [PIXEL_SIZE-1:0] Pix_367,input [PIXEL_SIZE-1:0] Pix_368,input [PIXEL_SIZE-1:0] Pix_369,input [PIXEL_SIZE-1:0] Pix_370,input [PIXEL_SIZE-1:0] Pix_371,input [PIXEL_SIZE-1:0] Pix_372,input [PIXEL_SIZE-1:0] Pix_373,input [PIXEL_SIZE-1:0] Pix_374,input [PIXEL_SIZE-1:0] Pix_375,input [PIXEL_SIZE-1:0] Pix_376,input [PIXEL_SIZE-1:0] Pix_377,input [PIXEL_SIZE-1:0] Pix_378,input [PIXEL_SIZE-1:0] Pix_379,input [PIXEL_SIZE-1:0] Pix_380,input [PIXEL_SIZE-1:0] Pix_381,input [PIXEL_SIZE-1:0] Pix_382,input [PIXEL_SIZE-1:0] Pix_383,input [PIXEL_SIZE-1:0] Pix_384,input [PIXEL_SIZE-1:0] Pix_385,input [PIXEL_SIZE-1:0] Pix_386,input [PIXEL_SIZE-1:0] Pix_387,input [PIXEL_SIZE-1:0] Pix_388,input [PIXEL_SIZE-1:0] Pix_389,input [PIXEL_SIZE-1:0] Pix_390,input [PIXEL_SIZE-1:0] Pix_391,input [PIXEL_SIZE-1:0] Pix_392,input [PIXEL_SIZE-1:0] Pix_393,input [PIXEL_SIZE-1:0] Pix_394,input [PIXEL_SIZE-1:0] Pix_395,input [PIXEL_SIZE-1:0] Pix_396,input [PIXEL_SIZE-1:0] Pix_397,input [PIXEL_SIZE-1:0] Pix_398,input [PIXEL_SIZE-1:0] Pix_399,input [PIXEL_SIZE-1:0] Pix_400,input [PIXEL_SIZE-1:0] Pix_401,input [PIXEL_SIZE-1:0] Pix_402,input [PIXEL_SIZE-1:0] Pix_403,input [PIXEL_SIZE-1:0] Pix_404,input [PIXEL_SIZE-1:0] Pix_405,input [PIXEL_SIZE-1:0] Pix_406,input [PIXEL_SIZE-1:0] Pix_407,input [PIXEL_SIZE-1:0] Pix_408,input [PIXEL_SIZE-1:0] Pix_409,input [PIXEL_SIZE-1:0] Pix_410,input [PIXEL_SIZE-1:0] Pix_411,input [PIXEL_SIZE-1:0] Pix_412,input [PIXEL_SIZE-1:0] Pix_413,input [PIXEL_SIZE-1:0] Pix_414,input [PIXEL_SIZE-1:0] Pix_415,input [PIXEL_SIZE-1:0] Pix_416,input [PIXEL_SIZE-1:0] Pix_417,input [PIXEL_SIZE-1:0] Pix_418,input [PIXEL_SIZE-1:0] Pix_419,input [PIXEL_SIZE-1:0] Pix_420,input [PIXEL_SIZE-1:0] Pix_421,input [PIXEL_SIZE-1:0] Pix_422,input [PIXEL_SIZE-1:0] Pix_423,input [PIXEL_SIZE-1:0] Pix_424,input [PIXEL_SIZE-1:0] Pix_425,input [PIXEL_SIZE-1:0] Pix_426,input [PIXEL_SIZE-1:0] Pix_427,input [PIXEL_SIZE-1:0] Pix_428,input [PIXEL_SIZE-1:0] Pix_429,input [PIXEL_SIZE-1:0] Pix_430,input [PIXEL_SIZE-1:0] Pix_431,input [PIXEL_SIZE-1:0] Pix_432,input [PIXEL_SIZE-1:0] Pix_433,input [PIXEL_SIZE-1:0] Pix_434,input [PIXEL_SIZE-1:0] Pix_435,input [PIXEL_SIZE-1:0] Pix_436,input [PIXEL_SIZE-1:0] Pix_437,input [PIXEL_SIZE-1:0] Pix_438,input [PIXEL_SIZE-1:0] Pix_439,input [PIXEL_SIZE-1:0] Pix_440,input [PIXEL_SIZE-1:0] Pix_441,input [PIXEL_SIZE-1:0] Pix_442,input [PIXEL_SIZE-1:0] Pix_443,input [PIXEL_SIZE-1:0] Pix_444,input [PIXEL_SIZE-1:0] Pix_445,input [PIXEL_SIZE-1:0] Pix_446,input [PIXEL_SIZE-1:0] Pix_447,input [PIXEL_SIZE-1:0] Pix_448,input [PIXEL_SIZE-1:0] Pix_449,input [PIXEL_SIZE-1:0] Pix_450,input [PIXEL_SIZE-1:0] Pix_451,input [PIXEL_SIZE-1:0] Pix_452,input [PIXEL_SIZE-1:0] Pix_453,input [PIXEL_SIZE-1:0] Pix_454,input [PIXEL_SIZE-1:0] Pix_455,input [PIXEL_SIZE-1:0] Pix_456,input [PIXEL_SIZE-1:0] Pix_457,input [PIXEL_SIZE-1:0] Pix_458,input [PIXEL_SIZE-1:0] Pix_459,input [PIXEL_SIZE-1:0] Pix_460,input [PIXEL_SIZE-1:0] Pix_461,input [PIXEL_SIZE-1:0] Pix_462,input [PIXEL_SIZE-1:0] Pix_463,input [PIXEL_SIZE-1:0] Pix_464,input [PIXEL_SIZE-1:0] Pix_465,input [PIXEL_SIZE-1:0] Pix_466,input [PIXEL_SIZE-1:0] Pix_467,input [PIXEL_SIZE-1:0] Pix_468,input [PIXEL_SIZE-1:0] Pix_469,input [PIXEL_SIZE-1:0] Pix_470,input [PIXEL_SIZE-1:0] Pix_471,input [PIXEL_SIZE-1:0] Pix_472,input [PIXEL_SIZE-1:0] Pix_473,input [PIXEL_SIZE-1:0] Pix_474,input [PIXEL_SIZE-1:0] Pix_475,input [PIXEL_SIZE-1:0] Pix_476,input [PIXEL_SIZE-1:0] Pix_477,input [PIXEL_SIZE-1:0] Pix_478,input [PIXEL_SIZE-1:0] Pix_479,input [PIXEL_SIZE-1:0] Pix_480,input [PIXEL_SIZE-1:0] Pix_481,input [PIXEL_SIZE-1:0] Pix_482,input [PIXEL_SIZE-1:0] Pix_483,input [PIXEL_SIZE-1:0] Pix_484,input [PIXEL_SIZE-1:0] Pix_485,input [PIXEL_SIZE-1:0] Pix_486,input [PIXEL_SIZE-1:0] Pix_487,input [PIXEL_SIZE-1:0] Pix_488,input [PIXEL_SIZE-1:0] Pix_489,input [PIXEL_SIZE-1:0] Pix_490,input [PIXEL_SIZE-1:0] Pix_491,input [PIXEL_SIZE-1:0] Pix_492,input [PIXEL_SIZE-1:0] Pix_493,input [PIXEL_SIZE-1:0] Pix_494,input [PIXEL_SIZE-1:0] Pix_495,input [PIXEL_SIZE-1:0] Pix_496,input [PIXEL_SIZE-1:0] Pix_497,input [PIXEL_SIZE-1:0] Pix_498,input [PIXEL_SIZE-1:0] Pix_499,input [PIXEL_SIZE-1:0] Pix_500,input [PIXEL_SIZE-1:0] Pix_501,input [PIXEL_SIZE-1:0] Pix_502,input [PIXEL_SIZE-1:0] Pix_503,input [PIXEL_SIZE-1:0] Pix_504,input [PIXEL_SIZE-1:0] Pix_505,input [PIXEL_SIZE-1:0] Pix_506,input [PIXEL_SIZE-1:0] Pix_507,input [PIXEL_SIZE-1:0] Pix_508,input [PIXEL_SIZE-1:0] Pix_509,input [PIXEL_SIZE-1:0] Pix_510,input [PIXEL_SIZE-1:0] Pix_511,input [PIXEL_SIZE-1:0] Pix_512,input [PIXEL_SIZE-1:0] Pix_513,input [PIXEL_SIZE-1:0] Pix_514,input [PIXEL_SIZE-1:0] Pix_515,input [PIXEL_SIZE-1:0] Pix_516,input [PIXEL_SIZE-1:0] Pix_517,input [PIXEL_SIZE-1:0] Pix_518,input [PIXEL_SIZE-1:0] Pix_519,input [PIXEL_SIZE-1:0] Pix_520,input [PIXEL_SIZE-1:0] Pix_521,input [PIXEL_SIZE-1:0] Pix_522,input [PIXEL_SIZE-1:0] Pix_523,input [PIXEL_SIZE-1:0] Pix_524,input [PIXEL_SIZE-1:0] Pix_525,input [PIXEL_SIZE-1:0] Pix_526,input [PIXEL_SIZE-1:0] Pix_527,input [PIXEL_SIZE-1:0] Pix_528,input [PIXEL_SIZE-1:0] Pix_529,input [PIXEL_SIZE-1:0] Pix_530,input [PIXEL_SIZE-1:0] Pix_531,input [PIXEL_SIZE-1:0] Pix_532,input [PIXEL_SIZE-1:0] Pix_533,input [PIXEL_SIZE-1:0] Pix_534,input [PIXEL_SIZE-1:0] Pix_535,input [PIXEL_SIZE-1:0] Pix_536,input [PIXEL_SIZE-1:0] Pix_537,input [PIXEL_SIZE-1:0] Pix_538,input [PIXEL_SIZE-1:0] Pix_539,input [PIXEL_SIZE-1:0] Pix_540,input [PIXEL_SIZE-1:0] Pix_541,input [PIXEL_SIZE-1:0] Pix_542,input [PIXEL_SIZE-1:0] Pix_543,input [PIXEL_SIZE-1:0] Pix_544,input [PIXEL_SIZE-1:0] Pix_545,input [PIXEL_SIZE-1:0] Pix_546,input [PIXEL_SIZE-1:0] Pix_547,input [PIXEL_SIZE-1:0] Pix_548,input [PIXEL_SIZE-1:0] Pix_549,input [PIXEL_SIZE-1:0] Pix_550,input [PIXEL_SIZE-1:0] Pix_551,input [PIXEL_SIZE-1:0] Pix_552,input [PIXEL_SIZE-1:0] Pix_553,input [PIXEL_SIZE-1:0] Pix_554,input [PIXEL_SIZE-1:0] Pix_555,input [PIXEL_SIZE-1:0] Pix_556,input [PIXEL_SIZE-1:0] Pix_557,input [PIXEL_SIZE-1:0] Pix_558,input [PIXEL_SIZE-1:0] Pix_559,input [PIXEL_SIZE-1:0] Pix_560,input [PIXEL_SIZE-1:0] Pix_561,input [PIXEL_SIZE-1:0] Pix_562,input [PIXEL_SIZE-1:0] Pix_563,input [PIXEL_SIZE-1:0] Pix_564,input [PIXEL_SIZE-1:0] Pix_565,input [PIXEL_SIZE-1:0] Pix_566,input [PIXEL_SIZE-1:0] Pix_567,input [PIXEL_SIZE-1:0] Pix_568,input [PIXEL_SIZE-1:0] Pix_569,input [PIXEL_SIZE-1:0] Pix_570,input [PIXEL_SIZE-1:0] Pix_571,input [PIXEL_SIZE-1:0] Pix_572,input [PIXEL_SIZE-1:0] Pix_573,input [PIXEL_SIZE-1:0] Pix_574,input [PIXEL_SIZE-1:0] Pix_575,input [PIXEL_SIZE-1:0] Pix_576,input [PIXEL_SIZE-1:0] Pix_577,input [PIXEL_SIZE-1:0] Pix_578,input [PIXEL_SIZE-1:0] Pix_579,input [PIXEL_SIZE-1:0] Pix_580,input [PIXEL_SIZE-1:0] Pix_581,input [PIXEL_SIZE-1:0] Pix_582,input [PIXEL_SIZE-1:0] Pix_583,input [PIXEL_SIZE-1:0] Pix_584,input [PIXEL_SIZE-1:0] Pix_585,input [PIXEL_SIZE-1:0] Pix_586,input [PIXEL_SIZE-1:0] Pix_587,input [PIXEL_SIZE-1:0] Pix_588,input [PIXEL_SIZE-1:0] Pix_589,input [PIXEL_SIZE-1:0] Pix_590,input [PIXEL_SIZE-1:0] Pix_591,input [PIXEL_SIZE-1:0] Pix_592,input [PIXEL_SIZE-1:0] Pix_593,input [PIXEL_SIZE-1:0] Pix_594,input [PIXEL_SIZE-1:0] Pix_595,input [PIXEL_SIZE-1:0] Pix_596,input [PIXEL_SIZE-1:0] Pix_597,input [PIXEL_SIZE-1:0] Pix_598,input [PIXEL_SIZE-1:0] Pix_599,input [PIXEL_SIZE-1:0] Pix_600,input [PIXEL_SIZE-1:0] Pix_601,input [PIXEL_SIZE-1:0] Pix_602,input [PIXEL_SIZE-1:0] Pix_603,input [PIXEL_SIZE-1:0] Pix_604,input [PIXEL_SIZE-1:0] Pix_605,input [PIXEL_SIZE-1:0] Pix_606,input [PIXEL_SIZE-1:0] Pix_607,input [PIXEL_SIZE-1:0] Pix_608,input [PIXEL_SIZE-1:0] Pix_609,input [PIXEL_SIZE-1:0] Pix_610,input [PIXEL_SIZE-1:0] Pix_611,input [PIXEL_SIZE-1:0] Pix_612,input [PIXEL_SIZE-1:0] Pix_613,input [PIXEL_SIZE-1:0] Pix_614,input [PIXEL_SIZE-1:0] Pix_615,input [PIXEL_SIZE-1:0] Pix_616,input [PIXEL_SIZE-1:0] Pix_617,input [PIXEL_SIZE-1:0] Pix_618,input [PIXEL_SIZE-1:0] Pix_619,input [PIXEL_SIZE-1:0] Pix_620,input [PIXEL_SIZE-1:0] Pix_621,input [PIXEL_SIZE-1:0] Pix_622,input [PIXEL_SIZE-1:0] Pix_623,input [PIXEL_SIZE-1:0] Pix_624,input [PIXEL_SIZE-1:0] Pix_625,input [PIXEL_SIZE-1:0] Pix_626,input [PIXEL_SIZE-1:0] Pix_627,input [PIXEL_SIZE-1:0] Pix_628,input [PIXEL_SIZE-1:0] Pix_629,input [PIXEL_SIZE-1:0] Pix_630,input [PIXEL_SIZE-1:0] Pix_631,input [PIXEL_SIZE-1:0] Pix_632,input [PIXEL_SIZE-1:0] Pix_633,input [PIXEL_SIZE-1:0] Pix_634,input [PIXEL_SIZE-1:0] Pix_635,input [PIXEL_SIZE-1:0] Pix_636,input [PIXEL_SIZE-1:0] Pix_637,input [PIXEL_SIZE-1:0] Pix_638,input [PIXEL_SIZE-1:0] Pix_639,input [PIXEL_SIZE-1:0] Pix_640,input [PIXEL_SIZE-1:0] Pix_641,input [PIXEL_SIZE-1:0] Pix_642,input [PIXEL_SIZE-1:0] Pix_643,input [PIXEL_SIZE-1:0] Pix_644,input [PIXEL_SIZE-1:0] Pix_645,input [PIXEL_SIZE-1:0] Pix_646,input [PIXEL_SIZE-1:0] Pix_647,input [PIXEL_SIZE-1:0] Pix_648,input [PIXEL_SIZE-1:0] Pix_649,input [PIXEL_SIZE-1:0] Pix_650,input [PIXEL_SIZE-1:0] Pix_651,input [PIXEL_SIZE-1:0] Pix_652,input [PIXEL_SIZE-1:0] Pix_653,input [PIXEL_SIZE-1:0] Pix_654,input [PIXEL_SIZE-1:0] Pix_655,input [PIXEL_SIZE-1:0] Pix_656,input [PIXEL_SIZE-1:0] Pix_657,input [PIXEL_SIZE-1:0] Pix_658,input [PIXEL_SIZE-1:0] Pix_659,input [PIXEL_SIZE-1:0] Pix_660,input [PIXEL_SIZE-1:0] Pix_661,input [PIXEL_SIZE-1:0] Pix_662,input [PIXEL_SIZE-1:0] Pix_663,input [PIXEL_SIZE-1:0] Pix_664,input [PIXEL_SIZE-1:0] Pix_665,input [PIXEL_SIZE-1:0] Pix_666,input [PIXEL_SIZE-1:0] Pix_667,input [PIXEL_SIZE-1:0] Pix_668,input [PIXEL_SIZE-1:0] Pix_669,input [PIXEL_SIZE-1:0] Pix_670,input [PIXEL_SIZE-1:0] Pix_671,input [PIXEL_SIZE-1:0] Pix_672,input [PIXEL_SIZE-1:0] Pix_673,input [PIXEL_SIZE-1:0] Pix_674,input [PIXEL_SIZE-1:0] Pix_675,input [PIXEL_SIZE-1:0] Pix_676,input [PIXEL_SIZE-1:0] Pix_677,input [PIXEL_SIZE-1:0] Pix_678,input [PIXEL_SIZE-1:0] Pix_679,input [PIXEL_SIZE-1:0] Pix_680,input [PIXEL_SIZE-1:0] Pix_681,input [PIXEL_SIZE-1:0] Pix_682,input [PIXEL_SIZE-1:0] Pix_683,input [PIXEL_SIZE-1:0] Pix_684,input [PIXEL_SIZE-1:0] Pix_685,input [PIXEL_SIZE-1:0] Pix_686,input [PIXEL_SIZE-1:0] Pix_687,input [PIXEL_SIZE-1:0] Pix_688,input [PIXEL_SIZE-1:0] Pix_689,input [PIXEL_SIZE-1:0] Pix_690,input [PIXEL_SIZE-1:0] Pix_691,input [PIXEL_SIZE-1:0] Pix_692,input [PIXEL_SIZE-1:0] Pix_693,input [PIXEL_SIZE-1:0] Pix_694,input [PIXEL_SIZE-1:0] Pix_695,input [PIXEL_SIZE-1:0] Pix_696,input [PIXEL_SIZE-1:0] Pix_697,input [PIXEL_SIZE-1:0] Pix_698,input [PIXEL_SIZE-1:0] Pix_699,input [PIXEL_SIZE-1:0] Pix_700,input [PIXEL_SIZE-1:0] Pix_701,input [PIXEL_SIZE-1:0] Pix_702,input [PIXEL_SIZE-1:0] Pix_703,input [PIXEL_SIZE-1:0] Pix_704,input [PIXEL_SIZE-1:0] Pix_705,input [PIXEL_SIZE-1:0] Pix_706,input [PIXEL_SIZE-1:0] Pix_707,input [PIXEL_SIZE-1:0] Pix_708,input [PIXEL_SIZE-1:0] Pix_709,input [PIXEL_SIZE-1:0] Pix_710,input [PIXEL_SIZE-1:0] Pix_711,input [PIXEL_SIZE-1:0] Pix_712,input [PIXEL_SIZE-1:0] Pix_713,input [PIXEL_SIZE-1:0] Pix_714,input [PIXEL_SIZE-1:0] Pix_715,input [PIXEL_SIZE-1:0] Pix_716,input [PIXEL_SIZE-1:0] Pix_717,input [PIXEL_SIZE-1:0] Pix_718,input [PIXEL_SIZE-1:0] Pix_719,input [PIXEL_SIZE-1:0] Pix_720,input [PIXEL_SIZE-1:0] Pix_721,input [PIXEL_SIZE-1:0] Pix_722,input [PIXEL_SIZE-1:0] Pix_723,input [PIXEL_SIZE-1:0] Pix_724,input [PIXEL_SIZE-1:0] Pix_725,input [PIXEL_SIZE-1:0] Pix_726,input [PIXEL_SIZE-1:0] Pix_727,input [PIXEL_SIZE-1:0] Pix_728,input [PIXEL_SIZE-1:0] Pix_729,input [PIXEL_SIZE-1:0] Pix_730,input [PIXEL_SIZE-1:0] Pix_731,input [PIXEL_SIZE-1:0] Pix_732,input [PIXEL_SIZE-1:0] Pix_733,input [PIXEL_SIZE-1:0] Pix_734,input [PIXEL_SIZE-1:0] Pix_735,input [PIXEL_SIZE-1:0] Pix_736,input [PIXEL_SIZE-1:0] Pix_737,input [PIXEL_SIZE-1:0] Pix_738,input [PIXEL_SIZE-1:0] Pix_739,input [PIXEL_SIZE-1:0] Pix_740,input [PIXEL_SIZE-1:0] Pix_741,input [PIXEL_SIZE-1:0] Pix_742,input [PIXEL_SIZE-1:0] Pix_743,input [PIXEL_SIZE-1:0] Pix_744,input [PIXEL_SIZE-1:0] Pix_745,input [PIXEL_SIZE-1:0] Pix_746,input [PIXEL_SIZE-1:0] Pix_747,input [PIXEL_SIZE-1:0] Pix_748,input [PIXEL_SIZE-1:0] Pix_749,input [PIXEL_SIZE-1:0] Pix_750,input [PIXEL_SIZE-1:0] Pix_751,input [PIXEL_SIZE-1:0] Pix_752,input [PIXEL_SIZE-1:0] Pix_753,input [PIXEL_SIZE-1:0] Pix_754,input [PIXEL_SIZE-1:0] Pix_755,input [PIXEL_SIZE-1:0] Pix_756,input [PIXEL_SIZE-1:0] Pix_757,input [PIXEL_SIZE-1:0] Pix_758,input [PIXEL_SIZE-1:0] Pix_759,input [PIXEL_SIZE-1:0] Pix_760,input [PIXEL_SIZE-1:0] Pix_761,input [PIXEL_SIZE-1:0] Pix_762,input [PIXEL_SIZE-1:0] Pix_763,input [PIXEL_SIZE-1:0] Pix_764,input [PIXEL_SIZE-1:0] Pix_765,input [PIXEL_SIZE-1:0] Pix_766,input [PIXEL_SIZE-1:0] Pix_767,input [PIXEL_SIZE-1:0] Pix_768,input [PIXEL_SIZE-1:0] Pix_769,input [PIXEL_SIZE-1:0] Pix_770,input [PIXEL_SIZE-1:0] Pix_771,input [PIXEL_SIZE-1:0] Pix_772,input [PIXEL_SIZE-1:0] Pix_773,input [PIXEL_SIZE-1:0] Pix_774,input [PIXEL_SIZE-1:0] Pix_775,input [PIXEL_SIZE-1:0] Pix_776,input [PIXEL_SIZE-1:0] Pix_777,input [PIXEL_SIZE-1:0] Pix_778,input [PIXEL_SIZE-1:0] Pix_779,input [PIXEL_SIZE-1:0] Pix_780,input [PIXEL_SIZE-1:0] Pix_781,input [PIXEL_SIZE-1:0] Pix_782,input [PIXEL_SIZE-1:0] Pix_783,input [PIXEL_SIZE-1:0] Pix_784,
output [3:0] Image_Number,
output Output_Valid
);

reg[PIXEL_SIZE-1:0] PixelsStore[0:PIXEL_N-1];
reg[WEIGHT_SIZE-1:0] WeightsStore[0:PIXEL_N-1][0:NEURONS-1];
reg[31:0] switchCounter;
reg ready;
reg internalReset;
wire[VAL_SIZE*NEURONS-1:0] value;

assign Output_Valid = ready;

always@(posedge clk)begin
	if(GlobalReset == 1'b0)begin
		switchCounter <= 0;
		ready = 1'b0;
		internalReset = 1'b0;
		PixelsStore[0]<=0;PixelsStore[1]<=0;PixelsStore[2]<=0;PixelsStore[3]<=0;PixelsStore[4]<=0;PixelsStore[5]<=0;PixelsStore[6]<=0;PixelsStore[7]<=0;PixelsStore[8]<=0;PixelsStore[9]<=0;PixelsStore[10]<=0;PixelsStore[11]<=0;PixelsStore[12]<=0;PixelsStore[13]<=0;PixelsStore[14]<=0;PixelsStore[15]<=0;PixelsStore[16]<=0;PixelsStore[17]<=0;PixelsStore[18]<=0;PixelsStore[19]<=0;PixelsStore[20]<=0;PixelsStore[21]<=0;PixelsStore[22]<=0;PixelsStore[23]<=0;PixelsStore[24]<=0;PixelsStore[25]<=0;PixelsStore[26]<=0;PixelsStore[27]<=0;PixelsStore[28]<=0;PixelsStore[29]<=0;PixelsStore[30]<=0;PixelsStore[31]<=0;PixelsStore[32]<=0;PixelsStore[33]<=0;PixelsStore[34]<=0;PixelsStore[35]<=0;PixelsStore[36]<=0;PixelsStore[37]<=0;PixelsStore[38]<=0;PixelsStore[39]<=0;PixelsStore[40]<=0;PixelsStore[41]<=0;PixelsStore[42]<=0;PixelsStore[43]<=0;PixelsStore[44]<=0;PixelsStore[45]<=0;PixelsStore[46]<=0;PixelsStore[47]<=0;PixelsStore[48]<=0;PixelsStore[49]<=0;PixelsStore[50]<=0;PixelsStore[51]<=0;PixelsStore[52]<=0;PixelsStore[53]<=0;PixelsStore[54]<=0;PixelsStore[55]<=0;PixelsStore[56]<=0;PixelsStore[57]<=0;PixelsStore[58]<=0;PixelsStore[59]<=0;PixelsStore[60]<=0;PixelsStore[61]<=0;PixelsStore[62]<=0;PixelsStore[63]<=0;PixelsStore[64]<=0;PixelsStore[65]<=0;PixelsStore[66]<=0;PixelsStore[67]<=0;PixelsStore[68]<=0;PixelsStore[69]<=0;PixelsStore[70]<=0;PixelsStore[71]<=0;PixelsStore[72]<=0;PixelsStore[73]<=0;PixelsStore[74]<=0;PixelsStore[75]<=0;PixelsStore[76]<=0;PixelsStore[77]<=0;PixelsStore[78]<=0;PixelsStore[79]<=0;PixelsStore[80]<=0;PixelsStore[81]<=0;PixelsStore[82]<=0;PixelsStore[83]<=0;PixelsStore[84]<=0;PixelsStore[85]<=0;PixelsStore[86]<=0;PixelsStore[87]<=0;PixelsStore[88]<=0;PixelsStore[89]<=0;PixelsStore[90]<=0;PixelsStore[91]<=0;PixelsStore[92]<=0;PixelsStore[93]<=0;PixelsStore[94]<=0;PixelsStore[95]<=0;PixelsStore[96]<=0;PixelsStore[97]<=0;PixelsStore[98]<=0;PixelsStore[99]<=0;PixelsStore[100]<=0;PixelsStore[101]<=0;PixelsStore[102]<=0;PixelsStore[103]<=0;PixelsStore[104]<=0;PixelsStore[105]<=0;PixelsStore[106]<=0;PixelsStore[107]<=0;PixelsStore[108]<=0;PixelsStore[109]<=0;PixelsStore[110]<=0;PixelsStore[111]<=0;PixelsStore[112]<=0;PixelsStore[113]<=0;PixelsStore[114]<=0;PixelsStore[115]<=0;PixelsStore[116]<=0;PixelsStore[117]<=0;PixelsStore[118]<=0;PixelsStore[119]<=0;PixelsStore[120]<=0;PixelsStore[121]<=0;PixelsStore[122]<=0;PixelsStore[123]<=0;PixelsStore[124]<=0;PixelsStore[125]<=0;PixelsStore[126]<=0;PixelsStore[127]<=0;PixelsStore[128]<=0;PixelsStore[129]<=0;PixelsStore[130]<=0;PixelsStore[131]<=0;PixelsStore[132]<=0;PixelsStore[133]<=0;PixelsStore[134]<=0;PixelsStore[135]<=0;PixelsStore[136]<=0;PixelsStore[137]<=0;PixelsStore[138]<=0;PixelsStore[139]<=0;PixelsStore[140]<=0;PixelsStore[141]<=0;PixelsStore[142]<=0;PixelsStore[143]<=0;PixelsStore[144]<=0;PixelsStore[145]<=0;PixelsStore[146]<=0;PixelsStore[147]<=0;PixelsStore[148]<=0;PixelsStore[149]<=0;PixelsStore[150]<=0;PixelsStore[151]<=0;PixelsStore[152]<=0;PixelsStore[153]<=0;PixelsStore[154]<=0;PixelsStore[155]<=0;PixelsStore[156]<=0;PixelsStore[157]<=0;PixelsStore[158]<=0;PixelsStore[159]<=0;PixelsStore[160]<=0;PixelsStore[161]<=0;PixelsStore[162]<=0;PixelsStore[163]<=0;PixelsStore[164]<=0;PixelsStore[165]<=0;PixelsStore[166]<=0;PixelsStore[167]<=0;PixelsStore[168]<=0;PixelsStore[169]<=0;PixelsStore[170]<=0;PixelsStore[171]<=0;PixelsStore[172]<=0;PixelsStore[173]<=0;PixelsStore[174]<=0;PixelsStore[175]<=0;PixelsStore[176]<=0;PixelsStore[177]<=0;PixelsStore[178]<=0;PixelsStore[179]<=0;PixelsStore[180]<=0;PixelsStore[181]<=0;PixelsStore[182]<=0;PixelsStore[183]<=0;PixelsStore[184]<=0;PixelsStore[185]<=0;PixelsStore[186]<=0;PixelsStore[187]<=0;PixelsStore[188]<=0;PixelsStore[189]<=0;PixelsStore[190]<=0;PixelsStore[191]<=0;PixelsStore[192]<=0;PixelsStore[193]<=0;PixelsStore[194]<=0;PixelsStore[195]<=0;PixelsStore[196]<=0;PixelsStore[197]<=0;PixelsStore[198]<=0;PixelsStore[199]<=0;PixelsStore[200]<=0;PixelsStore[201]<=0;PixelsStore[202]<=0;PixelsStore[203]<=0;PixelsStore[204]<=0;PixelsStore[205]<=0;PixelsStore[206]<=0;PixelsStore[207]<=0;PixelsStore[208]<=0;PixelsStore[209]<=0;PixelsStore[210]<=0;PixelsStore[211]<=0;PixelsStore[212]<=0;PixelsStore[213]<=0;PixelsStore[214]<=0;PixelsStore[215]<=0;PixelsStore[216]<=0;PixelsStore[217]<=0;PixelsStore[218]<=0;PixelsStore[219]<=0;PixelsStore[220]<=0;PixelsStore[221]<=0;PixelsStore[222]<=0;PixelsStore[223]<=0;PixelsStore[224]<=0;PixelsStore[225]<=0;PixelsStore[226]<=0;PixelsStore[227]<=0;PixelsStore[228]<=0;PixelsStore[229]<=0;PixelsStore[230]<=0;PixelsStore[231]<=0;PixelsStore[232]<=0;PixelsStore[233]<=0;PixelsStore[234]<=0;PixelsStore[235]<=0;PixelsStore[236]<=0;PixelsStore[237]<=0;PixelsStore[238]<=0;PixelsStore[239]<=0;PixelsStore[240]<=0;PixelsStore[241]<=0;PixelsStore[242]<=0;PixelsStore[243]<=0;PixelsStore[244]<=0;PixelsStore[245]<=0;PixelsStore[246]<=0;PixelsStore[247]<=0;PixelsStore[248]<=0;PixelsStore[249]<=0;PixelsStore[250]<=0;PixelsStore[251]<=0;PixelsStore[252]<=0;PixelsStore[253]<=0;PixelsStore[254]<=0;PixelsStore[255]<=0;PixelsStore[256]<=0;PixelsStore[257]<=0;PixelsStore[258]<=0;PixelsStore[259]<=0;PixelsStore[260]<=0;PixelsStore[261]<=0;PixelsStore[262]<=0;PixelsStore[263]<=0;PixelsStore[264]<=0;PixelsStore[265]<=0;PixelsStore[266]<=0;PixelsStore[267]<=0;PixelsStore[268]<=0;PixelsStore[269]<=0;PixelsStore[270]<=0;PixelsStore[271]<=0;PixelsStore[272]<=0;PixelsStore[273]<=0;PixelsStore[274]<=0;PixelsStore[275]<=0;PixelsStore[276]<=0;PixelsStore[277]<=0;PixelsStore[278]<=0;PixelsStore[279]<=0;PixelsStore[280]<=0;PixelsStore[281]<=0;PixelsStore[282]<=0;PixelsStore[283]<=0;PixelsStore[284]<=0;PixelsStore[285]<=0;PixelsStore[286]<=0;PixelsStore[287]<=0;PixelsStore[288]<=0;PixelsStore[289]<=0;PixelsStore[290]<=0;PixelsStore[291]<=0;PixelsStore[292]<=0;PixelsStore[293]<=0;PixelsStore[294]<=0;PixelsStore[295]<=0;PixelsStore[296]<=0;PixelsStore[297]<=0;PixelsStore[298]<=0;PixelsStore[299]<=0;PixelsStore[300]<=0;PixelsStore[301]<=0;PixelsStore[302]<=0;PixelsStore[303]<=0;PixelsStore[304]<=0;PixelsStore[305]<=0;PixelsStore[306]<=0;PixelsStore[307]<=0;PixelsStore[308]<=0;PixelsStore[309]<=0;PixelsStore[310]<=0;PixelsStore[311]<=0;PixelsStore[312]<=0;PixelsStore[313]<=0;PixelsStore[314]<=0;PixelsStore[315]<=0;PixelsStore[316]<=0;PixelsStore[317]<=0;PixelsStore[318]<=0;PixelsStore[319]<=0;PixelsStore[320]<=0;PixelsStore[321]<=0;PixelsStore[322]<=0;PixelsStore[323]<=0;PixelsStore[324]<=0;PixelsStore[325]<=0;PixelsStore[326]<=0;PixelsStore[327]<=0;PixelsStore[328]<=0;PixelsStore[329]<=0;PixelsStore[330]<=0;PixelsStore[331]<=0;PixelsStore[332]<=0;PixelsStore[333]<=0;PixelsStore[334]<=0;PixelsStore[335]<=0;PixelsStore[336]<=0;PixelsStore[337]<=0;PixelsStore[338]<=0;PixelsStore[339]<=0;PixelsStore[340]<=0;PixelsStore[341]<=0;PixelsStore[342]<=0;PixelsStore[343]<=0;PixelsStore[344]<=0;PixelsStore[345]<=0;PixelsStore[346]<=0;PixelsStore[347]<=0;PixelsStore[348]<=0;PixelsStore[349]<=0;PixelsStore[350]<=0;PixelsStore[351]<=0;PixelsStore[352]<=0;PixelsStore[353]<=0;PixelsStore[354]<=0;PixelsStore[355]<=0;PixelsStore[356]<=0;PixelsStore[357]<=0;PixelsStore[358]<=0;PixelsStore[359]<=0;PixelsStore[360]<=0;PixelsStore[361]<=0;PixelsStore[362]<=0;PixelsStore[363]<=0;PixelsStore[364]<=0;PixelsStore[365]<=0;PixelsStore[366]<=0;PixelsStore[367]<=0;PixelsStore[368]<=0;PixelsStore[369]<=0;PixelsStore[370]<=0;PixelsStore[371]<=0;PixelsStore[372]<=0;PixelsStore[373]<=0;PixelsStore[374]<=0;PixelsStore[375]<=0;PixelsStore[376]<=0;PixelsStore[377]<=0;PixelsStore[378]<=0;PixelsStore[379]<=0;PixelsStore[380]<=0;PixelsStore[381]<=0;PixelsStore[382]<=0;PixelsStore[383]<=0;PixelsStore[384]<=0;PixelsStore[385]<=0;PixelsStore[386]<=0;PixelsStore[387]<=0;PixelsStore[388]<=0;PixelsStore[389]<=0;PixelsStore[390]<=0;PixelsStore[391]<=0;PixelsStore[392]<=0;PixelsStore[393]<=0;PixelsStore[394]<=0;PixelsStore[395]<=0;PixelsStore[396]<=0;PixelsStore[397]<=0;PixelsStore[398]<=0;PixelsStore[399]<=0;PixelsStore[400]<=0;PixelsStore[401]<=0;PixelsStore[402]<=0;PixelsStore[403]<=0;PixelsStore[404]<=0;PixelsStore[405]<=0;PixelsStore[406]<=0;PixelsStore[407]<=0;PixelsStore[408]<=0;PixelsStore[409]<=0;PixelsStore[410]<=0;PixelsStore[411]<=0;PixelsStore[412]<=0;PixelsStore[413]<=0;PixelsStore[414]<=0;PixelsStore[415]<=0;PixelsStore[416]<=0;PixelsStore[417]<=0;PixelsStore[418]<=0;PixelsStore[419]<=0;PixelsStore[420]<=0;PixelsStore[421]<=0;PixelsStore[422]<=0;PixelsStore[423]<=0;PixelsStore[424]<=0;PixelsStore[425]<=0;PixelsStore[426]<=0;PixelsStore[427]<=0;PixelsStore[428]<=0;PixelsStore[429]<=0;PixelsStore[430]<=0;PixelsStore[431]<=0;PixelsStore[432]<=0;PixelsStore[433]<=0;PixelsStore[434]<=0;PixelsStore[435]<=0;PixelsStore[436]<=0;PixelsStore[437]<=0;PixelsStore[438]<=0;PixelsStore[439]<=0;PixelsStore[440]<=0;PixelsStore[441]<=0;PixelsStore[442]<=0;PixelsStore[443]<=0;PixelsStore[444]<=0;PixelsStore[445]<=0;PixelsStore[446]<=0;PixelsStore[447]<=0;PixelsStore[448]<=0;PixelsStore[449]<=0;PixelsStore[450]<=0;PixelsStore[451]<=0;PixelsStore[452]<=0;PixelsStore[453]<=0;PixelsStore[454]<=0;PixelsStore[455]<=0;PixelsStore[456]<=0;PixelsStore[457]<=0;PixelsStore[458]<=0;PixelsStore[459]<=0;PixelsStore[460]<=0;PixelsStore[461]<=0;PixelsStore[462]<=0;PixelsStore[463]<=0;PixelsStore[464]<=0;PixelsStore[465]<=0;PixelsStore[466]<=0;PixelsStore[467]<=0;PixelsStore[468]<=0;PixelsStore[469]<=0;PixelsStore[470]<=0;PixelsStore[471]<=0;PixelsStore[472]<=0;PixelsStore[473]<=0;PixelsStore[474]<=0;PixelsStore[475]<=0;PixelsStore[476]<=0;PixelsStore[477]<=0;PixelsStore[478]<=0;PixelsStore[479]<=0;PixelsStore[480]<=0;PixelsStore[481]<=0;PixelsStore[482]<=0;PixelsStore[483]<=0;PixelsStore[484]<=0;PixelsStore[485]<=0;PixelsStore[486]<=0;PixelsStore[487]<=0;PixelsStore[488]<=0;PixelsStore[489]<=0;PixelsStore[490]<=0;PixelsStore[491]<=0;PixelsStore[492]<=0;PixelsStore[493]<=0;PixelsStore[494]<=0;PixelsStore[495]<=0;PixelsStore[496]<=0;PixelsStore[497]<=0;PixelsStore[498]<=0;PixelsStore[499]<=0;PixelsStore[500]<=0;PixelsStore[501]<=0;PixelsStore[502]<=0;PixelsStore[503]<=0;PixelsStore[504]<=0;PixelsStore[505]<=0;PixelsStore[506]<=0;PixelsStore[507]<=0;PixelsStore[508]<=0;PixelsStore[509]<=0;PixelsStore[510]<=0;PixelsStore[511]<=0;PixelsStore[512]<=0;PixelsStore[513]<=0;PixelsStore[514]<=0;PixelsStore[515]<=0;PixelsStore[516]<=0;PixelsStore[517]<=0;PixelsStore[518]<=0;PixelsStore[519]<=0;PixelsStore[520]<=0;PixelsStore[521]<=0;PixelsStore[522]<=0;PixelsStore[523]<=0;PixelsStore[524]<=0;PixelsStore[525]<=0;PixelsStore[526]<=0;PixelsStore[527]<=0;PixelsStore[528]<=0;PixelsStore[529]<=0;PixelsStore[530]<=0;PixelsStore[531]<=0;PixelsStore[532]<=0;PixelsStore[533]<=0;PixelsStore[534]<=0;PixelsStore[535]<=0;PixelsStore[536]<=0;PixelsStore[537]<=0;PixelsStore[538]<=0;PixelsStore[539]<=0;PixelsStore[540]<=0;PixelsStore[541]<=0;PixelsStore[542]<=0;PixelsStore[543]<=0;PixelsStore[544]<=0;PixelsStore[545]<=0;PixelsStore[546]<=0;PixelsStore[547]<=0;PixelsStore[548]<=0;PixelsStore[549]<=0;PixelsStore[550]<=0;PixelsStore[551]<=0;PixelsStore[552]<=0;PixelsStore[553]<=0;PixelsStore[554]<=0;PixelsStore[555]<=0;PixelsStore[556]<=0;PixelsStore[557]<=0;PixelsStore[558]<=0;PixelsStore[559]<=0;PixelsStore[560]<=0;PixelsStore[561]<=0;PixelsStore[562]<=0;PixelsStore[563]<=0;PixelsStore[564]<=0;PixelsStore[565]<=0;PixelsStore[566]<=0;PixelsStore[567]<=0;PixelsStore[568]<=0;PixelsStore[569]<=0;PixelsStore[570]<=0;PixelsStore[571]<=0;PixelsStore[572]<=0;PixelsStore[573]<=0;PixelsStore[574]<=0;PixelsStore[575]<=0;PixelsStore[576]<=0;PixelsStore[577]<=0;PixelsStore[578]<=0;PixelsStore[579]<=0;PixelsStore[580]<=0;PixelsStore[581]<=0;PixelsStore[582]<=0;PixelsStore[583]<=0;PixelsStore[584]<=0;PixelsStore[585]<=0;PixelsStore[586]<=0;PixelsStore[587]<=0;PixelsStore[588]<=0;PixelsStore[589]<=0;PixelsStore[590]<=0;PixelsStore[591]<=0;PixelsStore[592]<=0;PixelsStore[593]<=0;PixelsStore[594]<=0;PixelsStore[595]<=0;PixelsStore[596]<=0;PixelsStore[597]<=0;PixelsStore[598]<=0;PixelsStore[599]<=0;PixelsStore[600]<=0;PixelsStore[601]<=0;PixelsStore[602]<=0;PixelsStore[603]<=0;PixelsStore[604]<=0;PixelsStore[605]<=0;PixelsStore[606]<=0;PixelsStore[607]<=0;PixelsStore[608]<=0;PixelsStore[609]<=0;PixelsStore[610]<=0;PixelsStore[611]<=0;PixelsStore[612]<=0;PixelsStore[613]<=0;PixelsStore[614]<=0;PixelsStore[615]<=0;PixelsStore[616]<=0;PixelsStore[617]<=0;PixelsStore[618]<=0;PixelsStore[619]<=0;PixelsStore[620]<=0;PixelsStore[621]<=0;PixelsStore[622]<=0;PixelsStore[623]<=0;PixelsStore[624]<=0;PixelsStore[625]<=0;PixelsStore[626]<=0;PixelsStore[627]<=0;PixelsStore[628]<=0;PixelsStore[629]<=0;PixelsStore[630]<=0;PixelsStore[631]<=0;PixelsStore[632]<=0;PixelsStore[633]<=0;PixelsStore[634]<=0;PixelsStore[635]<=0;PixelsStore[636]<=0;PixelsStore[637]<=0;PixelsStore[638]<=0;PixelsStore[639]<=0;PixelsStore[640]<=0;PixelsStore[641]<=0;PixelsStore[642]<=0;PixelsStore[643]<=0;PixelsStore[644]<=0;PixelsStore[645]<=0;PixelsStore[646]<=0;PixelsStore[647]<=0;PixelsStore[648]<=0;PixelsStore[649]<=0;PixelsStore[650]<=0;PixelsStore[651]<=0;PixelsStore[652]<=0;PixelsStore[653]<=0;PixelsStore[654]<=0;PixelsStore[655]<=0;PixelsStore[656]<=0;PixelsStore[657]<=0;PixelsStore[658]<=0;PixelsStore[659]<=0;PixelsStore[660]<=0;PixelsStore[661]<=0;PixelsStore[662]<=0;PixelsStore[663]<=0;PixelsStore[664]<=0;PixelsStore[665]<=0;PixelsStore[666]<=0;PixelsStore[667]<=0;PixelsStore[668]<=0;PixelsStore[669]<=0;PixelsStore[670]<=0;PixelsStore[671]<=0;PixelsStore[672]<=0;PixelsStore[673]<=0;PixelsStore[674]<=0;PixelsStore[675]<=0;PixelsStore[676]<=0;PixelsStore[677]<=0;PixelsStore[678]<=0;PixelsStore[679]<=0;PixelsStore[680]<=0;PixelsStore[681]<=0;PixelsStore[682]<=0;PixelsStore[683]<=0;PixelsStore[684]<=0;PixelsStore[685]<=0;PixelsStore[686]<=0;PixelsStore[687]<=0;PixelsStore[688]<=0;PixelsStore[689]<=0;PixelsStore[690]<=0;PixelsStore[691]<=0;PixelsStore[692]<=0;PixelsStore[693]<=0;PixelsStore[694]<=0;PixelsStore[695]<=0;PixelsStore[696]<=0;PixelsStore[697]<=0;PixelsStore[698]<=0;PixelsStore[699]<=0;PixelsStore[700]<=0;PixelsStore[701]<=0;PixelsStore[702]<=0;PixelsStore[703]<=0;PixelsStore[704]<=0;PixelsStore[705]<=0;PixelsStore[706]<=0;PixelsStore[707]<=0;PixelsStore[708]<=0;PixelsStore[709]<=0;PixelsStore[710]<=0;PixelsStore[711]<=0;PixelsStore[712]<=0;PixelsStore[713]<=0;PixelsStore[714]<=0;PixelsStore[715]<=0;PixelsStore[716]<=0;PixelsStore[717]<=0;PixelsStore[718]<=0;PixelsStore[719]<=0;PixelsStore[720]<=0;PixelsStore[721]<=0;PixelsStore[722]<=0;PixelsStore[723]<=0;PixelsStore[724]<=0;PixelsStore[725]<=0;PixelsStore[726]<=0;PixelsStore[727]<=0;PixelsStore[728]<=0;PixelsStore[729]<=0;PixelsStore[730]<=0;PixelsStore[731]<=0;PixelsStore[732]<=0;PixelsStore[733]<=0;PixelsStore[734]<=0;PixelsStore[735]<=0;PixelsStore[736]<=0;PixelsStore[737]<=0;PixelsStore[738]<=0;PixelsStore[739]<=0;PixelsStore[740]<=0;PixelsStore[741]<=0;PixelsStore[742]<=0;PixelsStore[743]<=0;PixelsStore[744]<=0;PixelsStore[745]<=0;PixelsStore[746]<=0;PixelsStore[747]<=0;PixelsStore[748]<=0;PixelsStore[749]<=0;PixelsStore[750]<=0;PixelsStore[751]<=0;PixelsStore[752]<=0;PixelsStore[753]<=0;PixelsStore[754]<=0;PixelsStore[755]<=0;PixelsStore[756]<=0;PixelsStore[757]<=0;PixelsStore[758]<=0;PixelsStore[759]<=0;PixelsStore[760]<=0;PixelsStore[761]<=0;PixelsStore[762]<=0;PixelsStore[763]<=0;PixelsStore[764]<=0;PixelsStore[765]<=0;PixelsStore[766]<=0;PixelsStore[767]<=0;PixelsStore[768]<=0;PixelsStore[769]<=0;PixelsStore[770]<=0;PixelsStore[771]<=0;PixelsStore[772]<=0;PixelsStore[773]<=0;PixelsStore[774]<=0;PixelsStore[775]<=0;PixelsStore[776]<=0;PixelsStore[777]<=0;PixelsStore[778]<=0;PixelsStore[779]<=0;PixelsStore[780]<=0;PixelsStore[781]<=0;PixelsStore[782]<=0;PixelsStore[783]<=0;PixelsStore[784]<=0;
		WeightsStore[0][0]<=0;WeightsStore[0][1]<=0;WeightsStore[0][2]<=0;WeightsStore[0][3]<=0;WeightsStore[0][4]<=0;WeightsStore[0][5]<=0;WeightsStore[0][6]<=0;WeightsStore[0][7]<=0;WeightsStore[0][8]<=0;WeightsStore[0][9]<=0;WeightsStore[0][10]<=0;WeightsStore[0][11]<=0;WeightsStore[0][12]<=0;WeightsStore[0][13]<=0;WeightsStore[0][14]<=0;WeightsStore[0][15]<=0;WeightsStore[0][16]<=0;WeightsStore[0][17]<=0;WeightsStore[0][18]<=0;WeightsStore[0][19]<=0;WeightsStore[0][20]<=0;WeightsStore[0][21]<=0;WeightsStore[0][22]<=0;WeightsStore[0][23]<=0;WeightsStore[0][24]<=0;WeightsStore[0][25]<=0;WeightsStore[0][26]<=0;WeightsStore[0][27]<=0;WeightsStore[0][28]<=0;WeightsStore[0][29]<=0;WeightsStore[0][30]<=0;WeightsStore[0][31]<=0;WeightsStore[0][32]<=0;WeightsStore[0][33]<=0;WeightsStore[0][34]<=0;WeightsStore[0][35]<=0;WeightsStore[0][36]<=0;WeightsStore[0][37]<=0;WeightsStore[0][38]<=0;WeightsStore[0][39]<=0;WeightsStore[0][40]<=0;WeightsStore[0][41]<=0;WeightsStore[0][42]<=0;WeightsStore[0][43]<=0;WeightsStore[0][44]<=0;WeightsStore[0][45]<=0;WeightsStore[0][46]<=0;WeightsStore[0][47]<=0;WeightsStore[0][48]<=0;WeightsStore[0][49]<=0;WeightsStore[0][50]<=0;WeightsStore[0][51]<=0;WeightsStore[0][52]<=0;WeightsStore[0][53]<=0;WeightsStore[0][54]<=0;WeightsStore[0][55]<=0;WeightsStore[0][56]<=0;WeightsStore[0][57]<=0;WeightsStore[0][58]<=0;WeightsStore[0][59]<=0;WeightsStore[0][60]<=0;WeightsStore[0][61]<=0;WeightsStore[0][62]<=0;WeightsStore[0][63]<=0;WeightsStore[0][64]<=0;WeightsStore[0][65]<=0;WeightsStore[0][66]<=0;WeightsStore[0][67]<=0;WeightsStore[0][68]<=0;WeightsStore[0][69]<=0;WeightsStore[0][70]<=0;WeightsStore[0][71]<=0;WeightsStore[0][72]<=0;WeightsStore[0][73]<=0;WeightsStore[0][74]<=0;WeightsStore[0][75]<=0;WeightsStore[0][76]<=0;WeightsStore[0][77]<=0;WeightsStore[0][78]<=0;WeightsStore[0][79]<=0;WeightsStore[0][80]<=0;WeightsStore[0][81]<=0;WeightsStore[0][82]<=0;WeightsStore[0][83]<=0;WeightsStore[0][84]<=0;WeightsStore[0][85]<=0;WeightsStore[0][86]<=0;WeightsStore[0][87]<=0;WeightsStore[0][88]<=0;WeightsStore[0][89]<=0;WeightsStore[0][90]<=0;WeightsStore[0][91]<=0;WeightsStore[0][92]<=0;WeightsStore[0][93]<=0;WeightsStore[0][94]<=0;WeightsStore[0][95]<=0;WeightsStore[0][96]<=0;WeightsStore[0][97]<=0;WeightsStore[0][98]<=0;WeightsStore[0][99]<=0;WeightsStore[0][100]<=0;WeightsStore[0][101]<=0;WeightsStore[0][102]<=0;WeightsStore[0][103]<=0;WeightsStore[0][104]<=0;WeightsStore[0][105]<=0;WeightsStore[0][106]<=0;WeightsStore[0][107]<=0;WeightsStore[0][108]<=0;WeightsStore[0][109]<=0;WeightsStore[0][110]<=0;WeightsStore[0][111]<=0;WeightsStore[0][112]<=0;WeightsStore[0][113]<=0;WeightsStore[0][114]<=0;WeightsStore[0][115]<=0;WeightsStore[0][116]<=0;WeightsStore[0][117]<=0;WeightsStore[0][118]<=0;WeightsStore[0][119]<=0;WeightsStore[0][120]<=0;WeightsStore[0][121]<=0;WeightsStore[0][122]<=0;WeightsStore[0][123]<=0;WeightsStore[0][124]<=0;WeightsStore[0][125]<=0;WeightsStore[0][126]<=0;WeightsStore[0][127]<=0;WeightsStore[0][128]<=0;WeightsStore[0][129]<=0;WeightsStore[0][130]<=0;WeightsStore[0][131]<=0;WeightsStore[0][132]<=0;WeightsStore[0][133]<=0;WeightsStore[0][134]<=0;WeightsStore[0][135]<=0;WeightsStore[0][136]<=0;WeightsStore[0][137]<=0;WeightsStore[0][138]<=0;WeightsStore[0][139]<=0;WeightsStore[0][140]<=0;WeightsStore[0][141]<=0;WeightsStore[0][142]<=0;WeightsStore[0][143]<=0;WeightsStore[0][144]<=0;WeightsStore[0][145]<=0;WeightsStore[0][146]<=0;WeightsStore[0][147]<=0;WeightsStore[0][148]<=0;WeightsStore[0][149]<=0;WeightsStore[0][150]<=0;WeightsStore[0][151]<=0;WeightsStore[0][152]<=0;WeightsStore[0][153]<=0;WeightsStore[0][154]<=0;WeightsStore[0][155]<=0;WeightsStore[0][156]<=0;WeightsStore[0][157]<=0;WeightsStore[0][158]<=0;WeightsStore[0][159]<=0;WeightsStore[0][160]<=0;WeightsStore[0][161]<=0;WeightsStore[0][162]<=0;WeightsStore[0][163]<=0;WeightsStore[0][164]<=0;WeightsStore[0][165]<=0;WeightsStore[0][166]<=0;WeightsStore[0][167]<=0;WeightsStore[0][168]<=0;WeightsStore[0][169]<=0;WeightsStore[0][170]<=0;WeightsStore[0][171]<=0;WeightsStore[0][172]<=0;WeightsStore[0][173]<=0;WeightsStore[0][174]<=0;WeightsStore[0][175]<=0;WeightsStore[0][176]<=0;WeightsStore[0][177]<=0;WeightsStore[0][178]<=0;WeightsStore[0][179]<=0;WeightsStore[0][180]<=0;WeightsStore[0][181]<=0;WeightsStore[0][182]<=0;WeightsStore[0][183]<=0;WeightsStore[0][184]<=0;WeightsStore[0][185]<=0;WeightsStore[0][186]<=0;WeightsStore[0][187]<=0;WeightsStore[0][188]<=0;WeightsStore[0][189]<=0;WeightsStore[0][190]<=0;WeightsStore[0][191]<=0;WeightsStore[0][192]<=0;WeightsStore[0][193]<=0;WeightsStore[0][194]<=0;WeightsStore[0][195]<=0;WeightsStore[0][196]<=0;WeightsStore[0][197]<=0;WeightsStore[0][198]<=0;WeightsStore[0][199]<=0;WeightsStore[0][200]<=0;WeightsStore[0][201]<=0;WeightsStore[0][202]<=0;WeightsStore[0][203]<=0;WeightsStore[0][204]<=0;WeightsStore[0][205]<=0;WeightsStore[0][206]<=0;WeightsStore[0][207]<=0;WeightsStore[0][208]<=0;WeightsStore[0][209]<=0;WeightsStore[0][210]<=0;WeightsStore[0][211]<=0;WeightsStore[0][212]<=0;WeightsStore[0][213]<=0;WeightsStore[0][214]<=0;WeightsStore[0][215]<=0;WeightsStore[0][216]<=0;WeightsStore[0][217]<=0;WeightsStore[0][218]<=0;WeightsStore[0][219]<=0;WeightsStore[0][220]<=0;WeightsStore[0][221]<=0;WeightsStore[0][222]<=0;WeightsStore[0][223]<=0;WeightsStore[0][224]<=0;WeightsStore[0][225]<=0;WeightsStore[0][226]<=0;WeightsStore[0][227]<=0;WeightsStore[0][228]<=0;WeightsStore[0][229]<=0;WeightsStore[0][230]<=0;WeightsStore[0][231]<=0;WeightsStore[0][232]<=0;WeightsStore[0][233]<=0;WeightsStore[0][234]<=0;WeightsStore[0][235]<=0;WeightsStore[0][236]<=0;WeightsStore[0][237]<=0;WeightsStore[0][238]<=0;WeightsStore[0][239]<=0;WeightsStore[0][240]<=0;WeightsStore[0][241]<=0;WeightsStore[0][242]<=0;WeightsStore[0][243]<=0;WeightsStore[0][244]<=0;WeightsStore[0][245]<=0;WeightsStore[0][246]<=0;WeightsStore[0][247]<=0;WeightsStore[0][248]<=0;WeightsStore[0][249]<=0;WeightsStore[0][250]<=0;WeightsStore[0][251]<=0;WeightsStore[0][252]<=0;WeightsStore[0][253]<=0;WeightsStore[0][254]<=0;WeightsStore[0][255]<=0;WeightsStore[0][256]<=0;WeightsStore[0][257]<=0;WeightsStore[0][258]<=0;WeightsStore[0][259]<=0;WeightsStore[0][260]<=0;WeightsStore[0][261]<=0;WeightsStore[0][262]<=0;WeightsStore[0][263]<=0;WeightsStore[0][264]<=0;WeightsStore[0][265]<=0;WeightsStore[0][266]<=0;WeightsStore[0][267]<=0;WeightsStore[0][268]<=0;WeightsStore[0][269]<=0;WeightsStore[0][270]<=0;WeightsStore[0][271]<=0;WeightsStore[0][272]<=0;WeightsStore[0][273]<=0;WeightsStore[0][274]<=0;WeightsStore[0][275]<=0;WeightsStore[0][276]<=0;WeightsStore[0][277]<=0;WeightsStore[0][278]<=0;WeightsStore[0][279]<=0;WeightsStore[0][280]<=0;WeightsStore[0][281]<=0;WeightsStore[0][282]<=0;WeightsStore[0][283]<=0;WeightsStore[0][284]<=0;WeightsStore[0][285]<=0;WeightsStore[0][286]<=0;WeightsStore[0][287]<=0;WeightsStore[0][288]<=0;WeightsStore[0][289]<=0;WeightsStore[0][290]<=0;WeightsStore[0][291]<=0;WeightsStore[0][292]<=0;WeightsStore[0][293]<=0;WeightsStore[0][294]<=0;WeightsStore[0][295]<=0;WeightsStore[0][296]<=0;WeightsStore[0][297]<=0;WeightsStore[0][298]<=0;WeightsStore[0][299]<=0;WeightsStore[0][300]<=0;WeightsStore[0][301]<=0;WeightsStore[0][302]<=0;WeightsStore[0][303]<=0;WeightsStore[0][304]<=0;WeightsStore[0][305]<=0;WeightsStore[0][306]<=0;WeightsStore[0][307]<=0;WeightsStore[0][308]<=0;WeightsStore[0][309]<=0;WeightsStore[0][310]<=0;WeightsStore[0][311]<=0;WeightsStore[0][312]<=0;WeightsStore[0][313]<=0;WeightsStore[0][314]<=0;WeightsStore[0][315]<=0;WeightsStore[0][316]<=0;WeightsStore[0][317]<=0;WeightsStore[0][318]<=0;WeightsStore[0][319]<=0;WeightsStore[0][320]<=0;WeightsStore[0][321]<=0;WeightsStore[0][322]<=0;WeightsStore[0][323]<=0;WeightsStore[0][324]<=0;WeightsStore[0][325]<=0;WeightsStore[0][326]<=0;WeightsStore[0][327]<=0;WeightsStore[0][328]<=0;WeightsStore[0][329]<=0;WeightsStore[0][330]<=0;WeightsStore[0][331]<=0;WeightsStore[0][332]<=0;WeightsStore[0][333]<=0;WeightsStore[0][334]<=0;WeightsStore[0][335]<=0;WeightsStore[0][336]<=0;WeightsStore[0][337]<=0;WeightsStore[0][338]<=0;WeightsStore[0][339]<=0;WeightsStore[0][340]<=0;WeightsStore[0][341]<=0;WeightsStore[0][342]<=0;WeightsStore[0][343]<=0;WeightsStore[0][344]<=0;WeightsStore[0][345]<=0;WeightsStore[0][346]<=0;WeightsStore[0][347]<=0;WeightsStore[0][348]<=0;WeightsStore[0][349]<=0;WeightsStore[0][350]<=0;WeightsStore[0][351]<=0;WeightsStore[0][352]<=0;WeightsStore[0][353]<=0;WeightsStore[0][354]<=0;WeightsStore[0][355]<=0;WeightsStore[0][356]<=0;WeightsStore[0][357]<=0;WeightsStore[0][358]<=0;WeightsStore[0][359]<=0;WeightsStore[0][360]<=0;WeightsStore[0][361]<=0;WeightsStore[0][362]<=0;WeightsStore[0][363]<=0;WeightsStore[0][364]<=0;WeightsStore[0][365]<=0;WeightsStore[0][366]<=0;WeightsStore[0][367]<=0;WeightsStore[0][368]<=0;WeightsStore[0][369]<=0;WeightsStore[0][370]<=0;WeightsStore[0][371]<=0;WeightsStore[0][372]<=0;WeightsStore[0][373]<=0;WeightsStore[0][374]<=0;WeightsStore[0][375]<=0;WeightsStore[0][376]<=0;WeightsStore[0][377]<=0;WeightsStore[0][378]<=0;WeightsStore[0][379]<=0;WeightsStore[0][380]<=0;WeightsStore[0][381]<=0;WeightsStore[0][382]<=0;WeightsStore[0][383]<=0;WeightsStore[0][384]<=0;WeightsStore[0][385]<=0;WeightsStore[0][386]<=0;WeightsStore[0][387]<=0;WeightsStore[0][388]<=0;WeightsStore[0][389]<=0;WeightsStore[0][390]<=0;WeightsStore[0][391]<=0;WeightsStore[0][392]<=0;WeightsStore[0][393]<=0;WeightsStore[0][394]<=0;WeightsStore[0][395]<=0;WeightsStore[0][396]<=0;WeightsStore[0][397]<=0;WeightsStore[0][398]<=0;WeightsStore[0][399]<=0;WeightsStore[0][400]<=0;WeightsStore[0][401]<=0;WeightsStore[0][402]<=0;WeightsStore[0][403]<=0;WeightsStore[0][404]<=0;WeightsStore[0][405]<=0;WeightsStore[0][406]<=0;WeightsStore[0][407]<=0;WeightsStore[0][408]<=0;WeightsStore[0][409]<=0;WeightsStore[0][410]<=0;WeightsStore[0][411]<=0;WeightsStore[0][412]<=0;WeightsStore[0][413]<=0;WeightsStore[0][414]<=0;WeightsStore[0][415]<=0;WeightsStore[0][416]<=0;WeightsStore[0][417]<=0;WeightsStore[0][418]<=0;WeightsStore[0][419]<=0;WeightsStore[0][420]<=0;WeightsStore[0][421]<=0;WeightsStore[0][422]<=0;WeightsStore[0][423]<=0;WeightsStore[0][424]<=0;WeightsStore[0][425]<=0;WeightsStore[0][426]<=0;WeightsStore[0][427]<=0;WeightsStore[0][428]<=0;WeightsStore[0][429]<=0;WeightsStore[0][430]<=0;WeightsStore[0][431]<=0;WeightsStore[0][432]<=0;WeightsStore[0][433]<=0;WeightsStore[0][434]<=0;WeightsStore[0][435]<=0;WeightsStore[0][436]<=0;WeightsStore[0][437]<=0;WeightsStore[0][438]<=0;WeightsStore[0][439]<=0;WeightsStore[0][440]<=0;WeightsStore[0][441]<=0;WeightsStore[0][442]<=0;WeightsStore[0][443]<=0;WeightsStore[0][444]<=0;WeightsStore[0][445]<=0;WeightsStore[0][446]<=0;WeightsStore[0][447]<=0;WeightsStore[0][448]<=0;WeightsStore[0][449]<=0;WeightsStore[0][450]<=0;WeightsStore[0][451]<=0;WeightsStore[0][452]<=0;WeightsStore[0][453]<=0;WeightsStore[0][454]<=0;WeightsStore[0][455]<=0;WeightsStore[0][456]<=0;WeightsStore[0][457]<=0;WeightsStore[0][458]<=0;WeightsStore[0][459]<=0;WeightsStore[0][460]<=0;WeightsStore[0][461]<=0;WeightsStore[0][462]<=0;WeightsStore[0][463]<=0;WeightsStore[0][464]<=0;WeightsStore[0][465]<=0;WeightsStore[0][466]<=0;WeightsStore[0][467]<=0;WeightsStore[0][468]<=0;WeightsStore[0][469]<=0;WeightsStore[0][470]<=0;WeightsStore[0][471]<=0;WeightsStore[0][472]<=0;WeightsStore[0][473]<=0;WeightsStore[0][474]<=0;WeightsStore[0][475]<=0;WeightsStore[0][476]<=0;WeightsStore[0][477]<=0;WeightsStore[0][478]<=0;WeightsStore[0][479]<=0;WeightsStore[0][480]<=0;WeightsStore[0][481]<=0;WeightsStore[0][482]<=0;WeightsStore[0][483]<=0;WeightsStore[0][484]<=0;WeightsStore[0][485]<=0;WeightsStore[0][486]<=0;WeightsStore[0][487]<=0;WeightsStore[0][488]<=0;WeightsStore[0][489]<=0;WeightsStore[0][490]<=0;WeightsStore[0][491]<=0;WeightsStore[0][492]<=0;WeightsStore[0][493]<=0;WeightsStore[0][494]<=0;WeightsStore[0][495]<=0;WeightsStore[0][496]<=0;WeightsStore[0][497]<=0;WeightsStore[0][498]<=0;WeightsStore[0][499]<=0;WeightsStore[0][500]<=0;WeightsStore[0][501]<=0;WeightsStore[0][502]<=0;WeightsStore[0][503]<=0;WeightsStore[0][504]<=0;WeightsStore[0][505]<=0;WeightsStore[0][506]<=0;WeightsStore[0][507]<=0;WeightsStore[0][508]<=0;WeightsStore[0][509]<=0;WeightsStore[0][510]<=0;WeightsStore[0][511]<=0;WeightsStore[0][512]<=0;WeightsStore[0][513]<=0;WeightsStore[0][514]<=0;WeightsStore[0][515]<=0;WeightsStore[0][516]<=0;WeightsStore[0][517]<=0;WeightsStore[0][518]<=0;WeightsStore[0][519]<=0;WeightsStore[0][520]<=0;WeightsStore[0][521]<=0;WeightsStore[0][522]<=0;WeightsStore[0][523]<=0;WeightsStore[0][524]<=0;WeightsStore[0][525]<=0;WeightsStore[0][526]<=0;WeightsStore[0][527]<=0;WeightsStore[0][528]<=0;WeightsStore[0][529]<=0;WeightsStore[0][530]<=0;WeightsStore[0][531]<=0;WeightsStore[0][532]<=0;WeightsStore[0][533]<=0;WeightsStore[0][534]<=0;WeightsStore[0][535]<=0;WeightsStore[0][536]<=0;WeightsStore[0][537]<=0;WeightsStore[0][538]<=0;WeightsStore[0][539]<=0;WeightsStore[0][540]<=0;WeightsStore[0][541]<=0;WeightsStore[0][542]<=0;WeightsStore[0][543]<=0;WeightsStore[0][544]<=0;WeightsStore[0][545]<=0;WeightsStore[0][546]<=0;WeightsStore[0][547]<=0;WeightsStore[0][548]<=0;WeightsStore[0][549]<=0;WeightsStore[0][550]<=0;WeightsStore[0][551]<=0;WeightsStore[0][552]<=0;WeightsStore[0][553]<=0;WeightsStore[0][554]<=0;WeightsStore[0][555]<=0;WeightsStore[0][556]<=0;WeightsStore[0][557]<=0;WeightsStore[0][558]<=0;WeightsStore[0][559]<=0;WeightsStore[0][560]<=0;WeightsStore[0][561]<=0;WeightsStore[0][562]<=0;WeightsStore[0][563]<=0;WeightsStore[0][564]<=0;WeightsStore[0][565]<=0;WeightsStore[0][566]<=0;WeightsStore[0][567]<=0;WeightsStore[0][568]<=0;WeightsStore[0][569]<=0;WeightsStore[0][570]<=0;WeightsStore[0][571]<=0;WeightsStore[0][572]<=0;WeightsStore[0][573]<=0;WeightsStore[0][574]<=0;WeightsStore[0][575]<=0;WeightsStore[0][576]<=0;WeightsStore[0][577]<=0;WeightsStore[0][578]<=0;WeightsStore[0][579]<=0;WeightsStore[0][580]<=0;WeightsStore[0][581]<=0;WeightsStore[0][582]<=0;WeightsStore[0][583]<=0;WeightsStore[0][584]<=0;WeightsStore[0][585]<=0;WeightsStore[0][586]<=0;WeightsStore[0][587]<=0;WeightsStore[0][588]<=0;WeightsStore[0][589]<=0;WeightsStore[0][590]<=0;WeightsStore[0][591]<=0;WeightsStore[0][592]<=0;WeightsStore[0][593]<=0;WeightsStore[0][594]<=0;WeightsStore[0][595]<=0;WeightsStore[0][596]<=0;WeightsStore[0][597]<=0;WeightsStore[0][598]<=0;WeightsStore[0][599]<=0;WeightsStore[0][600]<=0;WeightsStore[0][601]<=0;WeightsStore[0][602]<=0;WeightsStore[0][603]<=0;WeightsStore[0][604]<=0;WeightsStore[0][605]<=0;WeightsStore[0][606]<=0;WeightsStore[0][607]<=0;WeightsStore[0][608]<=0;WeightsStore[0][609]<=0;WeightsStore[0][610]<=0;WeightsStore[0][611]<=0;WeightsStore[0][612]<=0;WeightsStore[0][613]<=0;WeightsStore[0][614]<=0;WeightsStore[0][615]<=0;WeightsStore[0][616]<=0;WeightsStore[0][617]<=0;WeightsStore[0][618]<=0;WeightsStore[0][619]<=0;WeightsStore[0][620]<=0;WeightsStore[0][621]<=0;WeightsStore[0][622]<=0;WeightsStore[0][623]<=0;WeightsStore[0][624]<=0;WeightsStore[0][625]<=0;WeightsStore[0][626]<=0;WeightsStore[0][627]<=0;WeightsStore[0][628]<=0;WeightsStore[0][629]<=0;WeightsStore[0][630]<=0;WeightsStore[0][631]<=0;WeightsStore[0][632]<=0;WeightsStore[0][633]<=0;WeightsStore[0][634]<=0;WeightsStore[0][635]<=0;WeightsStore[0][636]<=0;WeightsStore[0][637]<=0;WeightsStore[0][638]<=0;WeightsStore[0][639]<=0;WeightsStore[0][640]<=0;WeightsStore[0][641]<=0;WeightsStore[0][642]<=0;WeightsStore[0][643]<=0;WeightsStore[0][644]<=0;WeightsStore[0][645]<=0;WeightsStore[0][646]<=0;WeightsStore[0][647]<=0;WeightsStore[0][648]<=0;WeightsStore[0][649]<=0;WeightsStore[0][650]<=0;WeightsStore[0][651]<=0;WeightsStore[0][652]<=0;WeightsStore[0][653]<=0;WeightsStore[0][654]<=0;WeightsStore[0][655]<=0;WeightsStore[0][656]<=0;WeightsStore[0][657]<=0;WeightsStore[0][658]<=0;WeightsStore[0][659]<=0;WeightsStore[0][660]<=0;WeightsStore[0][661]<=0;WeightsStore[0][662]<=0;WeightsStore[0][663]<=0;WeightsStore[0][664]<=0;WeightsStore[0][665]<=0;WeightsStore[0][666]<=0;WeightsStore[0][667]<=0;WeightsStore[0][668]<=0;WeightsStore[0][669]<=0;WeightsStore[0][670]<=0;WeightsStore[0][671]<=0;WeightsStore[0][672]<=0;WeightsStore[0][673]<=0;WeightsStore[0][674]<=0;WeightsStore[0][675]<=0;WeightsStore[0][676]<=0;WeightsStore[0][677]<=0;WeightsStore[0][678]<=0;WeightsStore[0][679]<=0;WeightsStore[0][680]<=0;WeightsStore[0][681]<=0;WeightsStore[0][682]<=0;WeightsStore[0][683]<=0;WeightsStore[0][684]<=0;WeightsStore[0][685]<=0;WeightsStore[0][686]<=0;WeightsStore[0][687]<=0;WeightsStore[0][688]<=0;WeightsStore[0][689]<=0;WeightsStore[0][690]<=0;WeightsStore[0][691]<=0;WeightsStore[0][692]<=0;WeightsStore[0][693]<=0;WeightsStore[0][694]<=0;WeightsStore[0][695]<=0;WeightsStore[0][696]<=0;WeightsStore[0][697]<=0;WeightsStore[0][698]<=0;WeightsStore[0][699]<=0;WeightsStore[0][700]<=0;WeightsStore[0][701]<=0;WeightsStore[0][702]<=0;WeightsStore[0][703]<=0;WeightsStore[0][704]<=0;WeightsStore[0][705]<=0;WeightsStore[0][706]<=0;WeightsStore[0][707]<=0;WeightsStore[0][708]<=0;WeightsStore[0][709]<=0;WeightsStore[0][710]<=0;WeightsStore[0][711]<=0;WeightsStore[0][712]<=0;WeightsStore[0][713]<=0;WeightsStore[0][714]<=0;WeightsStore[0][715]<=0;WeightsStore[0][716]<=0;WeightsStore[0][717]<=0;WeightsStore[0][718]<=0;WeightsStore[0][719]<=0;WeightsStore[0][720]<=0;WeightsStore[0][721]<=0;WeightsStore[0][722]<=0;WeightsStore[0][723]<=0;WeightsStore[0][724]<=0;WeightsStore[0][725]<=0;WeightsStore[0][726]<=0;WeightsStore[0][727]<=0;WeightsStore[0][728]<=0;WeightsStore[0][729]<=0;WeightsStore[0][730]<=0;WeightsStore[0][731]<=0;WeightsStore[0][732]<=0;WeightsStore[0][733]<=0;WeightsStore[0][734]<=0;WeightsStore[0][735]<=0;WeightsStore[0][736]<=0;WeightsStore[0][737]<=0;WeightsStore[0][738]<=0;WeightsStore[0][739]<=0;WeightsStore[0][740]<=0;WeightsStore[0][741]<=0;WeightsStore[0][742]<=0;WeightsStore[0][743]<=0;WeightsStore[0][744]<=0;WeightsStore[0][745]<=0;WeightsStore[0][746]<=0;WeightsStore[0][747]<=0;WeightsStore[0][748]<=0;WeightsStore[0][749]<=0;WeightsStore[0][750]<=0;WeightsStore[0][751]<=0;WeightsStore[0][752]<=0;WeightsStore[0][753]<=0;WeightsStore[0][754]<=0;WeightsStore[0][755]<=0;WeightsStore[0][756]<=0;WeightsStore[0][757]<=0;WeightsStore[0][758]<=0;WeightsStore[0][759]<=0;WeightsStore[0][760]<=0;WeightsStore[0][761]<=0;WeightsStore[0][762]<=0;WeightsStore[0][763]<=0;WeightsStore[0][764]<=0;WeightsStore[0][765]<=0;WeightsStore[0][766]<=0;WeightsStore[0][767]<=0;WeightsStore[0][768]<=0;WeightsStore[0][769]<=0;WeightsStore[0][770]<=0;WeightsStore[0][771]<=0;WeightsStore[0][772]<=0;WeightsStore[0][773]<=0;WeightsStore[0][774]<=0;WeightsStore[0][775]<=0;WeightsStore[0][776]<=0;WeightsStore[0][777]<=0;WeightsStore[0][778]<=0;WeightsStore[0][779]<=0;WeightsStore[0][780]<=0;WeightsStore[0][781]<=0;WeightsStore[0][782]<=0;WeightsStore[0][783]<=0;WeightsStore[0][784]<=0;WeightsStore[1][0]<=0;WeightsStore[1][1]<=0;WeightsStore[1][2]<=0;WeightsStore[1][3]<=0;WeightsStore[1][4]<=0;WeightsStore[1][5]<=0;WeightsStore[1][6]<=0;WeightsStore[1][7]<=0;WeightsStore[1][8]<=0;WeightsStore[1][9]<=0;WeightsStore[1][10]<=0;WeightsStore[1][11]<=0;WeightsStore[1][12]<=0;WeightsStore[1][13]<=0;WeightsStore[1][14]<=0;WeightsStore[1][15]<=0;WeightsStore[1][16]<=0;WeightsStore[1][17]<=0;WeightsStore[1][18]<=0;WeightsStore[1][19]<=0;WeightsStore[1][20]<=0;WeightsStore[1][21]<=0;WeightsStore[1][22]<=0;WeightsStore[1][23]<=0;WeightsStore[1][24]<=0;WeightsStore[1][25]<=0;WeightsStore[1][26]<=0;WeightsStore[1][27]<=0;WeightsStore[1][28]<=0;WeightsStore[1][29]<=0;WeightsStore[1][30]<=0;WeightsStore[1][31]<=0;WeightsStore[1][32]<=0;WeightsStore[1][33]<=0;WeightsStore[1][34]<=0;WeightsStore[1][35]<=0;WeightsStore[1][36]<=0;WeightsStore[1][37]<=0;WeightsStore[1][38]<=0;WeightsStore[1][39]<=0;WeightsStore[1][40]<=0;WeightsStore[1][41]<=0;WeightsStore[1][42]<=0;WeightsStore[1][43]<=0;WeightsStore[1][44]<=0;WeightsStore[1][45]<=0;WeightsStore[1][46]<=0;WeightsStore[1][47]<=0;WeightsStore[1][48]<=0;WeightsStore[1][49]<=0;WeightsStore[1][50]<=0;WeightsStore[1][51]<=0;WeightsStore[1][52]<=0;WeightsStore[1][53]<=0;WeightsStore[1][54]<=0;WeightsStore[1][55]<=0;WeightsStore[1][56]<=0;WeightsStore[1][57]<=0;WeightsStore[1][58]<=0;WeightsStore[1][59]<=0;WeightsStore[1][60]<=0;WeightsStore[1][61]<=0;WeightsStore[1][62]<=0;WeightsStore[1][63]<=0;WeightsStore[1][64]<=0;WeightsStore[1][65]<=0;WeightsStore[1][66]<=0;WeightsStore[1][67]<=0;WeightsStore[1][68]<=0;WeightsStore[1][69]<=0;WeightsStore[1][70]<=0;WeightsStore[1][71]<=0;WeightsStore[1][72]<=0;WeightsStore[1][73]<=0;WeightsStore[1][74]<=0;WeightsStore[1][75]<=0;WeightsStore[1][76]<=0;WeightsStore[1][77]<=0;WeightsStore[1][78]<=0;WeightsStore[1][79]<=0;WeightsStore[1][80]<=0;WeightsStore[1][81]<=0;WeightsStore[1][82]<=0;WeightsStore[1][83]<=0;WeightsStore[1][84]<=0;WeightsStore[1][85]<=0;WeightsStore[1][86]<=0;WeightsStore[1][87]<=0;WeightsStore[1][88]<=0;WeightsStore[1][89]<=0;WeightsStore[1][90]<=0;WeightsStore[1][91]<=0;WeightsStore[1][92]<=0;WeightsStore[1][93]<=0;WeightsStore[1][94]<=0;WeightsStore[1][95]<=0;WeightsStore[1][96]<=0;WeightsStore[1][97]<=0;WeightsStore[1][98]<=0;WeightsStore[1][99]<=0;WeightsStore[1][100]<=0;WeightsStore[1][101]<=0;WeightsStore[1][102]<=0;WeightsStore[1][103]<=0;WeightsStore[1][104]<=0;WeightsStore[1][105]<=0;WeightsStore[1][106]<=0;WeightsStore[1][107]<=0;WeightsStore[1][108]<=0;WeightsStore[1][109]<=0;WeightsStore[1][110]<=0;WeightsStore[1][111]<=0;WeightsStore[1][112]<=0;WeightsStore[1][113]<=0;WeightsStore[1][114]<=0;WeightsStore[1][115]<=0;WeightsStore[1][116]<=0;WeightsStore[1][117]<=0;WeightsStore[1][118]<=0;WeightsStore[1][119]<=0;WeightsStore[1][120]<=0;WeightsStore[1][121]<=0;WeightsStore[1][122]<=0;WeightsStore[1][123]<=0;WeightsStore[1][124]<=0;WeightsStore[1][125]<=0;WeightsStore[1][126]<=0;WeightsStore[1][127]<=0;WeightsStore[1][128]<=0;WeightsStore[1][129]<=0;WeightsStore[1][130]<=0;WeightsStore[1][131]<=0;WeightsStore[1][132]<=0;WeightsStore[1][133]<=0;WeightsStore[1][134]<=0;WeightsStore[1][135]<=0;WeightsStore[1][136]<=0;WeightsStore[1][137]<=0;WeightsStore[1][138]<=0;WeightsStore[1][139]<=0;WeightsStore[1][140]<=0;WeightsStore[1][141]<=0;WeightsStore[1][142]<=0;WeightsStore[1][143]<=0;WeightsStore[1][144]<=0;WeightsStore[1][145]<=0;WeightsStore[1][146]<=0;WeightsStore[1][147]<=0;WeightsStore[1][148]<=0;WeightsStore[1][149]<=0;WeightsStore[1][150]<=0;WeightsStore[1][151]<=0;WeightsStore[1][152]<=0;WeightsStore[1][153]<=0;WeightsStore[1][154]<=0;WeightsStore[1][155]<=0;WeightsStore[1][156]<=0;WeightsStore[1][157]<=0;WeightsStore[1][158]<=0;WeightsStore[1][159]<=0;WeightsStore[1][160]<=0;WeightsStore[1][161]<=0;WeightsStore[1][162]<=0;WeightsStore[1][163]<=0;WeightsStore[1][164]<=0;WeightsStore[1][165]<=0;WeightsStore[1][166]<=0;WeightsStore[1][167]<=0;WeightsStore[1][168]<=0;WeightsStore[1][169]<=0;WeightsStore[1][170]<=0;WeightsStore[1][171]<=0;WeightsStore[1][172]<=0;WeightsStore[1][173]<=0;WeightsStore[1][174]<=0;WeightsStore[1][175]<=0;WeightsStore[1][176]<=0;WeightsStore[1][177]<=0;WeightsStore[1][178]<=0;WeightsStore[1][179]<=0;WeightsStore[1][180]<=0;WeightsStore[1][181]<=0;WeightsStore[1][182]<=0;WeightsStore[1][183]<=0;WeightsStore[1][184]<=0;WeightsStore[1][185]<=0;WeightsStore[1][186]<=0;WeightsStore[1][187]<=0;WeightsStore[1][188]<=0;WeightsStore[1][189]<=0;WeightsStore[1][190]<=0;WeightsStore[1][191]<=0;WeightsStore[1][192]<=0;WeightsStore[1][193]<=0;WeightsStore[1][194]<=0;WeightsStore[1][195]<=0;WeightsStore[1][196]<=0;WeightsStore[1][197]<=0;WeightsStore[1][198]<=0;WeightsStore[1][199]<=0;WeightsStore[1][200]<=0;WeightsStore[1][201]<=0;WeightsStore[1][202]<=0;WeightsStore[1][203]<=0;WeightsStore[1][204]<=0;WeightsStore[1][205]<=0;WeightsStore[1][206]<=0;WeightsStore[1][207]<=0;WeightsStore[1][208]<=0;WeightsStore[1][209]<=0;WeightsStore[1][210]<=0;WeightsStore[1][211]<=0;WeightsStore[1][212]<=0;WeightsStore[1][213]<=0;WeightsStore[1][214]<=0;WeightsStore[1][215]<=0;WeightsStore[1][216]<=0;WeightsStore[1][217]<=0;WeightsStore[1][218]<=0;WeightsStore[1][219]<=0;WeightsStore[1][220]<=0;WeightsStore[1][221]<=0;WeightsStore[1][222]<=0;WeightsStore[1][223]<=0;WeightsStore[1][224]<=0;WeightsStore[1][225]<=0;WeightsStore[1][226]<=0;WeightsStore[1][227]<=0;WeightsStore[1][228]<=0;WeightsStore[1][229]<=0;WeightsStore[1][230]<=0;WeightsStore[1][231]<=0;WeightsStore[1][232]<=0;WeightsStore[1][233]<=0;WeightsStore[1][234]<=0;WeightsStore[1][235]<=0;WeightsStore[1][236]<=0;WeightsStore[1][237]<=0;WeightsStore[1][238]<=0;WeightsStore[1][239]<=0;WeightsStore[1][240]<=0;WeightsStore[1][241]<=0;WeightsStore[1][242]<=0;WeightsStore[1][243]<=0;WeightsStore[1][244]<=0;WeightsStore[1][245]<=0;WeightsStore[1][246]<=0;WeightsStore[1][247]<=0;WeightsStore[1][248]<=0;WeightsStore[1][249]<=0;WeightsStore[1][250]<=0;WeightsStore[1][251]<=0;WeightsStore[1][252]<=0;WeightsStore[1][253]<=0;WeightsStore[1][254]<=0;WeightsStore[1][255]<=0;WeightsStore[1][256]<=0;WeightsStore[1][257]<=0;WeightsStore[1][258]<=0;WeightsStore[1][259]<=0;WeightsStore[1][260]<=0;WeightsStore[1][261]<=0;WeightsStore[1][262]<=0;WeightsStore[1][263]<=0;WeightsStore[1][264]<=0;WeightsStore[1][265]<=0;WeightsStore[1][266]<=0;WeightsStore[1][267]<=0;WeightsStore[1][268]<=0;WeightsStore[1][269]<=0;WeightsStore[1][270]<=0;WeightsStore[1][271]<=0;WeightsStore[1][272]<=0;WeightsStore[1][273]<=0;WeightsStore[1][274]<=0;WeightsStore[1][275]<=0;WeightsStore[1][276]<=0;WeightsStore[1][277]<=0;WeightsStore[1][278]<=0;WeightsStore[1][279]<=0;WeightsStore[1][280]<=0;WeightsStore[1][281]<=0;WeightsStore[1][282]<=0;WeightsStore[1][283]<=0;WeightsStore[1][284]<=0;WeightsStore[1][285]<=0;WeightsStore[1][286]<=0;WeightsStore[1][287]<=0;WeightsStore[1][288]<=0;WeightsStore[1][289]<=0;WeightsStore[1][290]<=0;WeightsStore[1][291]<=0;WeightsStore[1][292]<=0;WeightsStore[1][293]<=0;WeightsStore[1][294]<=0;WeightsStore[1][295]<=0;WeightsStore[1][296]<=0;WeightsStore[1][297]<=0;WeightsStore[1][298]<=0;WeightsStore[1][299]<=0;WeightsStore[1][300]<=0;WeightsStore[1][301]<=0;WeightsStore[1][302]<=0;WeightsStore[1][303]<=0;WeightsStore[1][304]<=0;WeightsStore[1][305]<=0;WeightsStore[1][306]<=0;WeightsStore[1][307]<=0;WeightsStore[1][308]<=0;WeightsStore[1][309]<=0;WeightsStore[1][310]<=0;WeightsStore[1][311]<=0;WeightsStore[1][312]<=0;WeightsStore[1][313]<=0;WeightsStore[1][314]<=0;WeightsStore[1][315]<=0;WeightsStore[1][316]<=0;WeightsStore[1][317]<=0;WeightsStore[1][318]<=0;WeightsStore[1][319]<=0;WeightsStore[1][320]<=0;WeightsStore[1][321]<=0;WeightsStore[1][322]<=0;WeightsStore[1][323]<=0;WeightsStore[1][324]<=0;WeightsStore[1][325]<=0;WeightsStore[1][326]<=0;WeightsStore[1][327]<=0;WeightsStore[1][328]<=0;WeightsStore[1][329]<=0;WeightsStore[1][330]<=0;WeightsStore[1][331]<=0;WeightsStore[1][332]<=0;WeightsStore[1][333]<=0;WeightsStore[1][334]<=0;WeightsStore[1][335]<=0;WeightsStore[1][336]<=0;WeightsStore[1][337]<=0;WeightsStore[1][338]<=0;WeightsStore[1][339]<=0;WeightsStore[1][340]<=0;WeightsStore[1][341]<=0;WeightsStore[1][342]<=0;WeightsStore[1][343]<=0;WeightsStore[1][344]<=0;WeightsStore[1][345]<=0;WeightsStore[1][346]<=0;WeightsStore[1][347]<=0;WeightsStore[1][348]<=0;WeightsStore[1][349]<=0;WeightsStore[1][350]<=0;WeightsStore[1][351]<=0;WeightsStore[1][352]<=0;WeightsStore[1][353]<=0;WeightsStore[1][354]<=0;WeightsStore[1][355]<=0;WeightsStore[1][356]<=0;WeightsStore[1][357]<=0;WeightsStore[1][358]<=0;WeightsStore[1][359]<=0;WeightsStore[1][360]<=0;WeightsStore[1][361]<=0;WeightsStore[1][362]<=0;WeightsStore[1][363]<=0;WeightsStore[1][364]<=0;WeightsStore[1][365]<=0;WeightsStore[1][366]<=0;WeightsStore[1][367]<=0;WeightsStore[1][368]<=0;WeightsStore[1][369]<=0;WeightsStore[1][370]<=0;WeightsStore[1][371]<=0;WeightsStore[1][372]<=0;WeightsStore[1][373]<=0;WeightsStore[1][374]<=0;WeightsStore[1][375]<=0;WeightsStore[1][376]<=0;WeightsStore[1][377]<=0;WeightsStore[1][378]<=0;WeightsStore[1][379]<=0;WeightsStore[1][380]<=0;WeightsStore[1][381]<=0;WeightsStore[1][382]<=0;WeightsStore[1][383]<=0;WeightsStore[1][384]<=0;WeightsStore[1][385]<=0;WeightsStore[1][386]<=0;WeightsStore[1][387]<=0;WeightsStore[1][388]<=0;WeightsStore[1][389]<=0;WeightsStore[1][390]<=0;WeightsStore[1][391]<=0;WeightsStore[1][392]<=0;WeightsStore[1][393]<=0;WeightsStore[1][394]<=0;WeightsStore[1][395]<=0;WeightsStore[1][396]<=0;WeightsStore[1][397]<=0;WeightsStore[1][398]<=0;WeightsStore[1][399]<=0;WeightsStore[1][400]<=0;WeightsStore[1][401]<=0;WeightsStore[1][402]<=0;WeightsStore[1][403]<=0;WeightsStore[1][404]<=0;WeightsStore[1][405]<=0;WeightsStore[1][406]<=0;WeightsStore[1][407]<=0;WeightsStore[1][408]<=0;WeightsStore[1][409]<=0;WeightsStore[1][410]<=0;WeightsStore[1][411]<=0;WeightsStore[1][412]<=0;WeightsStore[1][413]<=0;WeightsStore[1][414]<=0;WeightsStore[1][415]<=0;WeightsStore[1][416]<=0;WeightsStore[1][417]<=0;WeightsStore[1][418]<=0;WeightsStore[1][419]<=0;WeightsStore[1][420]<=0;WeightsStore[1][421]<=0;WeightsStore[1][422]<=0;WeightsStore[1][423]<=0;WeightsStore[1][424]<=0;WeightsStore[1][425]<=0;WeightsStore[1][426]<=0;WeightsStore[1][427]<=0;WeightsStore[1][428]<=0;WeightsStore[1][429]<=0;WeightsStore[1][430]<=0;WeightsStore[1][431]<=0;WeightsStore[1][432]<=0;WeightsStore[1][433]<=0;WeightsStore[1][434]<=0;WeightsStore[1][435]<=0;WeightsStore[1][436]<=0;WeightsStore[1][437]<=0;WeightsStore[1][438]<=0;WeightsStore[1][439]<=0;WeightsStore[1][440]<=0;WeightsStore[1][441]<=0;WeightsStore[1][442]<=0;WeightsStore[1][443]<=0;WeightsStore[1][444]<=0;WeightsStore[1][445]<=0;WeightsStore[1][446]<=0;WeightsStore[1][447]<=0;WeightsStore[1][448]<=0;WeightsStore[1][449]<=0;WeightsStore[1][450]<=0;WeightsStore[1][451]<=0;WeightsStore[1][452]<=0;WeightsStore[1][453]<=0;WeightsStore[1][454]<=0;WeightsStore[1][455]<=0;WeightsStore[1][456]<=0;WeightsStore[1][457]<=0;WeightsStore[1][458]<=0;WeightsStore[1][459]<=0;WeightsStore[1][460]<=0;WeightsStore[1][461]<=0;WeightsStore[1][462]<=0;WeightsStore[1][463]<=0;WeightsStore[1][464]<=0;WeightsStore[1][465]<=0;WeightsStore[1][466]<=0;WeightsStore[1][467]<=0;WeightsStore[1][468]<=0;WeightsStore[1][469]<=0;WeightsStore[1][470]<=0;WeightsStore[1][471]<=0;WeightsStore[1][472]<=0;WeightsStore[1][473]<=0;WeightsStore[1][474]<=0;WeightsStore[1][475]<=0;WeightsStore[1][476]<=0;WeightsStore[1][477]<=0;WeightsStore[1][478]<=0;WeightsStore[1][479]<=0;WeightsStore[1][480]<=0;WeightsStore[1][481]<=0;WeightsStore[1][482]<=0;WeightsStore[1][483]<=0;WeightsStore[1][484]<=0;WeightsStore[1][485]<=0;WeightsStore[1][486]<=0;WeightsStore[1][487]<=0;WeightsStore[1][488]<=0;WeightsStore[1][489]<=0;WeightsStore[1][490]<=0;WeightsStore[1][491]<=0;WeightsStore[1][492]<=0;WeightsStore[1][493]<=0;WeightsStore[1][494]<=0;WeightsStore[1][495]<=0;WeightsStore[1][496]<=0;WeightsStore[1][497]<=0;WeightsStore[1][498]<=0;WeightsStore[1][499]<=0;WeightsStore[1][500]<=0;WeightsStore[1][501]<=0;WeightsStore[1][502]<=0;WeightsStore[1][503]<=0;WeightsStore[1][504]<=0;WeightsStore[1][505]<=0;WeightsStore[1][506]<=0;WeightsStore[1][507]<=0;WeightsStore[1][508]<=0;WeightsStore[1][509]<=0;WeightsStore[1][510]<=0;WeightsStore[1][511]<=0;WeightsStore[1][512]<=0;WeightsStore[1][513]<=0;WeightsStore[1][514]<=0;WeightsStore[1][515]<=0;WeightsStore[1][516]<=0;WeightsStore[1][517]<=0;WeightsStore[1][518]<=0;WeightsStore[1][519]<=0;WeightsStore[1][520]<=0;WeightsStore[1][521]<=0;WeightsStore[1][522]<=0;WeightsStore[1][523]<=0;WeightsStore[1][524]<=0;WeightsStore[1][525]<=0;WeightsStore[1][526]<=0;WeightsStore[1][527]<=0;WeightsStore[1][528]<=0;WeightsStore[1][529]<=0;WeightsStore[1][530]<=0;WeightsStore[1][531]<=0;WeightsStore[1][532]<=0;WeightsStore[1][533]<=0;WeightsStore[1][534]<=0;WeightsStore[1][535]<=0;WeightsStore[1][536]<=0;WeightsStore[1][537]<=0;WeightsStore[1][538]<=0;WeightsStore[1][539]<=0;WeightsStore[1][540]<=0;WeightsStore[1][541]<=0;WeightsStore[1][542]<=0;WeightsStore[1][543]<=0;WeightsStore[1][544]<=0;WeightsStore[1][545]<=0;WeightsStore[1][546]<=0;WeightsStore[1][547]<=0;WeightsStore[1][548]<=0;WeightsStore[1][549]<=0;WeightsStore[1][550]<=0;WeightsStore[1][551]<=0;WeightsStore[1][552]<=0;WeightsStore[1][553]<=0;WeightsStore[1][554]<=0;WeightsStore[1][555]<=0;WeightsStore[1][556]<=0;WeightsStore[1][557]<=0;WeightsStore[1][558]<=0;WeightsStore[1][559]<=0;WeightsStore[1][560]<=0;WeightsStore[1][561]<=0;WeightsStore[1][562]<=0;WeightsStore[1][563]<=0;WeightsStore[1][564]<=0;WeightsStore[1][565]<=0;WeightsStore[1][566]<=0;WeightsStore[1][567]<=0;WeightsStore[1][568]<=0;WeightsStore[1][569]<=0;WeightsStore[1][570]<=0;WeightsStore[1][571]<=0;WeightsStore[1][572]<=0;WeightsStore[1][573]<=0;WeightsStore[1][574]<=0;WeightsStore[1][575]<=0;WeightsStore[1][576]<=0;WeightsStore[1][577]<=0;WeightsStore[1][578]<=0;WeightsStore[1][579]<=0;WeightsStore[1][580]<=0;WeightsStore[1][581]<=0;WeightsStore[1][582]<=0;WeightsStore[1][583]<=0;WeightsStore[1][584]<=0;WeightsStore[1][585]<=0;WeightsStore[1][586]<=0;WeightsStore[1][587]<=0;WeightsStore[1][588]<=0;WeightsStore[1][589]<=0;WeightsStore[1][590]<=0;WeightsStore[1][591]<=0;WeightsStore[1][592]<=0;WeightsStore[1][593]<=0;WeightsStore[1][594]<=0;WeightsStore[1][595]<=0;WeightsStore[1][596]<=0;WeightsStore[1][597]<=0;WeightsStore[1][598]<=0;WeightsStore[1][599]<=0;WeightsStore[1][600]<=0;WeightsStore[1][601]<=0;WeightsStore[1][602]<=0;WeightsStore[1][603]<=0;WeightsStore[1][604]<=0;WeightsStore[1][605]<=0;WeightsStore[1][606]<=0;WeightsStore[1][607]<=0;WeightsStore[1][608]<=0;WeightsStore[1][609]<=0;WeightsStore[1][610]<=0;WeightsStore[1][611]<=0;WeightsStore[1][612]<=0;WeightsStore[1][613]<=0;WeightsStore[1][614]<=0;WeightsStore[1][615]<=0;WeightsStore[1][616]<=0;WeightsStore[1][617]<=0;WeightsStore[1][618]<=0;WeightsStore[1][619]<=0;WeightsStore[1][620]<=0;WeightsStore[1][621]<=0;WeightsStore[1][622]<=0;WeightsStore[1][623]<=0;WeightsStore[1][624]<=0;WeightsStore[1][625]<=0;WeightsStore[1][626]<=0;WeightsStore[1][627]<=0;WeightsStore[1][628]<=0;WeightsStore[1][629]<=0;WeightsStore[1][630]<=0;WeightsStore[1][631]<=0;WeightsStore[1][632]<=0;WeightsStore[1][633]<=0;WeightsStore[1][634]<=0;WeightsStore[1][635]<=0;WeightsStore[1][636]<=0;WeightsStore[1][637]<=0;WeightsStore[1][638]<=0;WeightsStore[1][639]<=0;WeightsStore[1][640]<=0;WeightsStore[1][641]<=0;WeightsStore[1][642]<=0;WeightsStore[1][643]<=0;WeightsStore[1][644]<=0;WeightsStore[1][645]<=0;WeightsStore[1][646]<=0;WeightsStore[1][647]<=0;WeightsStore[1][648]<=0;WeightsStore[1][649]<=0;WeightsStore[1][650]<=0;WeightsStore[1][651]<=0;WeightsStore[1][652]<=0;WeightsStore[1][653]<=0;WeightsStore[1][654]<=0;WeightsStore[1][655]<=0;WeightsStore[1][656]<=0;WeightsStore[1][657]<=0;WeightsStore[1][658]<=0;WeightsStore[1][659]<=0;WeightsStore[1][660]<=0;WeightsStore[1][661]<=0;WeightsStore[1][662]<=0;WeightsStore[1][663]<=0;WeightsStore[1][664]<=0;WeightsStore[1][665]<=0;WeightsStore[1][666]<=0;WeightsStore[1][667]<=0;WeightsStore[1][668]<=0;WeightsStore[1][669]<=0;WeightsStore[1][670]<=0;WeightsStore[1][671]<=0;WeightsStore[1][672]<=0;WeightsStore[1][673]<=0;WeightsStore[1][674]<=0;WeightsStore[1][675]<=0;WeightsStore[1][676]<=0;WeightsStore[1][677]<=0;WeightsStore[1][678]<=0;WeightsStore[1][679]<=0;WeightsStore[1][680]<=0;WeightsStore[1][681]<=0;WeightsStore[1][682]<=0;WeightsStore[1][683]<=0;WeightsStore[1][684]<=0;WeightsStore[1][685]<=0;WeightsStore[1][686]<=0;WeightsStore[1][687]<=0;WeightsStore[1][688]<=0;WeightsStore[1][689]<=0;WeightsStore[1][690]<=0;WeightsStore[1][691]<=0;WeightsStore[1][692]<=0;WeightsStore[1][693]<=0;WeightsStore[1][694]<=0;WeightsStore[1][695]<=0;WeightsStore[1][696]<=0;WeightsStore[1][697]<=0;WeightsStore[1][698]<=0;WeightsStore[1][699]<=0;WeightsStore[1][700]<=0;WeightsStore[1][701]<=0;WeightsStore[1][702]<=0;WeightsStore[1][703]<=0;WeightsStore[1][704]<=0;WeightsStore[1][705]<=0;WeightsStore[1][706]<=0;WeightsStore[1][707]<=0;WeightsStore[1][708]<=0;WeightsStore[1][709]<=0;WeightsStore[1][710]<=0;WeightsStore[1][711]<=0;WeightsStore[1][712]<=0;WeightsStore[1][713]<=0;WeightsStore[1][714]<=0;WeightsStore[1][715]<=0;WeightsStore[1][716]<=0;WeightsStore[1][717]<=0;WeightsStore[1][718]<=0;WeightsStore[1][719]<=0;WeightsStore[1][720]<=0;WeightsStore[1][721]<=0;WeightsStore[1][722]<=0;WeightsStore[1][723]<=0;WeightsStore[1][724]<=0;WeightsStore[1][725]<=0;WeightsStore[1][726]<=0;WeightsStore[1][727]<=0;WeightsStore[1][728]<=0;WeightsStore[1][729]<=0;WeightsStore[1][730]<=0;WeightsStore[1][731]<=0;WeightsStore[1][732]<=0;WeightsStore[1][733]<=0;WeightsStore[1][734]<=0;WeightsStore[1][735]<=0;WeightsStore[1][736]<=0;WeightsStore[1][737]<=0;WeightsStore[1][738]<=0;WeightsStore[1][739]<=0;WeightsStore[1][740]<=0;WeightsStore[1][741]<=0;WeightsStore[1][742]<=0;WeightsStore[1][743]<=0;WeightsStore[1][744]<=0;WeightsStore[1][745]<=0;WeightsStore[1][746]<=0;WeightsStore[1][747]<=0;WeightsStore[1][748]<=0;WeightsStore[1][749]<=0;WeightsStore[1][750]<=0;WeightsStore[1][751]<=0;WeightsStore[1][752]<=0;WeightsStore[1][753]<=0;WeightsStore[1][754]<=0;WeightsStore[1][755]<=0;WeightsStore[1][756]<=0;WeightsStore[1][757]<=0;WeightsStore[1][758]<=0;WeightsStore[1][759]<=0;WeightsStore[1][760]<=0;WeightsStore[1][761]<=0;WeightsStore[1][762]<=0;WeightsStore[1][763]<=0;WeightsStore[1][764]<=0;WeightsStore[1][765]<=0;WeightsStore[1][766]<=0;WeightsStore[1][767]<=0;WeightsStore[1][768]<=0;WeightsStore[1][769]<=0;WeightsStore[1][770]<=0;WeightsStore[1][771]<=0;WeightsStore[1][772]<=0;WeightsStore[1][773]<=0;WeightsStore[1][774]<=0;WeightsStore[1][775]<=0;WeightsStore[1][776]<=0;WeightsStore[1][777]<=0;WeightsStore[1][778]<=0;WeightsStore[1][779]<=0;WeightsStore[1][780]<=0;WeightsStore[1][781]<=0;WeightsStore[1][782]<=0;WeightsStore[1][783]<=0;WeightsStore[1][784]<=0;WeightsStore[2][0]<=0;WeightsStore[2][1]<=0;WeightsStore[2][2]<=0;WeightsStore[2][3]<=0;WeightsStore[2][4]<=0;WeightsStore[2][5]<=0;WeightsStore[2][6]<=0;WeightsStore[2][7]<=0;WeightsStore[2][8]<=0;WeightsStore[2][9]<=0;WeightsStore[2][10]<=0;WeightsStore[2][11]<=0;WeightsStore[2][12]<=0;WeightsStore[2][13]<=0;WeightsStore[2][14]<=0;WeightsStore[2][15]<=0;WeightsStore[2][16]<=0;WeightsStore[2][17]<=0;WeightsStore[2][18]<=0;WeightsStore[2][19]<=0;WeightsStore[2][20]<=0;WeightsStore[2][21]<=0;WeightsStore[2][22]<=0;WeightsStore[2][23]<=0;WeightsStore[2][24]<=0;WeightsStore[2][25]<=0;WeightsStore[2][26]<=0;WeightsStore[2][27]<=0;WeightsStore[2][28]<=0;WeightsStore[2][29]<=0;WeightsStore[2][30]<=0;WeightsStore[2][31]<=0;WeightsStore[2][32]<=0;WeightsStore[2][33]<=0;WeightsStore[2][34]<=0;WeightsStore[2][35]<=0;WeightsStore[2][36]<=0;WeightsStore[2][37]<=0;WeightsStore[2][38]<=0;WeightsStore[2][39]<=0;WeightsStore[2][40]<=0;WeightsStore[2][41]<=0;WeightsStore[2][42]<=0;WeightsStore[2][43]<=0;WeightsStore[2][44]<=0;WeightsStore[2][45]<=0;WeightsStore[2][46]<=0;WeightsStore[2][47]<=0;WeightsStore[2][48]<=0;WeightsStore[2][49]<=0;WeightsStore[2][50]<=0;WeightsStore[2][51]<=0;WeightsStore[2][52]<=0;WeightsStore[2][53]<=0;WeightsStore[2][54]<=0;WeightsStore[2][55]<=0;WeightsStore[2][56]<=0;WeightsStore[2][57]<=0;WeightsStore[2][58]<=0;WeightsStore[2][59]<=0;WeightsStore[2][60]<=0;WeightsStore[2][61]<=0;WeightsStore[2][62]<=0;WeightsStore[2][63]<=0;WeightsStore[2][64]<=0;WeightsStore[2][65]<=0;WeightsStore[2][66]<=0;WeightsStore[2][67]<=0;WeightsStore[2][68]<=0;WeightsStore[2][69]<=0;WeightsStore[2][70]<=0;WeightsStore[2][71]<=0;WeightsStore[2][72]<=0;WeightsStore[2][73]<=0;WeightsStore[2][74]<=0;WeightsStore[2][75]<=0;WeightsStore[2][76]<=0;WeightsStore[2][77]<=0;WeightsStore[2][78]<=0;WeightsStore[2][79]<=0;WeightsStore[2][80]<=0;WeightsStore[2][81]<=0;WeightsStore[2][82]<=0;WeightsStore[2][83]<=0;WeightsStore[2][84]<=0;WeightsStore[2][85]<=0;WeightsStore[2][86]<=0;WeightsStore[2][87]<=0;WeightsStore[2][88]<=0;WeightsStore[2][89]<=0;WeightsStore[2][90]<=0;WeightsStore[2][91]<=0;WeightsStore[2][92]<=0;WeightsStore[2][93]<=0;WeightsStore[2][94]<=0;WeightsStore[2][95]<=0;WeightsStore[2][96]<=0;WeightsStore[2][97]<=0;WeightsStore[2][98]<=0;WeightsStore[2][99]<=0;WeightsStore[2][100]<=0;WeightsStore[2][101]<=0;WeightsStore[2][102]<=0;WeightsStore[2][103]<=0;WeightsStore[2][104]<=0;WeightsStore[2][105]<=0;WeightsStore[2][106]<=0;WeightsStore[2][107]<=0;WeightsStore[2][108]<=0;WeightsStore[2][109]<=0;WeightsStore[2][110]<=0;WeightsStore[2][111]<=0;WeightsStore[2][112]<=0;WeightsStore[2][113]<=0;WeightsStore[2][114]<=0;WeightsStore[2][115]<=0;WeightsStore[2][116]<=0;WeightsStore[2][117]<=0;WeightsStore[2][118]<=0;WeightsStore[2][119]<=0;WeightsStore[2][120]<=0;WeightsStore[2][121]<=0;WeightsStore[2][122]<=0;WeightsStore[2][123]<=0;WeightsStore[2][124]<=0;WeightsStore[2][125]<=0;WeightsStore[2][126]<=0;WeightsStore[2][127]<=0;WeightsStore[2][128]<=0;WeightsStore[2][129]<=0;WeightsStore[2][130]<=0;WeightsStore[2][131]<=0;WeightsStore[2][132]<=0;WeightsStore[2][133]<=0;WeightsStore[2][134]<=0;WeightsStore[2][135]<=0;WeightsStore[2][136]<=0;WeightsStore[2][137]<=0;WeightsStore[2][138]<=0;WeightsStore[2][139]<=0;WeightsStore[2][140]<=0;WeightsStore[2][141]<=0;WeightsStore[2][142]<=0;WeightsStore[2][143]<=0;WeightsStore[2][144]<=0;WeightsStore[2][145]<=0;WeightsStore[2][146]<=0;WeightsStore[2][147]<=0;WeightsStore[2][148]<=0;WeightsStore[2][149]<=0;WeightsStore[2][150]<=0;WeightsStore[2][151]<=0;WeightsStore[2][152]<=0;WeightsStore[2][153]<=0;WeightsStore[2][154]<=0;WeightsStore[2][155]<=0;WeightsStore[2][156]<=0;WeightsStore[2][157]<=0;WeightsStore[2][158]<=0;WeightsStore[2][159]<=0;WeightsStore[2][160]<=0;WeightsStore[2][161]<=0;WeightsStore[2][162]<=0;WeightsStore[2][163]<=0;WeightsStore[2][164]<=0;WeightsStore[2][165]<=0;WeightsStore[2][166]<=0;WeightsStore[2][167]<=0;WeightsStore[2][168]<=0;WeightsStore[2][169]<=0;WeightsStore[2][170]<=0;WeightsStore[2][171]<=0;WeightsStore[2][172]<=0;WeightsStore[2][173]<=0;WeightsStore[2][174]<=0;WeightsStore[2][175]<=0;WeightsStore[2][176]<=0;WeightsStore[2][177]<=0;WeightsStore[2][178]<=0;WeightsStore[2][179]<=0;WeightsStore[2][180]<=0;WeightsStore[2][181]<=0;WeightsStore[2][182]<=0;WeightsStore[2][183]<=0;WeightsStore[2][184]<=0;WeightsStore[2][185]<=0;WeightsStore[2][186]<=0;WeightsStore[2][187]<=0;WeightsStore[2][188]<=0;WeightsStore[2][189]<=0;WeightsStore[2][190]<=0;WeightsStore[2][191]<=0;WeightsStore[2][192]<=0;WeightsStore[2][193]<=0;WeightsStore[2][194]<=0;WeightsStore[2][195]<=0;WeightsStore[2][196]<=0;WeightsStore[2][197]<=0;WeightsStore[2][198]<=0;WeightsStore[2][199]<=0;WeightsStore[2][200]<=0;WeightsStore[2][201]<=0;WeightsStore[2][202]<=0;WeightsStore[2][203]<=0;WeightsStore[2][204]<=0;WeightsStore[2][205]<=0;WeightsStore[2][206]<=0;WeightsStore[2][207]<=0;WeightsStore[2][208]<=0;WeightsStore[2][209]<=0;WeightsStore[2][210]<=0;WeightsStore[2][211]<=0;WeightsStore[2][212]<=0;WeightsStore[2][213]<=0;WeightsStore[2][214]<=0;WeightsStore[2][215]<=0;WeightsStore[2][216]<=0;WeightsStore[2][217]<=0;WeightsStore[2][218]<=0;WeightsStore[2][219]<=0;WeightsStore[2][220]<=0;WeightsStore[2][221]<=0;WeightsStore[2][222]<=0;WeightsStore[2][223]<=0;WeightsStore[2][224]<=0;WeightsStore[2][225]<=0;WeightsStore[2][226]<=0;WeightsStore[2][227]<=0;WeightsStore[2][228]<=0;WeightsStore[2][229]<=0;WeightsStore[2][230]<=0;WeightsStore[2][231]<=0;WeightsStore[2][232]<=0;WeightsStore[2][233]<=0;WeightsStore[2][234]<=0;WeightsStore[2][235]<=0;WeightsStore[2][236]<=0;WeightsStore[2][237]<=0;WeightsStore[2][238]<=0;WeightsStore[2][239]<=0;WeightsStore[2][240]<=0;WeightsStore[2][241]<=0;WeightsStore[2][242]<=0;WeightsStore[2][243]<=0;WeightsStore[2][244]<=0;WeightsStore[2][245]<=0;WeightsStore[2][246]<=0;WeightsStore[2][247]<=0;WeightsStore[2][248]<=0;WeightsStore[2][249]<=0;WeightsStore[2][250]<=0;WeightsStore[2][251]<=0;WeightsStore[2][252]<=0;WeightsStore[2][253]<=0;WeightsStore[2][254]<=0;WeightsStore[2][255]<=0;WeightsStore[2][256]<=0;WeightsStore[2][257]<=0;WeightsStore[2][258]<=0;WeightsStore[2][259]<=0;WeightsStore[2][260]<=0;WeightsStore[2][261]<=0;WeightsStore[2][262]<=0;WeightsStore[2][263]<=0;WeightsStore[2][264]<=0;WeightsStore[2][265]<=0;WeightsStore[2][266]<=0;WeightsStore[2][267]<=0;WeightsStore[2][268]<=0;WeightsStore[2][269]<=0;WeightsStore[2][270]<=0;WeightsStore[2][271]<=0;WeightsStore[2][272]<=0;WeightsStore[2][273]<=0;WeightsStore[2][274]<=0;WeightsStore[2][275]<=0;WeightsStore[2][276]<=0;WeightsStore[2][277]<=0;WeightsStore[2][278]<=0;WeightsStore[2][279]<=0;WeightsStore[2][280]<=0;WeightsStore[2][281]<=0;WeightsStore[2][282]<=0;WeightsStore[2][283]<=0;WeightsStore[2][284]<=0;WeightsStore[2][285]<=0;WeightsStore[2][286]<=0;WeightsStore[2][287]<=0;WeightsStore[2][288]<=0;WeightsStore[2][289]<=0;WeightsStore[2][290]<=0;WeightsStore[2][291]<=0;WeightsStore[2][292]<=0;WeightsStore[2][293]<=0;WeightsStore[2][294]<=0;WeightsStore[2][295]<=0;WeightsStore[2][296]<=0;WeightsStore[2][297]<=0;WeightsStore[2][298]<=0;WeightsStore[2][299]<=0;WeightsStore[2][300]<=0;WeightsStore[2][301]<=0;WeightsStore[2][302]<=0;WeightsStore[2][303]<=0;WeightsStore[2][304]<=0;WeightsStore[2][305]<=0;WeightsStore[2][306]<=0;WeightsStore[2][307]<=0;WeightsStore[2][308]<=0;WeightsStore[2][309]<=0;WeightsStore[2][310]<=0;WeightsStore[2][311]<=0;WeightsStore[2][312]<=0;WeightsStore[2][313]<=0;WeightsStore[2][314]<=0;WeightsStore[2][315]<=0;WeightsStore[2][316]<=0;WeightsStore[2][317]<=0;WeightsStore[2][318]<=0;WeightsStore[2][319]<=0;WeightsStore[2][320]<=0;WeightsStore[2][321]<=0;WeightsStore[2][322]<=0;WeightsStore[2][323]<=0;WeightsStore[2][324]<=0;WeightsStore[2][325]<=0;WeightsStore[2][326]<=0;WeightsStore[2][327]<=0;WeightsStore[2][328]<=0;WeightsStore[2][329]<=0;WeightsStore[2][330]<=0;WeightsStore[2][331]<=0;WeightsStore[2][332]<=0;WeightsStore[2][333]<=0;WeightsStore[2][334]<=0;WeightsStore[2][335]<=0;WeightsStore[2][336]<=0;WeightsStore[2][337]<=0;WeightsStore[2][338]<=0;WeightsStore[2][339]<=0;WeightsStore[2][340]<=0;WeightsStore[2][341]<=0;WeightsStore[2][342]<=0;WeightsStore[2][343]<=0;WeightsStore[2][344]<=0;WeightsStore[2][345]<=0;WeightsStore[2][346]<=0;WeightsStore[2][347]<=0;WeightsStore[2][348]<=0;WeightsStore[2][349]<=0;WeightsStore[2][350]<=0;WeightsStore[2][351]<=0;WeightsStore[2][352]<=0;WeightsStore[2][353]<=0;WeightsStore[2][354]<=0;WeightsStore[2][355]<=0;WeightsStore[2][356]<=0;WeightsStore[2][357]<=0;WeightsStore[2][358]<=0;WeightsStore[2][359]<=0;WeightsStore[2][360]<=0;WeightsStore[2][361]<=0;WeightsStore[2][362]<=0;WeightsStore[2][363]<=0;WeightsStore[2][364]<=0;WeightsStore[2][365]<=0;WeightsStore[2][366]<=0;WeightsStore[2][367]<=0;WeightsStore[2][368]<=0;WeightsStore[2][369]<=0;WeightsStore[2][370]<=0;WeightsStore[2][371]<=0;WeightsStore[2][372]<=0;WeightsStore[2][373]<=0;WeightsStore[2][374]<=0;WeightsStore[2][375]<=0;WeightsStore[2][376]<=0;WeightsStore[2][377]<=0;WeightsStore[2][378]<=0;WeightsStore[2][379]<=0;WeightsStore[2][380]<=0;WeightsStore[2][381]<=0;WeightsStore[2][382]<=0;WeightsStore[2][383]<=0;WeightsStore[2][384]<=0;WeightsStore[2][385]<=0;WeightsStore[2][386]<=0;WeightsStore[2][387]<=0;WeightsStore[2][388]<=0;WeightsStore[2][389]<=0;WeightsStore[2][390]<=0;WeightsStore[2][391]<=0;WeightsStore[2][392]<=0;WeightsStore[2][393]<=0;WeightsStore[2][394]<=0;WeightsStore[2][395]<=0;WeightsStore[2][396]<=0;WeightsStore[2][397]<=0;WeightsStore[2][398]<=0;WeightsStore[2][399]<=0;WeightsStore[2][400]<=0;WeightsStore[2][401]<=0;WeightsStore[2][402]<=0;WeightsStore[2][403]<=0;WeightsStore[2][404]<=0;WeightsStore[2][405]<=0;WeightsStore[2][406]<=0;WeightsStore[2][407]<=0;WeightsStore[2][408]<=0;WeightsStore[2][409]<=0;WeightsStore[2][410]<=0;WeightsStore[2][411]<=0;WeightsStore[2][412]<=0;WeightsStore[2][413]<=0;WeightsStore[2][414]<=0;WeightsStore[2][415]<=0;WeightsStore[2][416]<=0;WeightsStore[2][417]<=0;WeightsStore[2][418]<=0;WeightsStore[2][419]<=0;WeightsStore[2][420]<=0;WeightsStore[2][421]<=0;WeightsStore[2][422]<=0;WeightsStore[2][423]<=0;WeightsStore[2][424]<=0;WeightsStore[2][425]<=0;WeightsStore[2][426]<=0;WeightsStore[2][427]<=0;WeightsStore[2][428]<=0;WeightsStore[2][429]<=0;WeightsStore[2][430]<=0;WeightsStore[2][431]<=0;WeightsStore[2][432]<=0;WeightsStore[2][433]<=0;WeightsStore[2][434]<=0;WeightsStore[2][435]<=0;WeightsStore[2][436]<=0;WeightsStore[2][437]<=0;WeightsStore[2][438]<=0;WeightsStore[2][439]<=0;WeightsStore[2][440]<=0;WeightsStore[2][441]<=0;WeightsStore[2][442]<=0;WeightsStore[2][443]<=0;WeightsStore[2][444]<=0;WeightsStore[2][445]<=0;WeightsStore[2][446]<=0;WeightsStore[2][447]<=0;WeightsStore[2][448]<=0;WeightsStore[2][449]<=0;WeightsStore[2][450]<=0;WeightsStore[2][451]<=0;WeightsStore[2][452]<=0;WeightsStore[2][453]<=0;WeightsStore[2][454]<=0;WeightsStore[2][455]<=0;WeightsStore[2][456]<=0;WeightsStore[2][457]<=0;WeightsStore[2][458]<=0;WeightsStore[2][459]<=0;WeightsStore[2][460]<=0;WeightsStore[2][461]<=0;WeightsStore[2][462]<=0;WeightsStore[2][463]<=0;WeightsStore[2][464]<=0;WeightsStore[2][465]<=0;WeightsStore[2][466]<=0;WeightsStore[2][467]<=0;WeightsStore[2][468]<=0;WeightsStore[2][469]<=0;WeightsStore[2][470]<=0;WeightsStore[2][471]<=0;WeightsStore[2][472]<=0;WeightsStore[2][473]<=0;WeightsStore[2][474]<=0;WeightsStore[2][475]<=0;WeightsStore[2][476]<=0;WeightsStore[2][477]<=0;WeightsStore[2][478]<=0;WeightsStore[2][479]<=0;WeightsStore[2][480]<=0;WeightsStore[2][481]<=0;WeightsStore[2][482]<=0;WeightsStore[2][483]<=0;WeightsStore[2][484]<=0;WeightsStore[2][485]<=0;WeightsStore[2][486]<=0;WeightsStore[2][487]<=0;WeightsStore[2][488]<=0;WeightsStore[2][489]<=0;WeightsStore[2][490]<=0;WeightsStore[2][491]<=0;WeightsStore[2][492]<=0;WeightsStore[2][493]<=0;WeightsStore[2][494]<=0;WeightsStore[2][495]<=0;WeightsStore[2][496]<=0;WeightsStore[2][497]<=0;WeightsStore[2][498]<=0;WeightsStore[2][499]<=0;WeightsStore[2][500]<=0;WeightsStore[2][501]<=0;WeightsStore[2][502]<=0;WeightsStore[2][503]<=0;WeightsStore[2][504]<=0;WeightsStore[2][505]<=0;WeightsStore[2][506]<=0;WeightsStore[2][507]<=0;WeightsStore[2][508]<=0;WeightsStore[2][509]<=0;WeightsStore[2][510]<=0;WeightsStore[2][511]<=0;WeightsStore[2][512]<=0;WeightsStore[2][513]<=0;WeightsStore[2][514]<=0;WeightsStore[2][515]<=0;WeightsStore[2][516]<=0;WeightsStore[2][517]<=0;WeightsStore[2][518]<=0;WeightsStore[2][519]<=0;WeightsStore[2][520]<=0;WeightsStore[2][521]<=0;WeightsStore[2][522]<=0;WeightsStore[2][523]<=0;WeightsStore[2][524]<=0;WeightsStore[2][525]<=0;WeightsStore[2][526]<=0;WeightsStore[2][527]<=0;WeightsStore[2][528]<=0;WeightsStore[2][529]<=0;WeightsStore[2][530]<=0;WeightsStore[2][531]<=0;WeightsStore[2][532]<=0;WeightsStore[2][533]<=0;WeightsStore[2][534]<=0;WeightsStore[2][535]<=0;WeightsStore[2][536]<=0;WeightsStore[2][537]<=0;WeightsStore[2][538]<=0;WeightsStore[2][539]<=0;WeightsStore[2][540]<=0;WeightsStore[2][541]<=0;WeightsStore[2][542]<=0;WeightsStore[2][543]<=0;WeightsStore[2][544]<=0;WeightsStore[2][545]<=0;WeightsStore[2][546]<=0;WeightsStore[2][547]<=0;WeightsStore[2][548]<=0;WeightsStore[2][549]<=0;WeightsStore[2][550]<=0;WeightsStore[2][551]<=0;WeightsStore[2][552]<=0;WeightsStore[2][553]<=0;WeightsStore[2][554]<=0;WeightsStore[2][555]<=0;WeightsStore[2][556]<=0;WeightsStore[2][557]<=0;WeightsStore[2][558]<=0;WeightsStore[2][559]<=0;WeightsStore[2][560]<=0;WeightsStore[2][561]<=0;WeightsStore[2][562]<=0;WeightsStore[2][563]<=0;WeightsStore[2][564]<=0;WeightsStore[2][565]<=0;WeightsStore[2][566]<=0;WeightsStore[2][567]<=0;WeightsStore[2][568]<=0;WeightsStore[2][569]<=0;WeightsStore[2][570]<=0;WeightsStore[2][571]<=0;WeightsStore[2][572]<=0;WeightsStore[2][573]<=0;WeightsStore[2][574]<=0;WeightsStore[2][575]<=0;WeightsStore[2][576]<=0;WeightsStore[2][577]<=0;WeightsStore[2][578]<=0;WeightsStore[2][579]<=0;WeightsStore[2][580]<=0;WeightsStore[2][581]<=0;WeightsStore[2][582]<=0;WeightsStore[2][583]<=0;WeightsStore[2][584]<=0;WeightsStore[2][585]<=0;WeightsStore[2][586]<=0;WeightsStore[2][587]<=0;WeightsStore[2][588]<=0;WeightsStore[2][589]<=0;WeightsStore[2][590]<=0;WeightsStore[2][591]<=0;WeightsStore[2][592]<=0;WeightsStore[2][593]<=0;WeightsStore[2][594]<=0;WeightsStore[2][595]<=0;WeightsStore[2][596]<=0;WeightsStore[2][597]<=0;WeightsStore[2][598]<=0;WeightsStore[2][599]<=0;WeightsStore[2][600]<=0;WeightsStore[2][601]<=0;WeightsStore[2][602]<=0;WeightsStore[2][603]<=0;WeightsStore[2][604]<=0;WeightsStore[2][605]<=0;WeightsStore[2][606]<=0;WeightsStore[2][607]<=0;WeightsStore[2][608]<=0;WeightsStore[2][609]<=0;WeightsStore[2][610]<=0;WeightsStore[2][611]<=0;WeightsStore[2][612]<=0;WeightsStore[2][613]<=0;WeightsStore[2][614]<=0;WeightsStore[2][615]<=0;WeightsStore[2][616]<=0;WeightsStore[2][617]<=0;WeightsStore[2][618]<=0;WeightsStore[2][619]<=0;WeightsStore[2][620]<=0;WeightsStore[2][621]<=0;WeightsStore[2][622]<=0;WeightsStore[2][623]<=0;WeightsStore[2][624]<=0;WeightsStore[2][625]<=0;WeightsStore[2][626]<=0;WeightsStore[2][627]<=0;WeightsStore[2][628]<=0;WeightsStore[2][629]<=0;WeightsStore[2][630]<=0;WeightsStore[2][631]<=0;WeightsStore[2][632]<=0;WeightsStore[2][633]<=0;WeightsStore[2][634]<=0;WeightsStore[2][635]<=0;WeightsStore[2][636]<=0;WeightsStore[2][637]<=0;WeightsStore[2][638]<=0;WeightsStore[2][639]<=0;WeightsStore[2][640]<=0;WeightsStore[2][641]<=0;WeightsStore[2][642]<=0;WeightsStore[2][643]<=0;WeightsStore[2][644]<=0;WeightsStore[2][645]<=0;WeightsStore[2][646]<=0;WeightsStore[2][647]<=0;WeightsStore[2][648]<=0;WeightsStore[2][649]<=0;WeightsStore[2][650]<=0;WeightsStore[2][651]<=0;WeightsStore[2][652]<=0;WeightsStore[2][653]<=0;WeightsStore[2][654]<=0;WeightsStore[2][655]<=0;WeightsStore[2][656]<=0;WeightsStore[2][657]<=0;WeightsStore[2][658]<=0;WeightsStore[2][659]<=0;WeightsStore[2][660]<=0;WeightsStore[2][661]<=0;WeightsStore[2][662]<=0;WeightsStore[2][663]<=0;WeightsStore[2][664]<=0;WeightsStore[2][665]<=0;WeightsStore[2][666]<=0;WeightsStore[2][667]<=0;WeightsStore[2][668]<=0;WeightsStore[2][669]<=0;WeightsStore[2][670]<=0;WeightsStore[2][671]<=0;WeightsStore[2][672]<=0;WeightsStore[2][673]<=0;WeightsStore[2][674]<=0;WeightsStore[2][675]<=0;WeightsStore[2][676]<=0;WeightsStore[2][677]<=0;WeightsStore[2][678]<=0;WeightsStore[2][679]<=0;WeightsStore[2][680]<=0;WeightsStore[2][681]<=0;WeightsStore[2][682]<=0;WeightsStore[2][683]<=0;WeightsStore[2][684]<=0;WeightsStore[2][685]<=0;WeightsStore[2][686]<=0;WeightsStore[2][687]<=0;WeightsStore[2][688]<=0;WeightsStore[2][689]<=0;WeightsStore[2][690]<=0;WeightsStore[2][691]<=0;WeightsStore[2][692]<=0;WeightsStore[2][693]<=0;WeightsStore[2][694]<=0;WeightsStore[2][695]<=0;WeightsStore[2][696]<=0;WeightsStore[2][697]<=0;WeightsStore[2][698]<=0;WeightsStore[2][699]<=0;WeightsStore[2][700]<=0;WeightsStore[2][701]<=0;WeightsStore[2][702]<=0;WeightsStore[2][703]<=0;WeightsStore[2][704]<=0;WeightsStore[2][705]<=0;WeightsStore[2][706]<=0;WeightsStore[2][707]<=0;WeightsStore[2][708]<=0;WeightsStore[2][709]<=0;WeightsStore[2][710]<=0;WeightsStore[2][711]<=0;WeightsStore[2][712]<=0;WeightsStore[2][713]<=0;WeightsStore[2][714]<=0;WeightsStore[2][715]<=0;WeightsStore[2][716]<=0;WeightsStore[2][717]<=0;WeightsStore[2][718]<=0;WeightsStore[2][719]<=0;WeightsStore[2][720]<=0;WeightsStore[2][721]<=0;WeightsStore[2][722]<=0;WeightsStore[2][723]<=0;WeightsStore[2][724]<=0;WeightsStore[2][725]<=0;WeightsStore[2][726]<=0;WeightsStore[2][727]<=0;WeightsStore[2][728]<=0;WeightsStore[2][729]<=0;WeightsStore[2][730]<=0;WeightsStore[2][731]<=0;WeightsStore[2][732]<=0;WeightsStore[2][733]<=0;WeightsStore[2][734]<=0;WeightsStore[2][735]<=0;WeightsStore[2][736]<=0;WeightsStore[2][737]<=0;WeightsStore[2][738]<=0;WeightsStore[2][739]<=0;WeightsStore[2][740]<=0;WeightsStore[2][741]<=0;WeightsStore[2][742]<=0;WeightsStore[2][743]<=0;WeightsStore[2][744]<=0;WeightsStore[2][745]<=0;WeightsStore[2][746]<=0;WeightsStore[2][747]<=0;WeightsStore[2][748]<=0;WeightsStore[2][749]<=0;WeightsStore[2][750]<=0;WeightsStore[2][751]<=0;WeightsStore[2][752]<=0;WeightsStore[2][753]<=0;WeightsStore[2][754]<=0;WeightsStore[2][755]<=0;WeightsStore[2][756]<=0;WeightsStore[2][757]<=0;WeightsStore[2][758]<=0;WeightsStore[2][759]<=0;WeightsStore[2][760]<=0;WeightsStore[2][761]<=0;WeightsStore[2][762]<=0;WeightsStore[2][763]<=0;WeightsStore[2][764]<=0;WeightsStore[2][765]<=0;WeightsStore[2][766]<=0;WeightsStore[2][767]<=0;WeightsStore[2][768]<=0;WeightsStore[2][769]<=0;WeightsStore[2][770]<=0;WeightsStore[2][771]<=0;WeightsStore[2][772]<=0;WeightsStore[2][773]<=0;WeightsStore[2][774]<=0;WeightsStore[2][775]<=0;WeightsStore[2][776]<=0;WeightsStore[2][777]<=0;WeightsStore[2][778]<=0;WeightsStore[2][779]<=0;WeightsStore[2][780]<=0;WeightsStore[2][781]<=0;WeightsStore[2][782]<=0;WeightsStore[2][783]<=0;WeightsStore[2][784]<=0;WeightsStore[3][0]<=0;WeightsStore[3][1]<=0;WeightsStore[3][2]<=0;WeightsStore[3][3]<=0;WeightsStore[3][4]<=0;WeightsStore[3][5]<=0;WeightsStore[3][6]<=0;WeightsStore[3][7]<=0;WeightsStore[3][8]<=0;WeightsStore[3][9]<=0;WeightsStore[3][10]<=0;WeightsStore[3][11]<=0;WeightsStore[3][12]<=0;WeightsStore[3][13]<=0;WeightsStore[3][14]<=0;WeightsStore[3][15]<=0;WeightsStore[3][16]<=0;WeightsStore[3][17]<=0;WeightsStore[3][18]<=0;WeightsStore[3][19]<=0;WeightsStore[3][20]<=0;WeightsStore[3][21]<=0;WeightsStore[3][22]<=0;WeightsStore[3][23]<=0;WeightsStore[3][24]<=0;WeightsStore[3][25]<=0;WeightsStore[3][26]<=0;WeightsStore[3][27]<=0;WeightsStore[3][28]<=0;WeightsStore[3][29]<=0;WeightsStore[3][30]<=0;WeightsStore[3][31]<=0;WeightsStore[3][32]<=0;WeightsStore[3][33]<=0;WeightsStore[3][34]<=0;WeightsStore[3][35]<=0;WeightsStore[3][36]<=0;WeightsStore[3][37]<=0;WeightsStore[3][38]<=0;WeightsStore[3][39]<=0;WeightsStore[3][40]<=0;WeightsStore[3][41]<=0;WeightsStore[3][42]<=0;WeightsStore[3][43]<=0;WeightsStore[3][44]<=0;WeightsStore[3][45]<=0;WeightsStore[3][46]<=0;WeightsStore[3][47]<=0;WeightsStore[3][48]<=0;WeightsStore[3][49]<=0;WeightsStore[3][50]<=0;WeightsStore[3][51]<=0;WeightsStore[3][52]<=0;WeightsStore[3][53]<=0;WeightsStore[3][54]<=0;WeightsStore[3][55]<=0;WeightsStore[3][56]<=0;WeightsStore[3][57]<=0;WeightsStore[3][58]<=0;WeightsStore[3][59]<=0;WeightsStore[3][60]<=0;WeightsStore[3][61]<=0;WeightsStore[3][62]<=0;WeightsStore[3][63]<=0;WeightsStore[3][64]<=0;WeightsStore[3][65]<=0;WeightsStore[3][66]<=0;WeightsStore[3][67]<=0;WeightsStore[3][68]<=0;WeightsStore[3][69]<=0;WeightsStore[3][70]<=0;WeightsStore[3][71]<=0;WeightsStore[3][72]<=0;WeightsStore[3][73]<=0;WeightsStore[3][74]<=0;WeightsStore[3][75]<=0;WeightsStore[3][76]<=0;WeightsStore[3][77]<=0;WeightsStore[3][78]<=0;WeightsStore[3][79]<=0;WeightsStore[3][80]<=0;WeightsStore[3][81]<=0;WeightsStore[3][82]<=0;WeightsStore[3][83]<=0;WeightsStore[3][84]<=0;WeightsStore[3][85]<=0;WeightsStore[3][86]<=0;WeightsStore[3][87]<=0;WeightsStore[3][88]<=0;WeightsStore[3][89]<=0;WeightsStore[3][90]<=0;WeightsStore[3][91]<=0;WeightsStore[3][92]<=0;WeightsStore[3][93]<=0;WeightsStore[3][94]<=0;WeightsStore[3][95]<=0;WeightsStore[3][96]<=0;WeightsStore[3][97]<=0;WeightsStore[3][98]<=0;WeightsStore[3][99]<=0;WeightsStore[3][100]<=0;WeightsStore[3][101]<=0;WeightsStore[3][102]<=0;WeightsStore[3][103]<=0;WeightsStore[3][104]<=0;WeightsStore[3][105]<=0;WeightsStore[3][106]<=0;WeightsStore[3][107]<=0;WeightsStore[3][108]<=0;WeightsStore[3][109]<=0;WeightsStore[3][110]<=0;WeightsStore[3][111]<=0;WeightsStore[3][112]<=0;WeightsStore[3][113]<=0;WeightsStore[3][114]<=0;WeightsStore[3][115]<=0;WeightsStore[3][116]<=0;WeightsStore[3][117]<=0;WeightsStore[3][118]<=0;WeightsStore[3][119]<=0;WeightsStore[3][120]<=0;WeightsStore[3][121]<=0;WeightsStore[3][122]<=0;WeightsStore[3][123]<=0;WeightsStore[3][124]<=0;WeightsStore[3][125]<=0;WeightsStore[3][126]<=0;WeightsStore[3][127]<=0;WeightsStore[3][128]<=0;WeightsStore[3][129]<=0;WeightsStore[3][130]<=0;WeightsStore[3][131]<=0;WeightsStore[3][132]<=0;WeightsStore[3][133]<=0;WeightsStore[3][134]<=0;WeightsStore[3][135]<=0;WeightsStore[3][136]<=0;WeightsStore[3][137]<=0;WeightsStore[3][138]<=0;WeightsStore[3][139]<=0;WeightsStore[3][140]<=0;WeightsStore[3][141]<=0;WeightsStore[3][142]<=0;WeightsStore[3][143]<=0;WeightsStore[3][144]<=0;WeightsStore[3][145]<=0;WeightsStore[3][146]<=0;WeightsStore[3][147]<=0;WeightsStore[3][148]<=0;WeightsStore[3][149]<=0;WeightsStore[3][150]<=0;WeightsStore[3][151]<=0;WeightsStore[3][152]<=0;WeightsStore[3][153]<=0;WeightsStore[3][154]<=0;WeightsStore[3][155]<=0;WeightsStore[3][156]<=0;WeightsStore[3][157]<=0;WeightsStore[3][158]<=0;WeightsStore[3][159]<=0;WeightsStore[3][160]<=0;WeightsStore[3][161]<=0;WeightsStore[3][162]<=0;WeightsStore[3][163]<=0;WeightsStore[3][164]<=0;WeightsStore[3][165]<=0;WeightsStore[3][166]<=0;WeightsStore[3][167]<=0;WeightsStore[3][168]<=0;WeightsStore[3][169]<=0;WeightsStore[3][170]<=0;WeightsStore[3][171]<=0;WeightsStore[3][172]<=0;WeightsStore[3][173]<=0;WeightsStore[3][174]<=0;WeightsStore[3][175]<=0;WeightsStore[3][176]<=0;WeightsStore[3][177]<=0;WeightsStore[3][178]<=0;WeightsStore[3][179]<=0;WeightsStore[3][180]<=0;WeightsStore[3][181]<=0;WeightsStore[3][182]<=0;WeightsStore[3][183]<=0;WeightsStore[3][184]<=0;WeightsStore[3][185]<=0;WeightsStore[3][186]<=0;WeightsStore[3][187]<=0;WeightsStore[3][188]<=0;WeightsStore[3][189]<=0;WeightsStore[3][190]<=0;WeightsStore[3][191]<=0;WeightsStore[3][192]<=0;WeightsStore[3][193]<=0;WeightsStore[3][194]<=0;WeightsStore[3][195]<=0;WeightsStore[3][196]<=0;WeightsStore[3][197]<=0;WeightsStore[3][198]<=0;WeightsStore[3][199]<=0;WeightsStore[3][200]<=0;WeightsStore[3][201]<=0;WeightsStore[3][202]<=0;WeightsStore[3][203]<=0;WeightsStore[3][204]<=0;WeightsStore[3][205]<=0;WeightsStore[3][206]<=0;WeightsStore[3][207]<=0;WeightsStore[3][208]<=0;WeightsStore[3][209]<=0;WeightsStore[3][210]<=0;WeightsStore[3][211]<=0;WeightsStore[3][212]<=0;WeightsStore[3][213]<=0;WeightsStore[3][214]<=0;WeightsStore[3][215]<=0;WeightsStore[3][216]<=0;WeightsStore[3][217]<=0;WeightsStore[3][218]<=0;WeightsStore[3][219]<=0;WeightsStore[3][220]<=0;WeightsStore[3][221]<=0;WeightsStore[3][222]<=0;WeightsStore[3][223]<=0;WeightsStore[3][224]<=0;WeightsStore[3][225]<=0;WeightsStore[3][226]<=0;WeightsStore[3][227]<=0;WeightsStore[3][228]<=0;WeightsStore[3][229]<=0;WeightsStore[3][230]<=0;WeightsStore[3][231]<=0;WeightsStore[3][232]<=0;WeightsStore[3][233]<=0;WeightsStore[3][234]<=0;WeightsStore[3][235]<=0;WeightsStore[3][236]<=0;WeightsStore[3][237]<=0;WeightsStore[3][238]<=0;WeightsStore[3][239]<=0;WeightsStore[3][240]<=0;WeightsStore[3][241]<=0;WeightsStore[3][242]<=0;WeightsStore[3][243]<=0;WeightsStore[3][244]<=0;WeightsStore[3][245]<=0;WeightsStore[3][246]<=0;WeightsStore[3][247]<=0;WeightsStore[3][248]<=0;WeightsStore[3][249]<=0;WeightsStore[3][250]<=0;WeightsStore[3][251]<=0;WeightsStore[3][252]<=0;WeightsStore[3][253]<=0;WeightsStore[3][254]<=0;WeightsStore[3][255]<=0;WeightsStore[3][256]<=0;WeightsStore[3][257]<=0;WeightsStore[3][258]<=0;WeightsStore[3][259]<=0;WeightsStore[3][260]<=0;WeightsStore[3][261]<=0;WeightsStore[3][262]<=0;WeightsStore[3][263]<=0;WeightsStore[3][264]<=0;WeightsStore[3][265]<=0;WeightsStore[3][266]<=0;WeightsStore[3][267]<=0;WeightsStore[3][268]<=0;WeightsStore[3][269]<=0;WeightsStore[3][270]<=0;WeightsStore[3][271]<=0;WeightsStore[3][272]<=0;WeightsStore[3][273]<=0;WeightsStore[3][274]<=0;WeightsStore[3][275]<=0;WeightsStore[3][276]<=0;WeightsStore[3][277]<=0;WeightsStore[3][278]<=0;WeightsStore[3][279]<=0;WeightsStore[3][280]<=0;WeightsStore[3][281]<=0;WeightsStore[3][282]<=0;WeightsStore[3][283]<=0;WeightsStore[3][284]<=0;WeightsStore[3][285]<=0;WeightsStore[3][286]<=0;WeightsStore[3][287]<=0;WeightsStore[3][288]<=0;WeightsStore[3][289]<=0;WeightsStore[3][290]<=0;WeightsStore[3][291]<=0;WeightsStore[3][292]<=0;WeightsStore[3][293]<=0;WeightsStore[3][294]<=0;WeightsStore[3][295]<=0;WeightsStore[3][296]<=0;WeightsStore[3][297]<=0;WeightsStore[3][298]<=0;WeightsStore[3][299]<=0;WeightsStore[3][300]<=0;WeightsStore[3][301]<=0;WeightsStore[3][302]<=0;WeightsStore[3][303]<=0;WeightsStore[3][304]<=0;WeightsStore[3][305]<=0;WeightsStore[3][306]<=0;WeightsStore[3][307]<=0;WeightsStore[3][308]<=0;WeightsStore[3][309]<=0;WeightsStore[3][310]<=0;WeightsStore[3][311]<=0;WeightsStore[3][312]<=0;WeightsStore[3][313]<=0;WeightsStore[3][314]<=0;WeightsStore[3][315]<=0;WeightsStore[3][316]<=0;WeightsStore[3][317]<=0;WeightsStore[3][318]<=0;WeightsStore[3][319]<=0;WeightsStore[3][320]<=0;WeightsStore[3][321]<=0;WeightsStore[3][322]<=0;WeightsStore[3][323]<=0;WeightsStore[3][324]<=0;WeightsStore[3][325]<=0;WeightsStore[3][326]<=0;WeightsStore[3][327]<=0;WeightsStore[3][328]<=0;WeightsStore[3][329]<=0;WeightsStore[3][330]<=0;WeightsStore[3][331]<=0;WeightsStore[3][332]<=0;WeightsStore[3][333]<=0;WeightsStore[3][334]<=0;WeightsStore[3][335]<=0;WeightsStore[3][336]<=0;WeightsStore[3][337]<=0;WeightsStore[3][338]<=0;WeightsStore[3][339]<=0;WeightsStore[3][340]<=0;WeightsStore[3][341]<=0;WeightsStore[3][342]<=0;WeightsStore[3][343]<=0;WeightsStore[3][344]<=0;WeightsStore[3][345]<=0;WeightsStore[3][346]<=0;WeightsStore[3][347]<=0;WeightsStore[3][348]<=0;WeightsStore[3][349]<=0;WeightsStore[3][350]<=0;WeightsStore[3][351]<=0;WeightsStore[3][352]<=0;WeightsStore[3][353]<=0;WeightsStore[3][354]<=0;WeightsStore[3][355]<=0;WeightsStore[3][356]<=0;WeightsStore[3][357]<=0;WeightsStore[3][358]<=0;WeightsStore[3][359]<=0;WeightsStore[3][360]<=0;WeightsStore[3][361]<=0;WeightsStore[3][362]<=0;WeightsStore[3][363]<=0;WeightsStore[3][364]<=0;WeightsStore[3][365]<=0;WeightsStore[3][366]<=0;WeightsStore[3][367]<=0;WeightsStore[3][368]<=0;WeightsStore[3][369]<=0;WeightsStore[3][370]<=0;WeightsStore[3][371]<=0;WeightsStore[3][372]<=0;WeightsStore[3][373]<=0;WeightsStore[3][374]<=0;WeightsStore[3][375]<=0;WeightsStore[3][376]<=0;WeightsStore[3][377]<=0;WeightsStore[3][378]<=0;WeightsStore[3][379]<=0;WeightsStore[3][380]<=0;WeightsStore[3][381]<=0;WeightsStore[3][382]<=0;WeightsStore[3][383]<=0;WeightsStore[3][384]<=0;WeightsStore[3][385]<=0;WeightsStore[3][386]<=0;WeightsStore[3][387]<=0;WeightsStore[3][388]<=0;WeightsStore[3][389]<=0;WeightsStore[3][390]<=0;WeightsStore[3][391]<=0;WeightsStore[3][392]<=0;WeightsStore[3][393]<=0;WeightsStore[3][394]<=0;WeightsStore[3][395]<=0;WeightsStore[3][396]<=0;WeightsStore[3][397]<=0;WeightsStore[3][398]<=0;WeightsStore[3][399]<=0;WeightsStore[3][400]<=0;WeightsStore[3][401]<=0;WeightsStore[3][402]<=0;WeightsStore[3][403]<=0;WeightsStore[3][404]<=0;WeightsStore[3][405]<=0;WeightsStore[3][406]<=0;WeightsStore[3][407]<=0;WeightsStore[3][408]<=0;WeightsStore[3][409]<=0;WeightsStore[3][410]<=0;WeightsStore[3][411]<=0;WeightsStore[3][412]<=0;WeightsStore[3][413]<=0;WeightsStore[3][414]<=0;WeightsStore[3][415]<=0;WeightsStore[3][416]<=0;WeightsStore[3][417]<=0;WeightsStore[3][418]<=0;WeightsStore[3][419]<=0;WeightsStore[3][420]<=0;WeightsStore[3][421]<=0;WeightsStore[3][422]<=0;WeightsStore[3][423]<=0;WeightsStore[3][424]<=0;WeightsStore[3][425]<=0;WeightsStore[3][426]<=0;WeightsStore[3][427]<=0;WeightsStore[3][428]<=0;WeightsStore[3][429]<=0;WeightsStore[3][430]<=0;WeightsStore[3][431]<=0;WeightsStore[3][432]<=0;WeightsStore[3][433]<=0;WeightsStore[3][434]<=0;WeightsStore[3][435]<=0;WeightsStore[3][436]<=0;WeightsStore[3][437]<=0;WeightsStore[3][438]<=0;WeightsStore[3][439]<=0;WeightsStore[3][440]<=0;WeightsStore[3][441]<=0;WeightsStore[3][442]<=0;WeightsStore[3][443]<=0;WeightsStore[3][444]<=0;WeightsStore[3][445]<=0;WeightsStore[3][446]<=0;WeightsStore[3][447]<=0;WeightsStore[3][448]<=0;WeightsStore[3][449]<=0;WeightsStore[3][450]<=0;WeightsStore[3][451]<=0;WeightsStore[3][452]<=0;WeightsStore[3][453]<=0;WeightsStore[3][454]<=0;WeightsStore[3][455]<=0;WeightsStore[3][456]<=0;WeightsStore[3][457]<=0;WeightsStore[3][458]<=0;WeightsStore[3][459]<=0;WeightsStore[3][460]<=0;WeightsStore[3][461]<=0;WeightsStore[3][462]<=0;WeightsStore[3][463]<=0;WeightsStore[3][464]<=0;WeightsStore[3][465]<=0;WeightsStore[3][466]<=0;WeightsStore[3][467]<=0;WeightsStore[3][468]<=0;WeightsStore[3][469]<=0;WeightsStore[3][470]<=0;WeightsStore[3][471]<=0;WeightsStore[3][472]<=0;WeightsStore[3][473]<=0;WeightsStore[3][474]<=0;WeightsStore[3][475]<=0;WeightsStore[3][476]<=0;WeightsStore[3][477]<=0;WeightsStore[3][478]<=0;WeightsStore[3][479]<=0;WeightsStore[3][480]<=0;WeightsStore[3][481]<=0;WeightsStore[3][482]<=0;WeightsStore[3][483]<=0;WeightsStore[3][484]<=0;WeightsStore[3][485]<=0;WeightsStore[3][486]<=0;WeightsStore[3][487]<=0;WeightsStore[3][488]<=0;WeightsStore[3][489]<=0;WeightsStore[3][490]<=0;WeightsStore[3][491]<=0;WeightsStore[3][492]<=0;WeightsStore[3][493]<=0;WeightsStore[3][494]<=0;WeightsStore[3][495]<=0;WeightsStore[3][496]<=0;WeightsStore[3][497]<=0;WeightsStore[3][498]<=0;WeightsStore[3][499]<=0;WeightsStore[3][500]<=0;WeightsStore[3][501]<=0;WeightsStore[3][502]<=0;WeightsStore[3][503]<=0;WeightsStore[3][504]<=0;WeightsStore[3][505]<=0;WeightsStore[3][506]<=0;WeightsStore[3][507]<=0;WeightsStore[3][508]<=0;WeightsStore[3][509]<=0;WeightsStore[3][510]<=0;WeightsStore[3][511]<=0;WeightsStore[3][512]<=0;WeightsStore[3][513]<=0;WeightsStore[3][514]<=0;WeightsStore[3][515]<=0;WeightsStore[3][516]<=0;WeightsStore[3][517]<=0;WeightsStore[3][518]<=0;WeightsStore[3][519]<=0;WeightsStore[3][520]<=0;WeightsStore[3][521]<=0;WeightsStore[3][522]<=0;WeightsStore[3][523]<=0;WeightsStore[3][524]<=0;WeightsStore[3][525]<=0;WeightsStore[3][526]<=0;WeightsStore[3][527]<=0;WeightsStore[3][528]<=0;WeightsStore[3][529]<=0;WeightsStore[3][530]<=0;WeightsStore[3][531]<=0;WeightsStore[3][532]<=0;WeightsStore[3][533]<=0;WeightsStore[3][534]<=0;WeightsStore[3][535]<=0;WeightsStore[3][536]<=0;WeightsStore[3][537]<=0;WeightsStore[3][538]<=0;WeightsStore[3][539]<=0;WeightsStore[3][540]<=0;WeightsStore[3][541]<=0;WeightsStore[3][542]<=0;WeightsStore[3][543]<=0;WeightsStore[3][544]<=0;WeightsStore[3][545]<=0;WeightsStore[3][546]<=0;WeightsStore[3][547]<=0;WeightsStore[3][548]<=0;WeightsStore[3][549]<=0;WeightsStore[3][550]<=0;WeightsStore[3][551]<=0;WeightsStore[3][552]<=0;WeightsStore[3][553]<=0;WeightsStore[3][554]<=0;WeightsStore[3][555]<=0;WeightsStore[3][556]<=0;WeightsStore[3][557]<=0;WeightsStore[3][558]<=0;WeightsStore[3][559]<=0;WeightsStore[3][560]<=0;WeightsStore[3][561]<=0;WeightsStore[3][562]<=0;WeightsStore[3][563]<=0;WeightsStore[3][564]<=0;WeightsStore[3][565]<=0;WeightsStore[3][566]<=0;WeightsStore[3][567]<=0;WeightsStore[3][568]<=0;WeightsStore[3][569]<=0;WeightsStore[3][570]<=0;WeightsStore[3][571]<=0;WeightsStore[3][572]<=0;WeightsStore[3][573]<=0;WeightsStore[3][574]<=0;WeightsStore[3][575]<=0;WeightsStore[3][576]<=0;WeightsStore[3][577]<=0;WeightsStore[3][578]<=0;WeightsStore[3][579]<=0;WeightsStore[3][580]<=0;WeightsStore[3][581]<=0;WeightsStore[3][582]<=0;WeightsStore[3][583]<=0;WeightsStore[3][584]<=0;WeightsStore[3][585]<=0;WeightsStore[3][586]<=0;WeightsStore[3][587]<=0;WeightsStore[3][588]<=0;WeightsStore[3][589]<=0;WeightsStore[3][590]<=0;WeightsStore[3][591]<=0;WeightsStore[3][592]<=0;WeightsStore[3][593]<=0;WeightsStore[3][594]<=0;WeightsStore[3][595]<=0;WeightsStore[3][596]<=0;WeightsStore[3][597]<=0;WeightsStore[3][598]<=0;WeightsStore[3][599]<=0;WeightsStore[3][600]<=0;WeightsStore[3][601]<=0;WeightsStore[3][602]<=0;WeightsStore[3][603]<=0;WeightsStore[3][604]<=0;WeightsStore[3][605]<=0;WeightsStore[3][606]<=0;WeightsStore[3][607]<=0;WeightsStore[3][608]<=0;WeightsStore[3][609]<=0;WeightsStore[3][610]<=0;WeightsStore[3][611]<=0;WeightsStore[3][612]<=0;WeightsStore[3][613]<=0;WeightsStore[3][614]<=0;WeightsStore[3][615]<=0;WeightsStore[3][616]<=0;WeightsStore[3][617]<=0;WeightsStore[3][618]<=0;WeightsStore[3][619]<=0;WeightsStore[3][620]<=0;WeightsStore[3][621]<=0;WeightsStore[3][622]<=0;WeightsStore[3][623]<=0;WeightsStore[3][624]<=0;WeightsStore[3][625]<=0;WeightsStore[3][626]<=0;WeightsStore[3][627]<=0;WeightsStore[3][628]<=0;WeightsStore[3][629]<=0;WeightsStore[3][630]<=0;WeightsStore[3][631]<=0;WeightsStore[3][632]<=0;WeightsStore[3][633]<=0;WeightsStore[3][634]<=0;WeightsStore[3][635]<=0;WeightsStore[3][636]<=0;WeightsStore[3][637]<=0;WeightsStore[3][638]<=0;WeightsStore[3][639]<=0;WeightsStore[3][640]<=0;WeightsStore[3][641]<=0;WeightsStore[3][642]<=0;WeightsStore[3][643]<=0;WeightsStore[3][644]<=0;WeightsStore[3][645]<=0;WeightsStore[3][646]<=0;WeightsStore[3][647]<=0;WeightsStore[3][648]<=0;WeightsStore[3][649]<=0;WeightsStore[3][650]<=0;WeightsStore[3][651]<=0;WeightsStore[3][652]<=0;WeightsStore[3][653]<=0;WeightsStore[3][654]<=0;WeightsStore[3][655]<=0;WeightsStore[3][656]<=0;WeightsStore[3][657]<=0;WeightsStore[3][658]<=0;WeightsStore[3][659]<=0;WeightsStore[3][660]<=0;WeightsStore[3][661]<=0;WeightsStore[3][662]<=0;WeightsStore[3][663]<=0;WeightsStore[3][664]<=0;WeightsStore[3][665]<=0;WeightsStore[3][666]<=0;WeightsStore[3][667]<=0;WeightsStore[3][668]<=0;WeightsStore[3][669]<=0;WeightsStore[3][670]<=0;WeightsStore[3][671]<=0;WeightsStore[3][672]<=0;WeightsStore[3][673]<=0;WeightsStore[3][674]<=0;WeightsStore[3][675]<=0;WeightsStore[3][676]<=0;WeightsStore[3][677]<=0;WeightsStore[3][678]<=0;WeightsStore[3][679]<=0;WeightsStore[3][680]<=0;WeightsStore[3][681]<=0;WeightsStore[3][682]<=0;WeightsStore[3][683]<=0;WeightsStore[3][684]<=0;WeightsStore[3][685]<=0;WeightsStore[3][686]<=0;WeightsStore[3][687]<=0;WeightsStore[3][688]<=0;WeightsStore[3][689]<=0;WeightsStore[3][690]<=0;WeightsStore[3][691]<=0;WeightsStore[3][692]<=0;WeightsStore[3][693]<=0;WeightsStore[3][694]<=0;WeightsStore[3][695]<=0;WeightsStore[3][696]<=0;WeightsStore[3][697]<=0;WeightsStore[3][698]<=0;WeightsStore[3][699]<=0;WeightsStore[3][700]<=0;WeightsStore[3][701]<=0;WeightsStore[3][702]<=0;WeightsStore[3][703]<=0;WeightsStore[3][704]<=0;WeightsStore[3][705]<=0;WeightsStore[3][706]<=0;WeightsStore[3][707]<=0;WeightsStore[3][708]<=0;WeightsStore[3][709]<=0;WeightsStore[3][710]<=0;WeightsStore[3][711]<=0;WeightsStore[3][712]<=0;WeightsStore[3][713]<=0;WeightsStore[3][714]<=0;WeightsStore[3][715]<=0;WeightsStore[3][716]<=0;WeightsStore[3][717]<=0;WeightsStore[3][718]<=0;WeightsStore[3][719]<=0;WeightsStore[3][720]<=0;WeightsStore[3][721]<=0;WeightsStore[3][722]<=0;WeightsStore[3][723]<=0;WeightsStore[3][724]<=0;WeightsStore[3][725]<=0;WeightsStore[3][726]<=0;WeightsStore[3][727]<=0;WeightsStore[3][728]<=0;WeightsStore[3][729]<=0;WeightsStore[3][730]<=0;WeightsStore[3][731]<=0;WeightsStore[3][732]<=0;WeightsStore[3][733]<=0;WeightsStore[3][734]<=0;WeightsStore[3][735]<=0;WeightsStore[3][736]<=0;WeightsStore[3][737]<=0;WeightsStore[3][738]<=0;WeightsStore[3][739]<=0;WeightsStore[3][740]<=0;WeightsStore[3][741]<=0;WeightsStore[3][742]<=0;WeightsStore[3][743]<=0;WeightsStore[3][744]<=0;WeightsStore[3][745]<=0;WeightsStore[3][746]<=0;WeightsStore[3][747]<=0;WeightsStore[3][748]<=0;WeightsStore[3][749]<=0;WeightsStore[3][750]<=0;WeightsStore[3][751]<=0;WeightsStore[3][752]<=0;WeightsStore[3][753]<=0;WeightsStore[3][754]<=0;WeightsStore[3][755]<=0;WeightsStore[3][756]<=0;WeightsStore[3][757]<=0;WeightsStore[3][758]<=0;WeightsStore[3][759]<=0;WeightsStore[3][760]<=0;WeightsStore[3][761]<=0;WeightsStore[3][762]<=0;WeightsStore[3][763]<=0;WeightsStore[3][764]<=0;WeightsStore[3][765]<=0;WeightsStore[3][766]<=0;WeightsStore[3][767]<=0;WeightsStore[3][768]<=0;WeightsStore[3][769]<=0;WeightsStore[3][770]<=0;WeightsStore[3][771]<=0;WeightsStore[3][772]<=0;WeightsStore[3][773]<=0;WeightsStore[3][774]<=0;WeightsStore[3][775]<=0;WeightsStore[3][776]<=0;WeightsStore[3][777]<=0;WeightsStore[3][778]<=0;WeightsStore[3][779]<=0;WeightsStore[3][780]<=0;WeightsStore[3][781]<=0;WeightsStore[3][782]<=0;WeightsStore[3][783]<=0;WeightsStore[3][784]<=0;WeightsStore[4][0]<=0;WeightsStore[4][1]<=0;WeightsStore[4][2]<=0;WeightsStore[4][3]<=0;WeightsStore[4][4]<=0;WeightsStore[4][5]<=0;WeightsStore[4][6]<=0;WeightsStore[4][7]<=0;WeightsStore[4][8]<=0;WeightsStore[4][9]<=0;WeightsStore[4][10]<=0;WeightsStore[4][11]<=0;WeightsStore[4][12]<=0;WeightsStore[4][13]<=0;WeightsStore[4][14]<=0;WeightsStore[4][15]<=0;WeightsStore[4][16]<=0;WeightsStore[4][17]<=0;WeightsStore[4][18]<=0;WeightsStore[4][19]<=0;WeightsStore[4][20]<=0;WeightsStore[4][21]<=0;WeightsStore[4][22]<=0;WeightsStore[4][23]<=0;WeightsStore[4][24]<=0;WeightsStore[4][25]<=0;WeightsStore[4][26]<=0;WeightsStore[4][27]<=0;WeightsStore[4][28]<=0;WeightsStore[4][29]<=0;WeightsStore[4][30]<=0;WeightsStore[4][31]<=0;WeightsStore[4][32]<=0;WeightsStore[4][33]<=0;WeightsStore[4][34]<=0;WeightsStore[4][35]<=0;WeightsStore[4][36]<=0;WeightsStore[4][37]<=0;WeightsStore[4][38]<=0;WeightsStore[4][39]<=0;WeightsStore[4][40]<=0;WeightsStore[4][41]<=0;WeightsStore[4][42]<=0;WeightsStore[4][43]<=0;WeightsStore[4][44]<=0;WeightsStore[4][45]<=0;WeightsStore[4][46]<=0;WeightsStore[4][47]<=0;WeightsStore[4][48]<=0;WeightsStore[4][49]<=0;WeightsStore[4][50]<=0;WeightsStore[4][51]<=0;WeightsStore[4][52]<=0;WeightsStore[4][53]<=0;WeightsStore[4][54]<=0;WeightsStore[4][55]<=0;WeightsStore[4][56]<=0;WeightsStore[4][57]<=0;WeightsStore[4][58]<=0;WeightsStore[4][59]<=0;WeightsStore[4][60]<=0;WeightsStore[4][61]<=0;WeightsStore[4][62]<=0;WeightsStore[4][63]<=0;WeightsStore[4][64]<=0;WeightsStore[4][65]<=0;WeightsStore[4][66]<=0;WeightsStore[4][67]<=0;WeightsStore[4][68]<=0;WeightsStore[4][69]<=0;WeightsStore[4][70]<=0;WeightsStore[4][71]<=0;WeightsStore[4][72]<=0;WeightsStore[4][73]<=0;WeightsStore[4][74]<=0;WeightsStore[4][75]<=0;WeightsStore[4][76]<=0;WeightsStore[4][77]<=0;WeightsStore[4][78]<=0;WeightsStore[4][79]<=0;WeightsStore[4][80]<=0;WeightsStore[4][81]<=0;WeightsStore[4][82]<=0;WeightsStore[4][83]<=0;WeightsStore[4][84]<=0;WeightsStore[4][85]<=0;WeightsStore[4][86]<=0;WeightsStore[4][87]<=0;WeightsStore[4][88]<=0;WeightsStore[4][89]<=0;WeightsStore[4][90]<=0;WeightsStore[4][91]<=0;WeightsStore[4][92]<=0;WeightsStore[4][93]<=0;WeightsStore[4][94]<=0;WeightsStore[4][95]<=0;WeightsStore[4][96]<=0;WeightsStore[4][97]<=0;WeightsStore[4][98]<=0;WeightsStore[4][99]<=0;WeightsStore[4][100]<=0;WeightsStore[4][101]<=0;WeightsStore[4][102]<=0;WeightsStore[4][103]<=0;WeightsStore[4][104]<=0;WeightsStore[4][105]<=0;WeightsStore[4][106]<=0;WeightsStore[4][107]<=0;WeightsStore[4][108]<=0;WeightsStore[4][109]<=0;WeightsStore[4][110]<=0;WeightsStore[4][111]<=0;WeightsStore[4][112]<=0;WeightsStore[4][113]<=0;WeightsStore[4][114]<=0;WeightsStore[4][115]<=0;WeightsStore[4][116]<=0;WeightsStore[4][117]<=0;WeightsStore[4][118]<=0;WeightsStore[4][119]<=0;WeightsStore[4][120]<=0;WeightsStore[4][121]<=0;WeightsStore[4][122]<=0;WeightsStore[4][123]<=0;WeightsStore[4][124]<=0;WeightsStore[4][125]<=0;WeightsStore[4][126]<=0;WeightsStore[4][127]<=0;WeightsStore[4][128]<=0;WeightsStore[4][129]<=0;WeightsStore[4][130]<=0;WeightsStore[4][131]<=0;WeightsStore[4][132]<=0;WeightsStore[4][133]<=0;WeightsStore[4][134]<=0;WeightsStore[4][135]<=0;WeightsStore[4][136]<=0;WeightsStore[4][137]<=0;WeightsStore[4][138]<=0;WeightsStore[4][139]<=0;WeightsStore[4][140]<=0;WeightsStore[4][141]<=0;WeightsStore[4][142]<=0;WeightsStore[4][143]<=0;WeightsStore[4][144]<=0;WeightsStore[4][145]<=0;WeightsStore[4][146]<=0;WeightsStore[4][147]<=0;WeightsStore[4][148]<=0;WeightsStore[4][149]<=0;WeightsStore[4][150]<=0;WeightsStore[4][151]<=0;WeightsStore[4][152]<=0;WeightsStore[4][153]<=0;WeightsStore[4][154]<=0;WeightsStore[4][155]<=0;WeightsStore[4][156]<=0;WeightsStore[4][157]<=0;WeightsStore[4][158]<=0;WeightsStore[4][159]<=0;WeightsStore[4][160]<=0;WeightsStore[4][161]<=0;WeightsStore[4][162]<=0;WeightsStore[4][163]<=0;WeightsStore[4][164]<=0;WeightsStore[4][165]<=0;WeightsStore[4][166]<=0;WeightsStore[4][167]<=0;WeightsStore[4][168]<=0;WeightsStore[4][169]<=0;WeightsStore[4][170]<=0;WeightsStore[4][171]<=0;WeightsStore[4][172]<=0;WeightsStore[4][173]<=0;WeightsStore[4][174]<=0;WeightsStore[4][175]<=0;WeightsStore[4][176]<=0;WeightsStore[4][177]<=0;WeightsStore[4][178]<=0;WeightsStore[4][179]<=0;WeightsStore[4][180]<=0;WeightsStore[4][181]<=0;WeightsStore[4][182]<=0;WeightsStore[4][183]<=0;WeightsStore[4][184]<=0;WeightsStore[4][185]<=0;WeightsStore[4][186]<=0;WeightsStore[4][187]<=0;WeightsStore[4][188]<=0;WeightsStore[4][189]<=0;WeightsStore[4][190]<=0;WeightsStore[4][191]<=0;WeightsStore[4][192]<=0;WeightsStore[4][193]<=0;WeightsStore[4][194]<=0;WeightsStore[4][195]<=0;WeightsStore[4][196]<=0;WeightsStore[4][197]<=0;WeightsStore[4][198]<=0;WeightsStore[4][199]<=0;WeightsStore[4][200]<=0;WeightsStore[4][201]<=0;WeightsStore[4][202]<=0;WeightsStore[4][203]<=0;WeightsStore[4][204]<=0;WeightsStore[4][205]<=0;WeightsStore[4][206]<=0;WeightsStore[4][207]<=0;WeightsStore[4][208]<=0;WeightsStore[4][209]<=0;WeightsStore[4][210]<=0;WeightsStore[4][211]<=0;WeightsStore[4][212]<=0;WeightsStore[4][213]<=0;WeightsStore[4][214]<=0;WeightsStore[4][215]<=0;WeightsStore[4][216]<=0;WeightsStore[4][217]<=0;WeightsStore[4][218]<=0;WeightsStore[4][219]<=0;WeightsStore[4][220]<=0;WeightsStore[4][221]<=0;WeightsStore[4][222]<=0;WeightsStore[4][223]<=0;WeightsStore[4][224]<=0;WeightsStore[4][225]<=0;WeightsStore[4][226]<=0;WeightsStore[4][227]<=0;WeightsStore[4][228]<=0;WeightsStore[4][229]<=0;WeightsStore[4][230]<=0;WeightsStore[4][231]<=0;WeightsStore[4][232]<=0;WeightsStore[4][233]<=0;WeightsStore[4][234]<=0;WeightsStore[4][235]<=0;WeightsStore[4][236]<=0;WeightsStore[4][237]<=0;WeightsStore[4][238]<=0;WeightsStore[4][239]<=0;WeightsStore[4][240]<=0;WeightsStore[4][241]<=0;WeightsStore[4][242]<=0;WeightsStore[4][243]<=0;WeightsStore[4][244]<=0;WeightsStore[4][245]<=0;WeightsStore[4][246]<=0;WeightsStore[4][247]<=0;WeightsStore[4][248]<=0;WeightsStore[4][249]<=0;WeightsStore[4][250]<=0;WeightsStore[4][251]<=0;WeightsStore[4][252]<=0;WeightsStore[4][253]<=0;WeightsStore[4][254]<=0;WeightsStore[4][255]<=0;WeightsStore[4][256]<=0;WeightsStore[4][257]<=0;WeightsStore[4][258]<=0;WeightsStore[4][259]<=0;WeightsStore[4][260]<=0;WeightsStore[4][261]<=0;WeightsStore[4][262]<=0;WeightsStore[4][263]<=0;WeightsStore[4][264]<=0;WeightsStore[4][265]<=0;WeightsStore[4][266]<=0;WeightsStore[4][267]<=0;WeightsStore[4][268]<=0;WeightsStore[4][269]<=0;WeightsStore[4][270]<=0;WeightsStore[4][271]<=0;WeightsStore[4][272]<=0;WeightsStore[4][273]<=0;WeightsStore[4][274]<=0;WeightsStore[4][275]<=0;WeightsStore[4][276]<=0;WeightsStore[4][277]<=0;WeightsStore[4][278]<=0;WeightsStore[4][279]<=0;WeightsStore[4][280]<=0;WeightsStore[4][281]<=0;WeightsStore[4][282]<=0;WeightsStore[4][283]<=0;WeightsStore[4][284]<=0;WeightsStore[4][285]<=0;WeightsStore[4][286]<=0;WeightsStore[4][287]<=0;WeightsStore[4][288]<=0;WeightsStore[4][289]<=0;WeightsStore[4][290]<=0;WeightsStore[4][291]<=0;WeightsStore[4][292]<=0;WeightsStore[4][293]<=0;WeightsStore[4][294]<=0;WeightsStore[4][295]<=0;WeightsStore[4][296]<=0;WeightsStore[4][297]<=0;WeightsStore[4][298]<=0;WeightsStore[4][299]<=0;WeightsStore[4][300]<=0;WeightsStore[4][301]<=0;WeightsStore[4][302]<=0;WeightsStore[4][303]<=0;WeightsStore[4][304]<=0;WeightsStore[4][305]<=0;WeightsStore[4][306]<=0;WeightsStore[4][307]<=0;WeightsStore[4][308]<=0;WeightsStore[4][309]<=0;WeightsStore[4][310]<=0;WeightsStore[4][311]<=0;WeightsStore[4][312]<=0;WeightsStore[4][313]<=0;WeightsStore[4][314]<=0;WeightsStore[4][315]<=0;WeightsStore[4][316]<=0;WeightsStore[4][317]<=0;WeightsStore[4][318]<=0;WeightsStore[4][319]<=0;WeightsStore[4][320]<=0;WeightsStore[4][321]<=0;WeightsStore[4][322]<=0;WeightsStore[4][323]<=0;WeightsStore[4][324]<=0;WeightsStore[4][325]<=0;WeightsStore[4][326]<=0;WeightsStore[4][327]<=0;WeightsStore[4][328]<=0;WeightsStore[4][329]<=0;WeightsStore[4][330]<=0;WeightsStore[4][331]<=0;WeightsStore[4][332]<=0;WeightsStore[4][333]<=0;WeightsStore[4][334]<=0;WeightsStore[4][335]<=0;WeightsStore[4][336]<=0;WeightsStore[4][337]<=0;WeightsStore[4][338]<=0;WeightsStore[4][339]<=0;WeightsStore[4][340]<=0;WeightsStore[4][341]<=0;WeightsStore[4][342]<=0;WeightsStore[4][343]<=0;WeightsStore[4][344]<=0;WeightsStore[4][345]<=0;WeightsStore[4][346]<=0;WeightsStore[4][347]<=0;WeightsStore[4][348]<=0;WeightsStore[4][349]<=0;WeightsStore[4][350]<=0;WeightsStore[4][351]<=0;WeightsStore[4][352]<=0;WeightsStore[4][353]<=0;WeightsStore[4][354]<=0;WeightsStore[4][355]<=0;WeightsStore[4][356]<=0;WeightsStore[4][357]<=0;WeightsStore[4][358]<=0;WeightsStore[4][359]<=0;WeightsStore[4][360]<=0;WeightsStore[4][361]<=0;WeightsStore[4][362]<=0;WeightsStore[4][363]<=0;WeightsStore[4][364]<=0;WeightsStore[4][365]<=0;WeightsStore[4][366]<=0;WeightsStore[4][367]<=0;WeightsStore[4][368]<=0;WeightsStore[4][369]<=0;WeightsStore[4][370]<=0;WeightsStore[4][371]<=0;WeightsStore[4][372]<=0;WeightsStore[4][373]<=0;WeightsStore[4][374]<=0;WeightsStore[4][375]<=0;WeightsStore[4][376]<=0;WeightsStore[4][377]<=0;WeightsStore[4][378]<=0;WeightsStore[4][379]<=0;WeightsStore[4][380]<=0;WeightsStore[4][381]<=0;WeightsStore[4][382]<=0;WeightsStore[4][383]<=0;WeightsStore[4][384]<=0;WeightsStore[4][385]<=0;WeightsStore[4][386]<=0;WeightsStore[4][387]<=0;WeightsStore[4][388]<=0;WeightsStore[4][389]<=0;WeightsStore[4][390]<=0;WeightsStore[4][391]<=0;WeightsStore[4][392]<=0;WeightsStore[4][393]<=0;WeightsStore[4][394]<=0;WeightsStore[4][395]<=0;WeightsStore[4][396]<=0;WeightsStore[4][397]<=0;WeightsStore[4][398]<=0;WeightsStore[4][399]<=0;WeightsStore[4][400]<=0;WeightsStore[4][401]<=0;WeightsStore[4][402]<=0;WeightsStore[4][403]<=0;WeightsStore[4][404]<=0;WeightsStore[4][405]<=0;WeightsStore[4][406]<=0;WeightsStore[4][407]<=0;WeightsStore[4][408]<=0;WeightsStore[4][409]<=0;WeightsStore[4][410]<=0;WeightsStore[4][411]<=0;WeightsStore[4][412]<=0;WeightsStore[4][413]<=0;WeightsStore[4][414]<=0;WeightsStore[4][415]<=0;WeightsStore[4][416]<=0;WeightsStore[4][417]<=0;WeightsStore[4][418]<=0;WeightsStore[4][419]<=0;WeightsStore[4][420]<=0;WeightsStore[4][421]<=0;WeightsStore[4][422]<=0;WeightsStore[4][423]<=0;WeightsStore[4][424]<=0;WeightsStore[4][425]<=0;WeightsStore[4][426]<=0;WeightsStore[4][427]<=0;WeightsStore[4][428]<=0;WeightsStore[4][429]<=0;WeightsStore[4][430]<=0;WeightsStore[4][431]<=0;WeightsStore[4][432]<=0;WeightsStore[4][433]<=0;WeightsStore[4][434]<=0;WeightsStore[4][435]<=0;WeightsStore[4][436]<=0;WeightsStore[4][437]<=0;WeightsStore[4][438]<=0;WeightsStore[4][439]<=0;WeightsStore[4][440]<=0;WeightsStore[4][441]<=0;WeightsStore[4][442]<=0;WeightsStore[4][443]<=0;WeightsStore[4][444]<=0;WeightsStore[4][445]<=0;WeightsStore[4][446]<=0;WeightsStore[4][447]<=0;WeightsStore[4][448]<=0;WeightsStore[4][449]<=0;WeightsStore[4][450]<=0;WeightsStore[4][451]<=0;WeightsStore[4][452]<=0;WeightsStore[4][453]<=0;WeightsStore[4][454]<=0;WeightsStore[4][455]<=0;WeightsStore[4][456]<=0;WeightsStore[4][457]<=0;WeightsStore[4][458]<=0;WeightsStore[4][459]<=0;WeightsStore[4][460]<=0;WeightsStore[4][461]<=0;WeightsStore[4][462]<=0;WeightsStore[4][463]<=0;WeightsStore[4][464]<=0;WeightsStore[4][465]<=0;WeightsStore[4][466]<=0;WeightsStore[4][467]<=0;WeightsStore[4][468]<=0;WeightsStore[4][469]<=0;WeightsStore[4][470]<=0;WeightsStore[4][471]<=0;WeightsStore[4][472]<=0;WeightsStore[4][473]<=0;WeightsStore[4][474]<=0;WeightsStore[4][475]<=0;WeightsStore[4][476]<=0;WeightsStore[4][477]<=0;WeightsStore[4][478]<=0;WeightsStore[4][479]<=0;WeightsStore[4][480]<=0;WeightsStore[4][481]<=0;WeightsStore[4][482]<=0;WeightsStore[4][483]<=0;WeightsStore[4][484]<=0;WeightsStore[4][485]<=0;WeightsStore[4][486]<=0;WeightsStore[4][487]<=0;WeightsStore[4][488]<=0;WeightsStore[4][489]<=0;WeightsStore[4][490]<=0;WeightsStore[4][491]<=0;WeightsStore[4][492]<=0;WeightsStore[4][493]<=0;WeightsStore[4][494]<=0;WeightsStore[4][495]<=0;WeightsStore[4][496]<=0;WeightsStore[4][497]<=0;WeightsStore[4][498]<=0;WeightsStore[4][499]<=0;WeightsStore[4][500]<=0;WeightsStore[4][501]<=0;WeightsStore[4][502]<=0;WeightsStore[4][503]<=0;WeightsStore[4][504]<=0;WeightsStore[4][505]<=0;WeightsStore[4][506]<=0;WeightsStore[4][507]<=0;WeightsStore[4][508]<=0;WeightsStore[4][509]<=0;WeightsStore[4][510]<=0;WeightsStore[4][511]<=0;WeightsStore[4][512]<=0;WeightsStore[4][513]<=0;WeightsStore[4][514]<=0;WeightsStore[4][515]<=0;WeightsStore[4][516]<=0;WeightsStore[4][517]<=0;WeightsStore[4][518]<=0;WeightsStore[4][519]<=0;WeightsStore[4][520]<=0;WeightsStore[4][521]<=0;WeightsStore[4][522]<=0;WeightsStore[4][523]<=0;WeightsStore[4][524]<=0;WeightsStore[4][525]<=0;WeightsStore[4][526]<=0;WeightsStore[4][527]<=0;WeightsStore[4][528]<=0;WeightsStore[4][529]<=0;WeightsStore[4][530]<=0;WeightsStore[4][531]<=0;WeightsStore[4][532]<=0;WeightsStore[4][533]<=0;WeightsStore[4][534]<=0;WeightsStore[4][535]<=0;WeightsStore[4][536]<=0;WeightsStore[4][537]<=0;WeightsStore[4][538]<=0;WeightsStore[4][539]<=0;WeightsStore[4][540]<=0;WeightsStore[4][541]<=0;WeightsStore[4][542]<=0;WeightsStore[4][543]<=0;WeightsStore[4][544]<=0;WeightsStore[4][545]<=0;WeightsStore[4][546]<=0;WeightsStore[4][547]<=0;WeightsStore[4][548]<=0;WeightsStore[4][549]<=0;WeightsStore[4][550]<=0;WeightsStore[4][551]<=0;WeightsStore[4][552]<=0;WeightsStore[4][553]<=0;WeightsStore[4][554]<=0;WeightsStore[4][555]<=0;WeightsStore[4][556]<=0;WeightsStore[4][557]<=0;WeightsStore[4][558]<=0;WeightsStore[4][559]<=0;WeightsStore[4][560]<=0;WeightsStore[4][561]<=0;WeightsStore[4][562]<=0;WeightsStore[4][563]<=0;WeightsStore[4][564]<=0;WeightsStore[4][565]<=0;WeightsStore[4][566]<=0;WeightsStore[4][567]<=0;WeightsStore[4][568]<=0;WeightsStore[4][569]<=0;WeightsStore[4][570]<=0;WeightsStore[4][571]<=0;WeightsStore[4][572]<=0;WeightsStore[4][573]<=0;WeightsStore[4][574]<=0;WeightsStore[4][575]<=0;WeightsStore[4][576]<=0;WeightsStore[4][577]<=0;WeightsStore[4][578]<=0;WeightsStore[4][579]<=0;WeightsStore[4][580]<=0;WeightsStore[4][581]<=0;WeightsStore[4][582]<=0;WeightsStore[4][583]<=0;WeightsStore[4][584]<=0;WeightsStore[4][585]<=0;WeightsStore[4][586]<=0;WeightsStore[4][587]<=0;WeightsStore[4][588]<=0;WeightsStore[4][589]<=0;WeightsStore[4][590]<=0;WeightsStore[4][591]<=0;WeightsStore[4][592]<=0;WeightsStore[4][593]<=0;WeightsStore[4][594]<=0;WeightsStore[4][595]<=0;WeightsStore[4][596]<=0;WeightsStore[4][597]<=0;WeightsStore[4][598]<=0;WeightsStore[4][599]<=0;WeightsStore[4][600]<=0;WeightsStore[4][601]<=0;WeightsStore[4][602]<=0;WeightsStore[4][603]<=0;WeightsStore[4][604]<=0;WeightsStore[4][605]<=0;WeightsStore[4][606]<=0;WeightsStore[4][607]<=0;WeightsStore[4][608]<=0;WeightsStore[4][609]<=0;WeightsStore[4][610]<=0;WeightsStore[4][611]<=0;WeightsStore[4][612]<=0;WeightsStore[4][613]<=0;WeightsStore[4][614]<=0;WeightsStore[4][615]<=0;WeightsStore[4][616]<=0;WeightsStore[4][617]<=0;WeightsStore[4][618]<=0;WeightsStore[4][619]<=0;WeightsStore[4][620]<=0;WeightsStore[4][621]<=0;WeightsStore[4][622]<=0;WeightsStore[4][623]<=0;WeightsStore[4][624]<=0;WeightsStore[4][625]<=0;WeightsStore[4][626]<=0;WeightsStore[4][627]<=0;WeightsStore[4][628]<=0;WeightsStore[4][629]<=0;WeightsStore[4][630]<=0;WeightsStore[4][631]<=0;WeightsStore[4][632]<=0;WeightsStore[4][633]<=0;WeightsStore[4][634]<=0;WeightsStore[4][635]<=0;WeightsStore[4][636]<=0;WeightsStore[4][637]<=0;WeightsStore[4][638]<=0;WeightsStore[4][639]<=0;WeightsStore[4][640]<=0;WeightsStore[4][641]<=0;WeightsStore[4][642]<=0;WeightsStore[4][643]<=0;WeightsStore[4][644]<=0;WeightsStore[4][645]<=0;WeightsStore[4][646]<=0;WeightsStore[4][647]<=0;WeightsStore[4][648]<=0;WeightsStore[4][649]<=0;WeightsStore[4][650]<=0;WeightsStore[4][651]<=0;WeightsStore[4][652]<=0;WeightsStore[4][653]<=0;WeightsStore[4][654]<=0;WeightsStore[4][655]<=0;WeightsStore[4][656]<=0;WeightsStore[4][657]<=0;WeightsStore[4][658]<=0;WeightsStore[4][659]<=0;WeightsStore[4][660]<=0;WeightsStore[4][661]<=0;WeightsStore[4][662]<=0;WeightsStore[4][663]<=0;WeightsStore[4][664]<=0;WeightsStore[4][665]<=0;WeightsStore[4][666]<=0;WeightsStore[4][667]<=0;WeightsStore[4][668]<=0;WeightsStore[4][669]<=0;WeightsStore[4][670]<=0;WeightsStore[4][671]<=0;WeightsStore[4][672]<=0;WeightsStore[4][673]<=0;WeightsStore[4][674]<=0;WeightsStore[4][675]<=0;WeightsStore[4][676]<=0;WeightsStore[4][677]<=0;WeightsStore[4][678]<=0;WeightsStore[4][679]<=0;WeightsStore[4][680]<=0;WeightsStore[4][681]<=0;WeightsStore[4][682]<=0;WeightsStore[4][683]<=0;WeightsStore[4][684]<=0;WeightsStore[4][685]<=0;WeightsStore[4][686]<=0;WeightsStore[4][687]<=0;WeightsStore[4][688]<=0;WeightsStore[4][689]<=0;WeightsStore[4][690]<=0;WeightsStore[4][691]<=0;WeightsStore[4][692]<=0;WeightsStore[4][693]<=0;WeightsStore[4][694]<=0;WeightsStore[4][695]<=0;WeightsStore[4][696]<=0;WeightsStore[4][697]<=0;WeightsStore[4][698]<=0;WeightsStore[4][699]<=0;WeightsStore[4][700]<=0;WeightsStore[4][701]<=0;WeightsStore[4][702]<=0;WeightsStore[4][703]<=0;WeightsStore[4][704]<=0;WeightsStore[4][705]<=0;WeightsStore[4][706]<=0;WeightsStore[4][707]<=0;WeightsStore[4][708]<=0;WeightsStore[4][709]<=0;WeightsStore[4][710]<=0;WeightsStore[4][711]<=0;WeightsStore[4][712]<=0;WeightsStore[4][713]<=0;WeightsStore[4][714]<=0;WeightsStore[4][715]<=0;WeightsStore[4][716]<=0;WeightsStore[4][717]<=0;WeightsStore[4][718]<=0;WeightsStore[4][719]<=0;WeightsStore[4][720]<=0;WeightsStore[4][721]<=0;WeightsStore[4][722]<=0;WeightsStore[4][723]<=0;WeightsStore[4][724]<=0;WeightsStore[4][725]<=0;WeightsStore[4][726]<=0;WeightsStore[4][727]<=0;WeightsStore[4][728]<=0;WeightsStore[4][729]<=0;WeightsStore[4][730]<=0;WeightsStore[4][731]<=0;WeightsStore[4][732]<=0;WeightsStore[4][733]<=0;WeightsStore[4][734]<=0;WeightsStore[4][735]<=0;WeightsStore[4][736]<=0;WeightsStore[4][737]<=0;WeightsStore[4][738]<=0;WeightsStore[4][739]<=0;WeightsStore[4][740]<=0;WeightsStore[4][741]<=0;WeightsStore[4][742]<=0;WeightsStore[4][743]<=0;WeightsStore[4][744]<=0;WeightsStore[4][745]<=0;WeightsStore[4][746]<=0;WeightsStore[4][747]<=0;WeightsStore[4][748]<=0;WeightsStore[4][749]<=0;WeightsStore[4][750]<=0;WeightsStore[4][751]<=0;WeightsStore[4][752]<=0;WeightsStore[4][753]<=0;WeightsStore[4][754]<=0;WeightsStore[4][755]<=0;WeightsStore[4][756]<=0;WeightsStore[4][757]<=0;WeightsStore[4][758]<=0;WeightsStore[4][759]<=0;WeightsStore[4][760]<=0;WeightsStore[4][761]<=0;WeightsStore[4][762]<=0;WeightsStore[4][763]<=0;WeightsStore[4][764]<=0;WeightsStore[4][765]<=0;WeightsStore[4][766]<=0;WeightsStore[4][767]<=0;WeightsStore[4][768]<=0;WeightsStore[4][769]<=0;WeightsStore[4][770]<=0;WeightsStore[4][771]<=0;WeightsStore[4][772]<=0;WeightsStore[4][773]<=0;WeightsStore[4][774]<=0;WeightsStore[4][775]<=0;WeightsStore[4][776]<=0;WeightsStore[4][777]<=0;WeightsStore[4][778]<=0;WeightsStore[4][779]<=0;WeightsStore[4][780]<=0;WeightsStore[4][781]<=0;WeightsStore[4][782]<=0;WeightsStore[4][783]<=0;WeightsStore[4][784]<=0;WeightsStore[5][0]<=0;WeightsStore[5][1]<=0;WeightsStore[5][2]<=0;WeightsStore[5][3]<=0;WeightsStore[5][4]<=0;WeightsStore[5][5]<=0;WeightsStore[5][6]<=0;WeightsStore[5][7]<=0;WeightsStore[5][8]<=0;WeightsStore[5][9]<=0;WeightsStore[5][10]<=0;WeightsStore[5][11]<=0;WeightsStore[5][12]<=0;WeightsStore[5][13]<=0;WeightsStore[5][14]<=0;WeightsStore[5][15]<=0;WeightsStore[5][16]<=0;WeightsStore[5][17]<=0;WeightsStore[5][18]<=0;WeightsStore[5][19]<=0;WeightsStore[5][20]<=0;WeightsStore[5][21]<=0;WeightsStore[5][22]<=0;WeightsStore[5][23]<=0;WeightsStore[5][24]<=0;WeightsStore[5][25]<=0;WeightsStore[5][26]<=0;WeightsStore[5][27]<=0;WeightsStore[5][28]<=0;WeightsStore[5][29]<=0;WeightsStore[5][30]<=0;WeightsStore[5][31]<=0;WeightsStore[5][32]<=0;WeightsStore[5][33]<=0;WeightsStore[5][34]<=0;WeightsStore[5][35]<=0;WeightsStore[5][36]<=0;WeightsStore[5][37]<=0;WeightsStore[5][38]<=0;WeightsStore[5][39]<=0;WeightsStore[5][40]<=0;WeightsStore[5][41]<=0;WeightsStore[5][42]<=0;WeightsStore[5][43]<=0;WeightsStore[5][44]<=0;WeightsStore[5][45]<=0;WeightsStore[5][46]<=0;WeightsStore[5][47]<=0;WeightsStore[5][48]<=0;WeightsStore[5][49]<=0;WeightsStore[5][50]<=0;WeightsStore[5][51]<=0;WeightsStore[5][52]<=0;WeightsStore[5][53]<=0;WeightsStore[5][54]<=0;WeightsStore[5][55]<=0;WeightsStore[5][56]<=0;WeightsStore[5][57]<=0;WeightsStore[5][58]<=0;WeightsStore[5][59]<=0;WeightsStore[5][60]<=0;WeightsStore[5][61]<=0;WeightsStore[5][62]<=0;WeightsStore[5][63]<=0;WeightsStore[5][64]<=0;WeightsStore[5][65]<=0;WeightsStore[5][66]<=0;WeightsStore[5][67]<=0;WeightsStore[5][68]<=0;WeightsStore[5][69]<=0;WeightsStore[5][70]<=0;WeightsStore[5][71]<=0;WeightsStore[5][72]<=0;WeightsStore[5][73]<=0;WeightsStore[5][74]<=0;WeightsStore[5][75]<=0;WeightsStore[5][76]<=0;WeightsStore[5][77]<=0;WeightsStore[5][78]<=0;WeightsStore[5][79]<=0;WeightsStore[5][80]<=0;WeightsStore[5][81]<=0;WeightsStore[5][82]<=0;WeightsStore[5][83]<=0;WeightsStore[5][84]<=0;WeightsStore[5][85]<=0;WeightsStore[5][86]<=0;WeightsStore[5][87]<=0;WeightsStore[5][88]<=0;WeightsStore[5][89]<=0;WeightsStore[5][90]<=0;WeightsStore[5][91]<=0;WeightsStore[5][92]<=0;WeightsStore[5][93]<=0;WeightsStore[5][94]<=0;WeightsStore[5][95]<=0;WeightsStore[5][96]<=0;WeightsStore[5][97]<=0;WeightsStore[5][98]<=0;WeightsStore[5][99]<=0;WeightsStore[5][100]<=0;WeightsStore[5][101]<=0;WeightsStore[5][102]<=0;WeightsStore[5][103]<=0;WeightsStore[5][104]<=0;WeightsStore[5][105]<=0;WeightsStore[5][106]<=0;WeightsStore[5][107]<=0;WeightsStore[5][108]<=0;WeightsStore[5][109]<=0;WeightsStore[5][110]<=0;WeightsStore[5][111]<=0;WeightsStore[5][112]<=0;WeightsStore[5][113]<=0;WeightsStore[5][114]<=0;WeightsStore[5][115]<=0;WeightsStore[5][116]<=0;WeightsStore[5][117]<=0;WeightsStore[5][118]<=0;WeightsStore[5][119]<=0;WeightsStore[5][120]<=0;WeightsStore[5][121]<=0;WeightsStore[5][122]<=0;WeightsStore[5][123]<=0;WeightsStore[5][124]<=0;WeightsStore[5][125]<=0;WeightsStore[5][126]<=0;WeightsStore[5][127]<=0;WeightsStore[5][128]<=0;WeightsStore[5][129]<=0;WeightsStore[5][130]<=0;WeightsStore[5][131]<=0;WeightsStore[5][132]<=0;WeightsStore[5][133]<=0;WeightsStore[5][134]<=0;WeightsStore[5][135]<=0;WeightsStore[5][136]<=0;WeightsStore[5][137]<=0;WeightsStore[5][138]<=0;WeightsStore[5][139]<=0;WeightsStore[5][140]<=0;WeightsStore[5][141]<=0;WeightsStore[5][142]<=0;WeightsStore[5][143]<=0;WeightsStore[5][144]<=0;WeightsStore[5][145]<=0;WeightsStore[5][146]<=0;WeightsStore[5][147]<=0;WeightsStore[5][148]<=0;WeightsStore[5][149]<=0;WeightsStore[5][150]<=0;WeightsStore[5][151]<=0;WeightsStore[5][152]<=0;WeightsStore[5][153]<=0;WeightsStore[5][154]<=0;WeightsStore[5][155]<=0;WeightsStore[5][156]<=0;WeightsStore[5][157]<=0;WeightsStore[5][158]<=0;WeightsStore[5][159]<=0;WeightsStore[5][160]<=0;WeightsStore[5][161]<=0;WeightsStore[5][162]<=0;WeightsStore[5][163]<=0;WeightsStore[5][164]<=0;WeightsStore[5][165]<=0;WeightsStore[5][166]<=0;WeightsStore[5][167]<=0;WeightsStore[5][168]<=0;WeightsStore[5][169]<=0;WeightsStore[5][170]<=0;WeightsStore[5][171]<=0;WeightsStore[5][172]<=0;WeightsStore[5][173]<=0;WeightsStore[5][174]<=0;WeightsStore[5][175]<=0;WeightsStore[5][176]<=0;WeightsStore[5][177]<=0;WeightsStore[5][178]<=0;WeightsStore[5][179]<=0;WeightsStore[5][180]<=0;WeightsStore[5][181]<=0;WeightsStore[5][182]<=0;WeightsStore[5][183]<=0;WeightsStore[5][184]<=0;WeightsStore[5][185]<=0;WeightsStore[5][186]<=0;WeightsStore[5][187]<=0;WeightsStore[5][188]<=0;WeightsStore[5][189]<=0;WeightsStore[5][190]<=0;WeightsStore[5][191]<=0;WeightsStore[5][192]<=0;WeightsStore[5][193]<=0;WeightsStore[5][194]<=0;WeightsStore[5][195]<=0;WeightsStore[5][196]<=0;WeightsStore[5][197]<=0;WeightsStore[5][198]<=0;WeightsStore[5][199]<=0;WeightsStore[5][200]<=0;WeightsStore[5][201]<=0;WeightsStore[5][202]<=0;WeightsStore[5][203]<=0;WeightsStore[5][204]<=0;WeightsStore[5][205]<=0;WeightsStore[5][206]<=0;WeightsStore[5][207]<=0;WeightsStore[5][208]<=0;WeightsStore[5][209]<=0;WeightsStore[5][210]<=0;WeightsStore[5][211]<=0;WeightsStore[5][212]<=0;WeightsStore[5][213]<=0;WeightsStore[5][214]<=0;WeightsStore[5][215]<=0;WeightsStore[5][216]<=0;WeightsStore[5][217]<=0;WeightsStore[5][218]<=0;WeightsStore[5][219]<=0;WeightsStore[5][220]<=0;WeightsStore[5][221]<=0;WeightsStore[5][222]<=0;WeightsStore[5][223]<=0;WeightsStore[5][224]<=0;WeightsStore[5][225]<=0;WeightsStore[5][226]<=0;WeightsStore[5][227]<=0;WeightsStore[5][228]<=0;WeightsStore[5][229]<=0;WeightsStore[5][230]<=0;WeightsStore[5][231]<=0;WeightsStore[5][232]<=0;WeightsStore[5][233]<=0;WeightsStore[5][234]<=0;WeightsStore[5][235]<=0;WeightsStore[5][236]<=0;WeightsStore[5][237]<=0;WeightsStore[5][238]<=0;WeightsStore[5][239]<=0;WeightsStore[5][240]<=0;WeightsStore[5][241]<=0;WeightsStore[5][242]<=0;WeightsStore[5][243]<=0;WeightsStore[5][244]<=0;WeightsStore[5][245]<=0;WeightsStore[5][246]<=0;WeightsStore[5][247]<=0;WeightsStore[5][248]<=0;WeightsStore[5][249]<=0;WeightsStore[5][250]<=0;WeightsStore[5][251]<=0;WeightsStore[5][252]<=0;WeightsStore[5][253]<=0;WeightsStore[5][254]<=0;WeightsStore[5][255]<=0;WeightsStore[5][256]<=0;WeightsStore[5][257]<=0;WeightsStore[5][258]<=0;WeightsStore[5][259]<=0;WeightsStore[5][260]<=0;WeightsStore[5][261]<=0;WeightsStore[5][262]<=0;WeightsStore[5][263]<=0;WeightsStore[5][264]<=0;WeightsStore[5][265]<=0;WeightsStore[5][266]<=0;WeightsStore[5][267]<=0;WeightsStore[5][268]<=0;WeightsStore[5][269]<=0;WeightsStore[5][270]<=0;WeightsStore[5][271]<=0;WeightsStore[5][272]<=0;WeightsStore[5][273]<=0;WeightsStore[5][274]<=0;WeightsStore[5][275]<=0;WeightsStore[5][276]<=0;WeightsStore[5][277]<=0;WeightsStore[5][278]<=0;WeightsStore[5][279]<=0;WeightsStore[5][280]<=0;WeightsStore[5][281]<=0;WeightsStore[5][282]<=0;WeightsStore[5][283]<=0;WeightsStore[5][284]<=0;WeightsStore[5][285]<=0;WeightsStore[5][286]<=0;WeightsStore[5][287]<=0;WeightsStore[5][288]<=0;WeightsStore[5][289]<=0;WeightsStore[5][290]<=0;WeightsStore[5][291]<=0;WeightsStore[5][292]<=0;WeightsStore[5][293]<=0;WeightsStore[5][294]<=0;WeightsStore[5][295]<=0;WeightsStore[5][296]<=0;WeightsStore[5][297]<=0;WeightsStore[5][298]<=0;WeightsStore[5][299]<=0;WeightsStore[5][300]<=0;WeightsStore[5][301]<=0;WeightsStore[5][302]<=0;WeightsStore[5][303]<=0;WeightsStore[5][304]<=0;WeightsStore[5][305]<=0;WeightsStore[5][306]<=0;WeightsStore[5][307]<=0;WeightsStore[5][308]<=0;WeightsStore[5][309]<=0;WeightsStore[5][310]<=0;WeightsStore[5][311]<=0;WeightsStore[5][312]<=0;WeightsStore[5][313]<=0;WeightsStore[5][314]<=0;WeightsStore[5][315]<=0;WeightsStore[5][316]<=0;WeightsStore[5][317]<=0;WeightsStore[5][318]<=0;WeightsStore[5][319]<=0;WeightsStore[5][320]<=0;WeightsStore[5][321]<=0;WeightsStore[5][322]<=0;WeightsStore[5][323]<=0;WeightsStore[5][324]<=0;WeightsStore[5][325]<=0;WeightsStore[5][326]<=0;WeightsStore[5][327]<=0;WeightsStore[5][328]<=0;WeightsStore[5][329]<=0;WeightsStore[5][330]<=0;WeightsStore[5][331]<=0;WeightsStore[5][332]<=0;WeightsStore[5][333]<=0;WeightsStore[5][334]<=0;WeightsStore[5][335]<=0;WeightsStore[5][336]<=0;WeightsStore[5][337]<=0;WeightsStore[5][338]<=0;WeightsStore[5][339]<=0;WeightsStore[5][340]<=0;WeightsStore[5][341]<=0;WeightsStore[5][342]<=0;WeightsStore[5][343]<=0;WeightsStore[5][344]<=0;WeightsStore[5][345]<=0;WeightsStore[5][346]<=0;WeightsStore[5][347]<=0;WeightsStore[5][348]<=0;WeightsStore[5][349]<=0;WeightsStore[5][350]<=0;WeightsStore[5][351]<=0;WeightsStore[5][352]<=0;WeightsStore[5][353]<=0;WeightsStore[5][354]<=0;WeightsStore[5][355]<=0;WeightsStore[5][356]<=0;WeightsStore[5][357]<=0;WeightsStore[5][358]<=0;WeightsStore[5][359]<=0;WeightsStore[5][360]<=0;WeightsStore[5][361]<=0;WeightsStore[5][362]<=0;WeightsStore[5][363]<=0;WeightsStore[5][364]<=0;WeightsStore[5][365]<=0;WeightsStore[5][366]<=0;WeightsStore[5][367]<=0;WeightsStore[5][368]<=0;WeightsStore[5][369]<=0;WeightsStore[5][370]<=0;WeightsStore[5][371]<=0;WeightsStore[5][372]<=0;WeightsStore[5][373]<=0;WeightsStore[5][374]<=0;WeightsStore[5][375]<=0;WeightsStore[5][376]<=0;WeightsStore[5][377]<=0;WeightsStore[5][378]<=0;WeightsStore[5][379]<=0;WeightsStore[5][380]<=0;WeightsStore[5][381]<=0;WeightsStore[5][382]<=0;WeightsStore[5][383]<=0;WeightsStore[5][384]<=0;WeightsStore[5][385]<=0;WeightsStore[5][386]<=0;WeightsStore[5][387]<=0;WeightsStore[5][388]<=0;WeightsStore[5][389]<=0;WeightsStore[5][390]<=0;WeightsStore[5][391]<=0;WeightsStore[5][392]<=0;WeightsStore[5][393]<=0;WeightsStore[5][394]<=0;WeightsStore[5][395]<=0;WeightsStore[5][396]<=0;WeightsStore[5][397]<=0;WeightsStore[5][398]<=0;WeightsStore[5][399]<=0;WeightsStore[5][400]<=0;WeightsStore[5][401]<=0;WeightsStore[5][402]<=0;WeightsStore[5][403]<=0;WeightsStore[5][404]<=0;WeightsStore[5][405]<=0;WeightsStore[5][406]<=0;WeightsStore[5][407]<=0;WeightsStore[5][408]<=0;WeightsStore[5][409]<=0;WeightsStore[5][410]<=0;WeightsStore[5][411]<=0;WeightsStore[5][412]<=0;WeightsStore[5][413]<=0;WeightsStore[5][414]<=0;WeightsStore[5][415]<=0;WeightsStore[5][416]<=0;WeightsStore[5][417]<=0;WeightsStore[5][418]<=0;WeightsStore[5][419]<=0;WeightsStore[5][420]<=0;WeightsStore[5][421]<=0;WeightsStore[5][422]<=0;WeightsStore[5][423]<=0;WeightsStore[5][424]<=0;WeightsStore[5][425]<=0;WeightsStore[5][426]<=0;WeightsStore[5][427]<=0;WeightsStore[5][428]<=0;WeightsStore[5][429]<=0;WeightsStore[5][430]<=0;WeightsStore[5][431]<=0;WeightsStore[5][432]<=0;WeightsStore[5][433]<=0;WeightsStore[5][434]<=0;WeightsStore[5][435]<=0;WeightsStore[5][436]<=0;WeightsStore[5][437]<=0;WeightsStore[5][438]<=0;WeightsStore[5][439]<=0;WeightsStore[5][440]<=0;WeightsStore[5][441]<=0;WeightsStore[5][442]<=0;WeightsStore[5][443]<=0;WeightsStore[5][444]<=0;WeightsStore[5][445]<=0;WeightsStore[5][446]<=0;WeightsStore[5][447]<=0;WeightsStore[5][448]<=0;WeightsStore[5][449]<=0;WeightsStore[5][450]<=0;WeightsStore[5][451]<=0;WeightsStore[5][452]<=0;WeightsStore[5][453]<=0;WeightsStore[5][454]<=0;WeightsStore[5][455]<=0;WeightsStore[5][456]<=0;WeightsStore[5][457]<=0;WeightsStore[5][458]<=0;WeightsStore[5][459]<=0;WeightsStore[5][460]<=0;WeightsStore[5][461]<=0;WeightsStore[5][462]<=0;WeightsStore[5][463]<=0;WeightsStore[5][464]<=0;WeightsStore[5][465]<=0;WeightsStore[5][466]<=0;WeightsStore[5][467]<=0;WeightsStore[5][468]<=0;WeightsStore[5][469]<=0;WeightsStore[5][470]<=0;WeightsStore[5][471]<=0;WeightsStore[5][472]<=0;WeightsStore[5][473]<=0;WeightsStore[5][474]<=0;WeightsStore[5][475]<=0;WeightsStore[5][476]<=0;WeightsStore[5][477]<=0;WeightsStore[5][478]<=0;WeightsStore[5][479]<=0;WeightsStore[5][480]<=0;WeightsStore[5][481]<=0;WeightsStore[5][482]<=0;WeightsStore[5][483]<=0;WeightsStore[5][484]<=0;WeightsStore[5][485]<=0;WeightsStore[5][486]<=0;WeightsStore[5][487]<=0;WeightsStore[5][488]<=0;WeightsStore[5][489]<=0;WeightsStore[5][490]<=0;WeightsStore[5][491]<=0;WeightsStore[5][492]<=0;WeightsStore[5][493]<=0;WeightsStore[5][494]<=0;WeightsStore[5][495]<=0;WeightsStore[5][496]<=0;WeightsStore[5][497]<=0;WeightsStore[5][498]<=0;WeightsStore[5][499]<=0;WeightsStore[5][500]<=0;WeightsStore[5][501]<=0;WeightsStore[5][502]<=0;WeightsStore[5][503]<=0;WeightsStore[5][504]<=0;WeightsStore[5][505]<=0;WeightsStore[5][506]<=0;WeightsStore[5][507]<=0;WeightsStore[5][508]<=0;WeightsStore[5][509]<=0;WeightsStore[5][510]<=0;WeightsStore[5][511]<=0;WeightsStore[5][512]<=0;WeightsStore[5][513]<=0;WeightsStore[5][514]<=0;WeightsStore[5][515]<=0;WeightsStore[5][516]<=0;WeightsStore[5][517]<=0;WeightsStore[5][518]<=0;WeightsStore[5][519]<=0;WeightsStore[5][520]<=0;WeightsStore[5][521]<=0;WeightsStore[5][522]<=0;WeightsStore[5][523]<=0;WeightsStore[5][524]<=0;WeightsStore[5][525]<=0;WeightsStore[5][526]<=0;WeightsStore[5][527]<=0;WeightsStore[5][528]<=0;WeightsStore[5][529]<=0;WeightsStore[5][530]<=0;WeightsStore[5][531]<=0;WeightsStore[5][532]<=0;WeightsStore[5][533]<=0;WeightsStore[5][534]<=0;WeightsStore[5][535]<=0;WeightsStore[5][536]<=0;WeightsStore[5][537]<=0;WeightsStore[5][538]<=0;WeightsStore[5][539]<=0;WeightsStore[5][540]<=0;WeightsStore[5][541]<=0;WeightsStore[5][542]<=0;WeightsStore[5][543]<=0;WeightsStore[5][544]<=0;WeightsStore[5][545]<=0;WeightsStore[5][546]<=0;WeightsStore[5][547]<=0;WeightsStore[5][548]<=0;WeightsStore[5][549]<=0;WeightsStore[5][550]<=0;WeightsStore[5][551]<=0;WeightsStore[5][552]<=0;WeightsStore[5][553]<=0;WeightsStore[5][554]<=0;WeightsStore[5][555]<=0;WeightsStore[5][556]<=0;WeightsStore[5][557]<=0;WeightsStore[5][558]<=0;WeightsStore[5][559]<=0;WeightsStore[5][560]<=0;WeightsStore[5][561]<=0;WeightsStore[5][562]<=0;WeightsStore[5][563]<=0;WeightsStore[5][564]<=0;WeightsStore[5][565]<=0;WeightsStore[5][566]<=0;WeightsStore[5][567]<=0;WeightsStore[5][568]<=0;WeightsStore[5][569]<=0;WeightsStore[5][570]<=0;WeightsStore[5][571]<=0;WeightsStore[5][572]<=0;WeightsStore[5][573]<=0;WeightsStore[5][574]<=0;WeightsStore[5][575]<=0;WeightsStore[5][576]<=0;WeightsStore[5][577]<=0;WeightsStore[5][578]<=0;WeightsStore[5][579]<=0;WeightsStore[5][580]<=0;WeightsStore[5][581]<=0;WeightsStore[5][582]<=0;WeightsStore[5][583]<=0;WeightsStore[5][584]<=0;WeightsStore[5][585]<=0;WeightsStore[5][586]<=0;WeightsStore[5][587]<=0;WeightsStore[5][588]<=0;WeightsStore[5][589]<=0;WeightsStore[5][590]<=0;WeightsStore[5][591]<=0;WeightsStore[5][592]<=0;WeightsStore[5][593]<=0;WeightsStore[5][594]<=0;WeightsStore[5][595]<=0;WeightsStore[5][596]<=0;WeightsStore[5][597]<=0;WeightsStore[5][598]<=0;WeightsStore[5][599]<=0;WeightsStore[5][600]<=0;WeightsStore[5][601]<=0;WeightsStore[5][602]<=0;WeightsStore[5][603]<=0;WeightsStore[5][604]<=0;WeightsStore[5][605]<=0;WeightsStore[5][606]<=0;WeightsStore[5][607]<=0;WeightsStore[5][608]<=0;WeightsStore[5][609]<=0;WeightsStore[5][610]<=0;WeightsStore[5][611]<=0;WeightsStore[5][612]<=0;WeightsStore[5][613]<=0;WeightsStore[5][614]<=0;WeightsStore[5][615]<=0;WeightsStore[5][616]<=0;WeightsStore[5][617]<=0;WeightsStore[5][618]<=0;WeightsStore[5][619]<=0;WeightsStore[5][620]<=0;WeightsStore[5][621]<=0;WeightsStore[5][622]<=0;WeightsStore[5][623]<=0;WeightsStore[5][624]<=0;WeightsStore[5][625]<=0;WeightsStore[5][626]<=0;WeightsStore[5][627]<=0;WeightsStore[5][628]<=0;WeightsStore[5][629]<=0;WeightsStore[5][630]<=0;WeightsStore[5][631]<=0;WeightsStore[5][632]<=0;WeightsStore[5][633]<=0;WeightsStore[5][634]<=0;WeightsStore[5][635]<=0;WeightsStore[5][636]<=0;WeightsStore[5][637]<=0;WeightsStore[5][638]<=0;WeightsStore[5][639]<=0;WeightsStore[5][640]<=0;WeightsStore[5][641]<=0;WeightsStore[5][642]<=0;WeightsStore[5][643]<=0;WeightsStore[5][644]<=0;WeightsStore[5][645]<=0;WeightsStore[5][646]<=0;WeightsStore[5][647]<=0;WeightsStore[5][648]<=0;WeightsStore[5][649]<=0;WeightsStore[5][650]<=0;WeightsStore[5][651]<=0;WeightsStore[5][652]<=0;WeightsStore[5][653]<=0;WeightsStore[5][654]<=0;WeightsStore[5][655]<=0;WeightsStore[5][656]<=0;WeightsStore[5][657]<=0;WeightsStore[5][658]<=0;WeightsStore[5][659]<=0;WeightsStore[5][660]<=0;WeightsStore[5][661]<=0;WeightsStore[5][662]<=0;WeightsStore[5][663]<=0;WeightsStore[5][664]<=0;WeightsStore[5][665]<=0;WeightsStore[5][666]<=0;WeightsStore[5][667]<=0;WeightsStore[5][668]<=0;WeightsStore[5][669]<=0;WeightsStore[5][670]<=0;WeightsStore[5][671]<=0;WeightsStore[5][672]<=0;WeightsStore[5][673]<=0;WeightsStore[5][674]<=0;WeightsStore[5][675]<=0;WeightsStore[5][676]<=0;WeightsStore[5][677]<=0;WeightsStore[5][678]<=0;WeightsStore[5][679]<=0;WeightsStore[5][680]<=0;WeightsStore[5][681]<=0;WeightsStore[5][682]<=0;WeightsStore[5][683]<=0;WeightsStore[5][684]<=0;WeightsStore[5][685]<=0;WeightsStore[5][686]<=0;WeightsStore[5][687]<=0;WeightsStore[5][688]<=0;WeightsStore[5][689]<=0;WeightsStore[5][690]<=0;WeightsStore[5][691]<=0;WeightsStore[5][692]<=0;WeightsStore[5][693]<=0;WeightsStore[5][694]<=0;WeightsStore[5][695]<=0;WeightsStore[5][696]<=0;WeightsStore[5][697]<=0;WeightsStore[5][698]<=0;WeightsStore[5][699]<=0;WeightsStore[5][700]<=0;WeightsStore[5][701]<=0;WeightsStore[5][702]<=0;WeightsStore[5][703]<=0;WeightsStore[5][704]<=0;WeightsStore[5][705]<=0;WeightsStore[5][706]<=0;WeightsStore[5][707]<=0;WeightsStore[5][708]<=0;WeightsStore[5][709]<=0;WeightsStore[5][710]<=0;WeightsStore[5][711]<=0;WeightsStore[5][712]<=0;WeightsStore[5][713]<=0;WeightsStore[5][714]<=0;WeightsStore[5][715]<=0;WeightsStore[5][716]<=0;WeightsStore[5][717]<=0;WeightsStore[5][718]<=0;WeightsStore[5][719]<=0;WeightsStore[5][720]<=0;WeightsStore[5][721]<=0;WeightsStore[5][722]<=0;WeightsStore[5][723]<=0;WeightsStore[5][724]<=0;WeightsStore[5][725]<=0;WeightsStore[5][726]<=0;WeightsStore[5][727]<=0;WeightsStore[5][728]<=0;WeightsStore[5][729]<=0;WeightsStore[5][730]<=0;WeightsStore[5][731]<=0;WeightsStore[5][732]<=0;WeightsStore[5][733]<=0;WeightsStore[5][734]<=0;WeightsStore[5][735]<=0;WeightsStore[5][736]<=0;WeightsStore[5][737]<=0;WeightsStore[5][738]<=0;WeightsStore[5][739]<=0;WeightsStore[5][740]<=0;WeightsStore[5][741]<=0;WeightsStore[5][742]<=0;WeightsStore[5][743]<=0;WeightsStore[5][744]<=0;WeightsStore[5][745]<=0;WeightsStore[5][746]<=0;WeightsStore[5][747]<=0;WeightsStore[5][748]<=0;WeightsStore[5][749]<=0;WeightsStore[5][750]<=0;WeightsStore[5][751]<=0;WeightsStore[5][752]<=0;WeightsStore[5][753]<=0;WeightsStore[5][754]<=0;WeightsStore[5][755]<=0;WeightsStore[5][756]<=0;WeightsStore[5][757]<=0;WeightsStore[5][758]<=0;WeightsStore[5][759]<=0;WeightsStore[5][760]<=0;WeightsStore[5][761]<=0;WeightsStore[5][762]<=0;WeightsStore[5][763]<=0;WeightsStore[5][764]<=0;WeightsStore[5][765]<=0;WeightsStore[5][766]<=0;WeightsStore[5][767]<=0;WeightsStore[5][768]<=0;WeightsStore[5][769]<=0;WeightsStore[5][770]<=0;WeightsStore[5][771]<=0;WeightsStore[5][772]<=0;WeightsStore[5][773]<=0;WeightsStore[5][774]<=0;WeightsStore[5][775]<=0;WeightsStore[5][776]<=0;WeightsStore[5][777]<=0;WeightsStore[5][778]<=0;WeightsStore[5][779]<=0;WeightsStore[5][780]<=0;WeightsStore[5][781]<=0;WeightsStore[5][782]<=0;WeightsStore[5][783]<=0;WeightsStore[5][784]<=0;WeightsStore[6][0]<=0;WeightsStore[6][1]<=0;WeightsStore[6][2]<=0;WeightsStore[6][3]<=0;WeightsStore[6][4]<=0;WeightsStore[6][5]<=0;WeightsStore[6][6]<=0;WeightsStore[6][7]<=0;WeightsStore[6][8]<=0;WeightsStore[6][9]<=0;WeightsStore[6][10]<=0;WeightsStore[6][11]<=0;WeightsStore[6][12]<=0;WeightsStore[6][13]<=0;WeightsStore[6][14]<=0;WeightsStore[6][15]<=0;WeightsStore[6][16]<=0;WeightsStore[6][17]<=0;WeightsStore[6][18]<=0;WeightsStore[6][19]<=0;WeightsStore[6][20]<=0;WeightsStore[6][21]<=0;WeightsStore[6][22]<=0;WeightsStore[6][23]<=0;WeightsStore[6][24]<=0;WeightsStore[6][25]<=0;WeightsStore[6][26]<=0;WeightsStore[6][27]<=0;WeightsStore[6][28]<=0;WeightsStore[6][29]<=0;WeightsStore[6][30]<=0;WeightsStore[6][31]<=0;WeightsStore[6][32]<=0;WeightsStore[6][33]<=0;WeightsStore[6][34]<=0;WeightsStore[6][35]<=0;WeightsStore[6][36]<=0;WeightsStore[6][37]<=0;WeightsStore[6][38]<=0;WeightsStore[6][39]<=0;WeightsStore[6][40]<=0;WeightsStore[6][41]<=0;WeightsStore[6][42]<=0;WeightsStore[6][43]<=0;WeightsStore[6][44]<=0;WeightsStore[6][45]<=0;WeightsStore[6][46]<=0;WeightsStore[6][47]<=0;WeightsStore[6][48]<=0;WeightsStore[6][49]<=0;WeightsStore[6][50]<=0;WeightsStore[6][51]<=0;WeightsStore[6][52]<=0;WeightsStore[6][53]<=0;WeightsStore[6][54]<=0;WeightsStore[6][55]<=0;WeightsStore[6][56]<=0;WeightsStore[6][57]<=0;WeightsStore[6][58]<=0;WeightsStore[6][59]<=0;WeightsStore[6][60]<=0;WeightsStore[6][61]<=0;WeightsStore[6][62]<=0;WeightsStore[6][63]<=0;WeightsStore[6][64]<=0;WeightsStore[6][65]<=0;WeightsStore[6][66]<=0;WeightsStore[6][67]<=0;WeightsStore[6][68]<=0;WeightsStore[6][69]<=0;WeightsStore[6][70]<=0;WeightsStore[6][71]<=0;WeightsStore[6][72]<=0;WeightsStore[6][73]<=0;WeightsStore[6][74]<=0;WeightsStore[6][75]<=0;WeightsStore[6][76]<=0;WeightsStore[6][77]<=0;WeightsStore[6][78]<=0;WeightsStore[6][79]<=0;WeightsStore[6][80]<=0;WeightsStore[6][81]<=0;WeightsStore[6][82]<=0;WeightsStore[6][83]<=0;WeightsStore[6][84]<=0;WeightsStore[6][85]<=0;WeightsStore[6][86]<=0;WeightsStore[6][87]<=0;WeightsStore[6][88]<=0;WeightsStore[6][89]<=0;WeightsStore[6][90]<=0;WeightsStore[6][91]<=0;WeightsStore[6][92]<=0;WeightsStore[6][93]<=0;WeightsStore[6][94]<=0;WeightsStore[6][95]<=0;WeightsStore[6][96]<=0;WeightsStore[6][97]<=0;WeightsStore[6][98]<=0;WeightsStore[6][99]<=0;WeightsStore[6][100]<=0;WeightsStore[6][101]<=0;WeightsStore[6][102]<=0;WeightsStore[6][103]<=0;WeightsStore[6][104]<=0;WeightsStore[6][105]<=0;WeightsStore[6][106]<=0;WeightsStore[6][107]<=0;WeightsStore[6][108]<=0;WeightsStore[6][109]<=0;WeightsStore[6][110]<=0;WeightsStore[6][111]<=0;WeightsStore[6][112]<=0;WeightsStore[6][113]<=0;WeightsStore[6][114]<=0;WeightsStore[6][115]<=0;WeightsStore[6][116]<=0;WeightsStore[6][117]<=0;WeightsStore[6][118]<=0;WeightsStore[6][119]<=0;WeightsStore[6][120]<=0;WeightsStore[6][121]<=0;WeightsStore[6][122]<=0;WeightsStore[6][123]<=0;WeightsStore[6][124]<=0;WeightsStore[6][125]<=0;WeightsStore[6][126]<=0;WeightsStore[6][127]<=0;WeightsStore[6][128]<=0;WeightsStore[6][129]<=0;WeightsStore[6][130]<=0;WeightsStore[6][131]<=0;WeightsStore[6][132]<=0;WeightsStore[6][133]<=0;WeightsStore[6][134]<=0;WeightsStore[6][135]<=0;WeightsStore[6][136]<=0;WeightsStore[6][137]<=0;WeightsStore[6][138]<=0;WeightsStore[6][139]<=0;WeightsStore[6][140]<=0;WeightsStore[6][141]<=0;WeightsStore[6][142]<=0;WeightsStore[6][143]<=0;WeightsStore[6][144]<=0;WeightsStore[6][145]<=0;WeightsStore[6][146]<=0;WeightsStore[6][147]<=0;WeightsStore[6][148]<=0;WeightsStore[6][149]<=0;WeightsStore[6][150]<=0;WeightsStore[6][151]<=0;WeightsStore[6][152]<=0;WeightsStore[6][153]<=0;WeightsStore[6][154]<=0;WeightsStore[6][155]<=0;WeightsStore[6][156]<=0;WeightsStore[6][157]<=0;WeightsStore[6][158]<=0;WeightsStore[6][159]<=0;WeightsStore[6][160]<=0;WeightsStore[6][161]<=0;WeightsStore[6][162]<=0;WeightsStore[6][163]<=0;WeightsStore[6][164]<=0;WeightsStore[6][165]<=0;WeightsStore[6][166]<=0;WeightsStore[6][167]<=0;WeightsStore[6][168]<=0;WeightsStore[6][169]<=0;WeightsStore[6][170]<=0;WeightsStore[6][171]<=0;WeightsStore[6][172]<=0;WeightsStore[6][173]<=0;WeightsStore[6][174]<=0;WeightsStore[6][175]<=0;WeightsStore[6][176]<=0;WeightsStore[6][177]<=0;WeightsStore[6][178]<=0;WeightsStore[6][179]<=0;WeightsStore[6][180]<=0;WeightsStore[6][181]<=0;WeightsStore[6][182]<=0;WeightsStore[6][183]<=0;WeightsStore[6][184]<=0;WeightsStore[6][185]<=0;WeightsStore[6][186]<=0;WeightsStore[6][187]<=0;WeightsStore[6][188]<=0;WeightsStore[6][189]<=0;WeightsStore[6][190]<=0;WeightsStore[6][191]<=0;WeightsStore[6][192]<=0;WeightsStore[6][193]<=0;WeightsStore[6][194]<=0;WeightsStore[6][195]<=0;WeightsStore[6][196]<=0;WeightsStore[6][197]<=0;WeightsStore[6][198]<=0;WeightsStore[6][199]<=0;WeightsStore[6][200]<=0;WeightsStore[6][201]<=0;WeightsStore[6][202]<=0;WeightsStore[6][203]<=0;WeightsStore[6][204]<=0;WeightsStore[6][205]<=0;WeightsStore[6][206]<=0;WeightsStore[6][207]<=0;WeightsStore[6][208]<=0;WeightsStore[6][209]<=0;WeightsStore[6][210]<=0;WeightsStore[6][211]<=0;WeightsStore[6][212]<=0;WeightsStore[6][213]<=0;WeightsStore[6][214]<=0;WeightsStore[6][215]<=0;WeightsStore[6][216]<=0;WeightsStore[6][217]<=0;WeightsStore[6][218]<=0;WeightsStore[6][219]<=0;WeightsStore[6][220]<=0;WeightsStore[6][221]<=0;WeightsStore[6][222]<=0;WeightsStore[6][223]<=0;WeightsStore[6][224]<=0;WeightsStore[6][225]<=0;WeightsStore[6][226]<=0;WeightsStore[6][227]<=0;WeightsStore[6][228]<=0;WeightsStore[6][229]<=0;WeightsStore[6][230]<=0;WeightsStore[6][231]<=0;WeightsStore[6][232]<=0;WeightsStore[6][233]<=0;WeightsStore[6][234]<=0;WeightsStore[6][235]<=0;WeightsStore[6][236]<=0;WeightsStore[6][237]<=0;WeightsStore[6][238]<=0;WeightsStore[6][239]<=0;WeightsStore[6][240]<=0;WeightsStore[6][241]<=0;WeightsStore[6][242]<=0;WeightsStore[6][243]<=0;WeightsStore[6][244]<=0;WeightsStore[6][245]<=0;WeightsStore[6][246]<=0;WeightsStore[6][247]<=0;WeightsStore[6][248]<=0;WeightsStore[6][249]<=0;WeightsStore[6][250]<=0;WeightsStore[6][251]<=0;WeightsStore[6][252]<=0;WeightsStore[6][253]<=0;WeightsStore[6][254]<=0;WeightsStore[6][255]<=0;WeightsStore[6][256]<=0;WeightsStore[6][257]<=0;WeightsStore[6][258]<=0;WeightsStore[6][259]<=0;WeightsStore[6][260]<=0;WeightsStore[6][261]<=0;WeightsStore[6][262]<=0;WeightsStore[6][263]<=0;WeightsStore[6][264]<=0;WeightsStore[6][265]<=0;WeightsStore[6][266]<=0;WeightsStore[6][267]<=0;WeightsStore[6][268]<=0;WeightsStore[6][269]<=0;WeightsStore[6][270]<=0;WeightsStore[6][271]<=0;WeightsStore[6][272]<=0;WeightsStore[6][273]<=0;WeightsStore[6][274]<=0;WeightsStore[6][275]<=0;WeightsStore[6][276]<=0;WeightsStore[6][277]<=0;WeightsStore[6][278]<=0;WeightsStore[6][279]<=0;WeightsStore[6][280]<=0;WeightsStore[6][281]<=0;WeightsStore[6][282]<=0;WeightsStore[6][283]<=0;WeightsStore[6][284]<=0;WeightsStore[6][285]<=0;WeightsStore[6][286]<=0;WeightsStore[6][287]<=0;WeightsStore[6][288]<=0;WeightsStore[6][289]<=0;WeightsStore[6][290]<=0;WeightsStore[6][291]<=0;WeightsStore[6][292]<=0;WeightsStore[6][293]<=0;WeightsStore[6][294]<=0;WeightsStore[6][295]<=0;WeightsStore[6][296]<=0;WeightsStore[6][297]<=0;WeightsStore[6][298]<=0;WeightsStore[6][299]<=0;WeightsStore[6][300]<=0;WeightsStore[6][301]<=0;WeightsStore[6][302]<=0;WeightsStore[6][303]<=0;WeightsStore[6][304]<=0;WeightsStore[6][305]<=0;WeightsStore[6][306]<=0;WeightsStore[6][307]<=0;WeightsStore[6][308]<=0;WeightsStore[6][309]<=0;WeightsStore[6][310]<=0;WeightsStore[6][311]<=0;WeightsStore[6][312]<=0;WeightsStore[6][313]<=0;WeightsStore[6][314]<=0;WeightsStore[6][315]<=0;WeightsStore[6][316]<=0;WeightsStore[6][317]<=0;WeightsStore[6][318]<=0;WeightsStore[6][319]<=0;WeightsStore[6][320]<=0;WeightsStore[6][321]<=0;WeightsStore[6][322]<=0;WeightsStore[6][323]<=0;WeightsStore[6][324]<=0;WeightsStore[6][325]<=0;WeightsStore[6][326]<=0;WeightsStore[6][327]<=0;WeightsStore[6][328]<=0;WeightsStore[6][329]<=0;WeightsStore[6][330]<=0;WeightsStore[6][331]<=0;WeightsStore[6][332]<=0;WeightsStore[6][333]<=0;WeightsStore[6][334]<=0;WeightsStore[6][335]<=0;WeightsStore[6][336]<=0;WeightsStore[6][337]<=0;WeightsStore[6][338]<=0;WeightsStore[6][339]<=0;WeightsStore[6][340]<=0;WeightsStore[6][341]<=0;WeightsStore[6][342]<=0;WeightsStore[6][343]<=0;WeightsStore[6][344]<=0;WeightsStore[6][345]<=0;WeightsStore[6][346]<=0;WeightsStore[6][347]<=0;WeightsStore[6][348]<=0;WeightsStore[6][349]<=0;WeightsStore[6][350]<=0;WeightsStore[6][351]<=0;WeightsStore[6][352]<=0;WeightsStore[6][353]<=0;WeightsStore[6][354]<=0;WeightsStore[6][355]<=0;WeightsStore[6][356]<=0;WeightsStore[6][357]<=0;WeightsStore[6][358]<=0;WeightsStore[6][359]<=0;WeightsStore[6][360]<=0;WeightsStore[6][361]<=0;WeightsStore[6][362]<=0;WeightsStore[6][363]<=0;WeightsStore[6][364]<=0;WeightsStore[6][365]<=0;WeightsStore[6][366]<=0;WeightsStore[6][367]<=0;WeightsStore[6][368]<=0;WeightsStore[6][369]<=0;WeightsStore[6][370]<=0;WeightsStore[6][371]<=0;WeightsStore[6][372]<=0;WeightsStore[6][373]<=0;WeightsStore[6][374]<=0;WeightsStore[6][375]<=0;WeightsStore[6][376]<=0;WeightsStore[6][377]<=0;WeightsStore[6][378]<=0;WeightsStore[6][379]<=0;WeightsStore[6][380]<=0;WeightsStore[6][381]<=0;WeightsStore[6][382]<=0;WeightsStore[6][383]<=0;WeightsStore[6][384]<=0;WeightsStore[6][385]<=0;WeightsStore[6][386]<=0;WeightsStore[6][387]<=0;WeightsStore[6][388]<=0;WeightsStore[6][389]<=0;WeightsStore[6][390]<=0;WeightsStore[6][391]<=0;WeightsStore[6][392]<=0;WeightsStore[6][393]<=0;WeightsStore[6][394]<=0;WeightsStore[6][395]<=0;WeightsStore[6][396]<=0;WeightsStore[6][397]<=0;WeightsStore[6][398]<=0;WeightsStore[6][399]<=0;WeightsStore[6][400]<=0;WeightsStore[6][401]<=0;WeightsStore[6][402]<=0;WeightsStore[6][403]<=0;WeightsStore[6][404]<=0;WeightsStore[6][405]<=0;WeightsStore[6][406]<=0;WeightsStore[6][407]<=0;WeightsStore[6][408]<=0;WeightsStore[6][409]<=0;WeightsStore[6][410]<=0;WeightsStore[6][411]<=0;WeightsStore[6][412]<=0;WeightsStore[6][413]<=0;WeightsStore[6][414]<=0;WeightsStore[6][415]<=0;WeightsStore[6][416]<=0;WeightsStore[6][417]<=0;WeightsStore[6][418]<=0;WeightsStore[6][419]<=0;WeightsStore[6][420]<=0;WeightsStore[6][421]<=0;WeightsStore[6][422]<=0;WeightsStore[6][423]<=0;WeightsStore[6][424]<=0;WeightsStore[6][425]<=0;WeightsStore[6][426]<=0;WeightsStore[6][427]<=0;WeightsStore[6][428]<=0;WeightsStore[6][429]<=0;WeightsStore[6][430]<=0;WeightsStore[6][431]<=0;WeightsStore[6][432]<=0;WeightsStore[6][433]<=0;WeightsStore[6][434]<=0;WeightsStore[6][435]<=0;WeightsStore[6][436]<=0;WeightsStore[6][437]<=0;WeightsStore[6][438]<=0;WeightsStore[6][439]<=0;WeightsStore[6][440]<=0;WeightsStore[6][441]<=0;WeightsStore[6][442]<=0;WeightsStore[6][443]<=0;WeightsStore[6][444]<=0;WeightsStore[6][445]<=0;WeightsStore[6][446]<=0;WeightsStore[6][447]<=0;WeightsStore[6][448]<=0;WeightsStore[6][449]<=0;WeightsStore[6][450]<=0;WeightsStore[6][451]<=0;WeightsStore[6][452]<=0;WeightsStore[6][453]<=0;WeightsStore[6][454]<=0;WeightsStore[6][455]<=0;WeightsStore[6][456]<=0;WeightsStore[6][457]<=0;WeightsStore[6][458]<=0;WeightsStore[6][459]<=0;WeightsStore[6][460]<=0;WeightsStore[6][461]<=0;WeightsStore[6][462]<=0;WeightsStore[6][463]<=0;WeightsStore[6][464]<=0;WeightsStore[6][465]<=0;WeightsStore[6][466]<=0;WeightsStore[6][467]<=0;WeightsStore[6][468]<=0;WeightsStore[6][469]<=0;WeightsStore[6][470]<=0;WeightsStore[6][471]<=0;WeightsStore[6][472]<=0;WeightsStore[6][473]<=0;WeightsStore[6][474]<=0;WeightsStore[6][475]<=0;WeightsStore[6][476]<=0;WeightsStore[6][477]<=0;WeightsStore[6][478]<=0;WeightsStore[6][479]<=0;WeightsStore[6][480]<=0;WeightsStore[6][481]<=0;WeightsStore[6][482]<=0;WeightsStore[6][483]<=0;WeightsStore[6][484]<=0;WeightsStore[6][485]<=0;WeightsStore[6][486]<=0;WeightsStore[6][487]<=0;WeightsStore[6][488]<=0;WeightsStore[6][489]<=0;WeightsStore[6][490]<=0;WeightsStore[6][491]<=0;WeightsStore[6][492]<=0;WeightsStore[6][493]<=0;WeightsStore[6][494]<=0;WeightsStore[6][495]<=0;WeightsStore[6][496]<=0;WeightsStore[6][497]<=0;WeightsStore[6][498]<=0;WeightsStore[6][499]<=0;WeightsStore[6][500]<=0;WeightsStore[6][501]<=0;WeightsStore[6][502]<=0;WeightsStore[6][503]<=0;WeightsStore[6][504]<=0;WeightsStore[6][505]<=0;WeightsStore[6][506]<=0;WeightsStore[6][507]<=0;WeightsStore[6][508]<=0;WeightsStore[6][509]<=0;WeightsStore[6][510]<=0;WeightsStore[6][511]<=0;WeightsStore[6][512]<=0;WeightsStore[6][513]<=0;WeightsStore[6][514]<=0;WeightsStore[6][515]<=0;WeightsStore[6][516]<=0;WeightsStore[6][517]<=0;WeightsStore[6][518]<=0;WeightsStore[6][519]<=0;WeightsStore[6][520]<=0;WeightsStore[6][521]<=0;WeightsStore[6][522]<=0;WeightsStore[6][523]<=0;WeightsStore[6][524]<=0;WeightsStore[6][525]<=0;WeightsStore[6][526]<=0;WeightsStore[6][527]<=0;WeightsStore[6][528]<=0;WeightsStore[6][529]<=0;WeightsStore[6][530]<=0;WeightsStore[6][531]<=0;WeightsStore[6][532]<=0;WeightsStore[6][533]<=0;WeightsStore[6][534]<=0;WeightsStore[6][535]<=0;WeightsStore[6][536]<=0;WeightsStore[6][537]<=0;WeightsStore[6][538]<=0;WeightsStore[6][539]<=0;WeightsStore[6][540]<=0;WeightsStore[6][541]<=0;WeightsStore[6][542]<=0;WeightsStore[6][543]<=0;WeightsStore[6][544]<=0;WeightsStore[6][545]<=0;WeightsStore[6][546]<=0;WeightsStore[6][547]<=0;WeightsStore[6][548]<=0;WeightsStore[6][549]<=0;WeightsStore[6][550]<=0;WeightsStore[6][551]<=0;WeightsStore[6][552]<=0;WeightsStore[6][553]<=0;WeightsStore[6][554]<=0;WeightsStore[6][555]<=0;WeightsStore[6][556]<=0;WeightsStore[6][557]<=0;WeightsStore[6][558]<=0;WeightsStore[6][559]<=0;WeightsStore[6][560]<=0;WeightsStore[6][561]<=0;WeightsStore[6][562]<=0;WeightsStore[6][563]<=0;WeightsStore[6][564]<=0;WeightsStore[6][565]<=0;WeightsStore[6][566]<=0;WeightsStore[6][567]<=0;WeightsStore[6][568]<=0;WeightsStore[6][569]<=0;WeightsStore[6][570]<=0;WeightsStore[6][571]<=0;WeightsStore[6][572]<=0;WeightsStore[6][573]<=0;WeightsStore[6][574]<=0;WeightsStore[6][575]<=0;WeightsStore[6][576]<=0;WeightsStore[6][577]<=0;WeightsStore[6][578]<=0;WeightsStore[6][579]<=0;WeightsStore[6][580]<=0;WeightsStore[6][581]<=0;WeightsStore[6][582]<=0;WeightsStore[6][583]<=0;WeightsStore[6][584]<=0;WeightsStore[6][585]<=0;WeightsStore[6][586]<=0;WeightsStore[6][587]<=0;WeightsStore[6][588]<=0;WeightsStore[6][589]<=0;WeightsStore[6][590]<=0;WeightsStore[6][591]<=0;WeightsStore[6][592]<=0;WeightsStore[6][593]<=0;WeightsStore[6][594]<=0;WeightsStore[6][595]<=0;WeightsStore[6][596]<=0;WeightsStore[6][597]<=0;WeightsStore[6][598]<=0;WeightsStore[6][599]<=0;WeightsStore[6][600]<=0;WeightsStore[6][601]<=0;WeightsStore[6][602]<=0;WeightsStore[6][603]<=0;WeightsStore[6][604]<=0;WeightsStore[6][605]<=0;WeightsStore[6][606]<=0;WeightsStore[6][607]<=0;WeightsStore[6][608]<=0;WeightsStore[6][609]<=0;WeightsStore[6][610]<=0;WeightsStore[6][611]<=0;WeightsStore[6][612]<=0;WeightsStore[6][613]<=0;WeightsStore[6][614]<=0;WeightsStore[6][615]<=0;WeightsStore[6][616]<=0;WeightsStore[6][617]<=0;WeightsStore[6][618]<=0;WeightsStore[6][619]<=0;WeightsStore[6][620]<=0;WeightsStore[6][621]<=0;WeightsStore[6][622]<=0;WeightsStore[6][623]<=0;WeightsStore[6][624]<=0;WeightsStore[6][625]<=0;WeightsStore[6][626]<=0;WeightsStore[6][627]<=0;WeightsStore[6][628]<=0;WeightsStore[6][629]<=0;WeightsStore[6][630]<=0;WeightsStore[6][631]<=0;WeightsStore[6][632]<=0;WeightsStore[6][633]<=0;WeightsStore[6][634]<=0;WeightsStore[6][635]<=0;WeightsStore[6][636]<=0;WeightsStore[6][637]<=0;WeightsStore[6][638]<=0;WeightsStore[6][639]<=0;WeightsStore[6][640]<=0;WeightsStore[6][641]<=0;WeightsStore[6][642]<=0;WeightsStore[6][643]<=0;WeightsStore[6][644]<=0;WeightsStore[6][645]<=0;WeightsStore[6][646]<=0;WeightsStore[6][647]<=0;WeightsStore[6][648]<=0;WeightsStore[6][649]<=0;WeightsStore[6][650]<=0;WeightsStore[6][651]<=0;WeightsStore[6][652]<=0;WeightsStore[6][653]<=0;WeightsStore[6][654]<=0;WeightsStore[6][655]<=0;WeightsStore[6][656]<=0;WeightsStore[6][657]<=0;WeightsStore[6][658]<=0;WeightsStore[6][659]<=0;WeightsStore[6][660]<=0;WeightsStore[6][661]<=0;WeightsStore[6][662]<=0;WeightsStore[6][663]<=0;WeightsStore[6][664]<=0;WeightsStore[6][665]<=0;WeightsStore[6][666]<=0;WeightsStore[6][667]<=0;WeightsStore[6][668]<=0;WeightsStore[6][669]<=0;WeightsStore[6][670]<=0;WeightsStore[6][671]<=0;WeightsStore[6][672]<=0;WeightsStore[6][673]<=0;WeightsStore[6][674]<=0;WeightsStore[6][675]<=0;WeightsStore[6][676]<=0;WeightsStore[6][677]<=0;WeightsStore[6][678]<=0;WeightsStore[6][679]<=0;WeightsStore[6][680]<=0;WeightsStore[6][681]<=0;WeightsStore[6][682]<=0;WeightsStore[6][683]<=0;WeightsStore[6][684]<=0;WeightsStore[6][685]<=0;WeightsStore[6][686]<=0;WeightsStore[6][687]<=0;WeightsStore[6][688]<=0;WeightsStore[6][689]<=0;WeightsStore[6][690]<=0;WeightsStore[6][691]<=0;WeightsStore[6][692]<=0;WeightsStore[6][693]<=0;WeightsStore[6][694]<=0;WeightsStore[6][695]<=0;WeightsStore[6][696]<=0;WeightsStore[6][697]<=0;WeightsStore[6][698]<=0;WeightsStore[6][699]<=0;WeightsStore[6][700]<=0;WeightsStore[6][701]<=0;WeightsStore[6][702]<=0;WeightsStore[6][703]<=0;WeightsStore[6][704]<=0;WeightsStore[6][705]<=0;WeightsStore[6][706]<=0;WeightsStore[6][707]<=0;WeightsStore[6][708]<=0;WeightsStore[6][709]<=0;WeightsStore[6][710]<=0;WeightsStore[6][711]<=0;WeightsStore[6][712]<=0;WeightsStore[6][713]<=0;WeightsStore[6][714]<=0;WeightsStore[6][715]<=0;WeightsStore[6][716]<=0;WeightsStore[6][717]<=0;WeightsStore[6][718]<=0;WeightsStore[6][719]<=0;WeightsStore[6][720]<=0;WeightsStore[6][721]<=0;WeightsStore[6][722]<=0;WeightsStore[6][723]<=0;WeightsStore[6][724]<=0;WeightsStore[6][725]<=0;WeightsStore[6][726]<=0;WeightsStore[6][727]<=0;WeightsStore[6][728]<=0;WeightsStore[6][729]<=0;WeightsStore[6][730]<=0;WeightsStore[6][731]<=0;WeightsStore[6][732]<=0;WeightsStore[6][733]<=0;WeightsStore[6][734]<=0;WeightsStore[6][735]<=0;WeightsStore[6][736]<=0;WeightsStore[6][737]<=0;WeightsStore[6][738]<=0;WeightsStore[6][739]<=0;WeightsStore[6][740]<=0;WeightsStore[6][741]<=0;WeightsStore[6][742]<=0;WeightsStore[6][743]<=0;WeightsStore[6][744]<=0;WeightsStore[6][745]<=0;WeightsStore[6][746]<=0;WeightsStore[6][747]<=0;WeightsStore[6][748]<=0;WeightsStore[6][749]<=0;WeightsStore[6][750]<=0;WeightsStore[6][751]<=0;WeightsStore[6][752]<=0;WeightsStore[6][753]<=0;WeightsStore[6][754]<=0;WeightsStore[6][755]<=0;WeightsStore[6][756]<=0;WeightsStore[6][757]<=0;WeightsStore[6][758]<=0;WeightsStore[6][759]<=0;WeightsStore[6][760]<=0;WeightsStore[6][761]<=0;WeightsStore[6][762]<=0;WeightsStore[6][763]<=0;WeightsStore[6][764]<=0;WeightsStore[6][765]<=0;WeightsStore[6][766]<=0;WeightsStore[6][767]<=0;WeightsStore[6][768]<=0;WeightsStore[6][769]<=0;WeightsStore[6][770]<=0;WeightsStore[6][771]<=0;WeightsStore[6][772]<=0;WeightsStore[6][773]<=0;WeightsStore[6][774]<=0;WeightsStore[6][775]<=0;WeightsStore[6][776]<=0;WeightsStore[6][777]<=0;WeightsStore[6][778]<=0;WeightsStore[6][779]<=0;WeightsStore[6][780]<=0;WeightsStore[6][781]<=0;WeightsStore[6][782]<=0;WeightsStore[6][783]<=0;WeightsStore[6][784]<=0;WeightsStore[7][0]<=0;WeightsStore[7][1]<=0;WeightsStore[7][2]<=0;WeightsStore[7][3]<=0;WeightsStore[7][4]<=0;WeightsStore[7][5]<=0;WeightsStore[7][6]<=0;WeightsStore[7][7]<=0;WeightsStore[7][8]<=0;WeightsStore[7][9]<=0;WeightsStore[7][10]<=0;WeightsStore[7][11]<=0;WeightsStore[7][12]<=0;WeightsStore[7][13]<=0;WeightsStore[7][14]<=0;WeightsStore[7][15]<=0;WeightsStore[7][16]<=0;WeightsStore[7][17]<=0;WeightsStore[7][18]<=0;WeightsStore[7][19]<=0;WeightsStore[7][20]<=0;WeightsStore[7][21]<=0;WeightsStore[7][22]<=0;WeightsStore[7][23]<=0;WeightsStore[7][24]<=0;WeightsStore[7][25]<=0;WeightsStore[7][26]<=0;WeightsStore[7][27]<=0;WeightsStore[7][28]<=0;WeightsStore[7][29]<=0;WeightsStore[7][30]<=0;WeightsStore[7][31]<=0;WeightsStore[7][32]<=0;WeightsStore[7][33]<=0;WeightsStore[7][34]<=0;WeightsStore[7][35]<=0;WeightsStore[7][36]<=0;WeightsStore[7][37]<=0;WeightsStore[7][38]<=0;WeightsStore[7][39]<=0;WeightsStore[7][40]<=0;WeightsStore[7][41]<=0;WeightsStore[7][42]<=0;WeightsStore[7][43]<=0;WeightsStore[7][44]<=0;WeightsStore[7][45]<=0;WeightsStore[7][46]<=0;WeightsStore[7][47]<=0;WeightsStore[7][48]<=0;WeightsStore[7][49]<=0;WeightsStore[7][50]<=0;WeightsStore[7][51]<=0;WeightsStore[7][52]<=0;WeightsStore[7][53]<=0;WeightsStore[7][54]<=0;WeightsStore[7][55]<=0;WeightsStore[7][56]<=0;WeightsStore[7][57]<=0;WeightsStore[7][58]<=0;WeightsStore[7][59]<=0;WeightsStore[7][60]<=0;WeightsStore[7][61]<=0;WeightsStore[7][62]<=0;WeightsStore[7][63]<=0;WeightsStore[7][64]<=0;WeightsStore[7][65]<=0;WeightsStore[7][66]<=0;WeightsStore[7][67]<=0;WeightsStore[7][68]<=0;WeightsStore[7][69]<=0;WeightsStore[7][70]<=0;WeightsStore[7][71]<=0;WeightsStore[7][72]<=0;WeightsStore[7][73]<=0;WeightsStore[7][74]<=0;WeightsStore[7][75]<=0;WeightsStore[7][76]<=0;WeightsStore[7][77]<=0;WeightsStore[7][78]<=0;WeightsStore[7][79]<=0;WeightsStore[7][80]<=0;WeightsStore[7][81]<=0;WeightsStore[7][82]<=0;WeightsStore[7][83]<=0;WeightsStore[7][84]<=0;WeightsStore[7][85]<=0;WeightsStore[7][86]<=0;WeightsStore[7][87]<=0;WeightsStore[7][88]<=0;WeightsStore[7][89]<=0;WeightsStore[7][90]<=0;WeightsStore[7][91]<=0;WeightsStore[7][92]<=0;WeightsStore[7][93]<=0;WeightsStore[7][94]<=0;WeightsStore[7][95]<=0;WeightsStore[7][96]<=0;WeightsStore[7][97]<=0;WeightsStore[7][98]<=0;WeightsStore[7][99]<=0;WeightsStore[7][100]<=0;WeightsStore[7][101]<=0;WeightsStore[7][102]<=0;WeightsStore[7][103]<=0;WeightsStore[7][104]<=0;WeightsStore[7][105]<=0;WeightsStore[7][106]<=0;WeightsStore[7][107]<=0;WeightsStore[7][108]<=0;WeightsStore[7][109]<=0;WeightsStore[7][110]<=0;WeightsStore[7][111]<=0;WeightsStore[7][112]<=0;WeightsStore[7][113]<=0;WeightsStore[7][114]<=0;WeightsStore[7][115]<=0;WeightsStore[7][116]<=0;WeightsStore[7][117]<=0;WeightsStore[7][118]<=0;WeightsStore[7][119]<=0;WeightsStore[7][120]<=0;WeightsStore[7][121]<=0;WeightsStore[7][122]<=0;WeightsStore[7][123]<=0;WeightsStore[7][124]<=0;WeightsStore[7][125]<=0;WeightsStore[7][126]<=0;WeightsStore[7][127]<=0;WeightsStore[7][128]<=0;WeightsStore[7][129]<=0;WeightsStore[7][130]<=0;WeightsStore[7][131]<=0;WeightsStore[7][132]<=0;WeightsStore[7][133]<=0;WeightsStore[7][134]<=0;WeightsStore[7][135]<=0;WeightsStore[7][136]<=0;WeightsStore[7][137]<=0;WeightsStore[7][138]<=0;WeightsStore[7][139]<=0;WeightsStore[7][140]<=0;WeightsStore[7][141]<=0;WeightsStore[7][142]<=0;WeightsStore[7][143]<=0;WeightsStore[7][144]<=0;WeightsStore[7][145]<=0;WeightsStore[7][146]<=0;WeightsStore[7][147]<=0;WeightsStore[7][148]<=0;WeightsStore[7][149]<=0;WeightsStore[7][150]<=0;WeightsStore[7][151]<=0;WeightsStore[7][152]<=0;WeightsStore[7][153]<=0;WeightsStore[7][154]<=0;WeightsStore[7][155]<=0;WeightsStore[7][156]<=0;WeightsStore[7][157]<=0;WeightsStore[7][158]<=0;WeightsStore[7][159]<=0;WeightsStore[7][160]<=0;WeightsStore[7][161]<=0;WeightsStore[7][162]<=0;WeightsStore[7][163]<=0;WeightsStore[7][164]<=0;WeightsStore[7][165]<=0;WeightsStore[7][166]<=0;WeightsStore[7][167]<=0;WeightsStore[7][168]<=0;WeightsStore[7][169]<=0;WeightsStore[7][170]<=0;WeightsStore[7][171]<=0;WeightsStore[7][172]<=0;WeightsStore[7][173]<=0;WeightsStore[7][174]<=0;WeightsStore[7][175]<=0;WeightsStore[7][176]<=0;WeightsStore[7][177]<=0;WeightsStore[7][178]<=0;WeightsStore[7][179]<=0;WeightsStore[7][180]<=0;WeightsStore[7][181]<=0;WeightsStore[7][182]<=0;WeightsStore[7][183]<=0;WeightsStore[7][184]<=0;WeightsStore[7][185]<=0;WeightsStore[7][186]<=0;WeightsStore[7][187]<=0;WeightsStore[7][188]<=0;WeightsStore[7][189]<=0;WeightsStore[7][190]<=0;WeightsStore[7][191]<=0;WeightsStore[7][192]<=0;WeightsStore[7][193]<=0;WeightsStore[7][194]<=0;WeightsStore[7][195]<=0;WeightsStore[7][196]<=0;WeightsStore[7][197]<=0;WeightsStore[7][198]<=0;WeightsStore[7][199]<=0;WeightsStore[7][200]<=0;WeightsStore[7][201]<=0;WeightsStore[7][202]<=0;WeightsStore[7][203]<=0;WeightsStore[7][204]<=0;WeightsStore[7][205]<=0;WeightsStore[7][206]<=0;WeightsStore[7][207]<=0;WeightsStore[7][208]<=0;WeightsStore[7][209]<=0;WeightsStore[7][210]<=0;WeightsStore[7][211]<=0;WeightsStore[7][212]<=0;WeightsStore[7][213]<=0;WeightsStore[7][214]<=0;WeightsStore[7][215]<=0;WeightsStore[7][216]<=0;WeightsStore[7][217]<=0;WeightsStore[7][218]<=0;WeightsStore[7][219]<=0;WeightsStore[7][220]<=0;WeightsStore[7][221]<=0;WeightsStore[7][222]<=0;WeightsStore[7][223]<=0;WeightsStore[7][224]<=0;WeightsStore[7][225]<=0;WeightsStore[7][226]<=0;WeightsStore[7][227]<=0;WeightsStore[7][228]<=0;WeightsStore[7][229]<=0;WeightsStore[7][230]<=0;WeightsStore[7][231]<=0;WeightsStore[7][232]<=0;WeightsStore[7][233]<=0;WeightsStore[7][234]<=0;WeightsStore[7][235]<=0;WeightsStore[7][236]<=0;WeightsStore[7][237]<=0;WeightsStore[7][238]<=0;WeightsStore[7][239]<=0;WeightsStore[7][240]<=0;WeightsStore[7][241]<=0;WeightsStore[7][242]<=0;WeightsStore[7][243]<=0;WeightsStore[7][244]<=0;WeightsStore[7][245]<=0;WeightsStore[7][246]<=0;WeightsStore[7][247]<=0;WeightsStore[7][248]<=0;WeightsStore[7][249]<=0;WeightsStore[7][250]<=0;WeightsStore[7][251]<=0;WeightsStore[7][252]<=0;WeightsStore[7][253]<=0;WeightsStore[7][254]<=0;WeightsStore[7][255]<=0;WeightsStore[7][256]<=0;WeightsStore[7][257]<=0;WeightsStore[7][258]<=0;WeightsStore[7][259]<=0;WeightsStore[7][260]<=0;WeightsStore[7][261]<=0;WeightsStore[7][262]<=0;WeightsStore[7][263]<=0;WeightsStore[7][264]<=0;WeightsStore[7][265]<=0;WeightsStore[7][266]<=0;WeightsStore[7][267]<=0;WeightsStore[7][268]<=0;WeightsStore[7][269]<=0;WeightsStore[7][270]<=0;WeightsStore[7][271]<=0;WeightsStore[7][272]<=0;WeightsStore[7][273]<=0;WeightsStore[7][274]<=0;WeightsStore[7][275]<=0;WeightsStore[7][276]<=0;WeightsStore[7][277]<=0;WeightsStore[7][278]<=0;WeightsStore[7][279]<=0;WeightsStore[7][280]<=0;WeightsStore[7][281]<=0;WeightsStore[7][282]<=0;WeightsStore[7][283]<=0;WeightsStore[7][284]<=0;WeightsStore[7][285]<=0;WeightsStore[7][286]<=0;WeightsStore[7][287]<=0;WeightsStore[7][288]<=0;WeightsStore[7][289]<=0;WeightsStore[7][290]<=0;WeightsStore[7][291]<=0;WeightsStore[7][292]<=0;WeightsStore[7][293]<=0;WeightsStore[7][294]<=0;WeightsStore[7][295]<=0;WeightsStore[7][296]<=0;WeightsStore[7][297]<=0;WeightsStore[7][298]<=0;WeightsStore[7][299]<=0;WeightsStore[7][300]<=0;WeightsStore[7][301]<=0;WeightsStore[7][302]<=0;WeightsStore[7][303]<=0;WeightsStore[7][304]<=0;WeightsStore[7][305]<=0;WeightsStore[7][306]<=0;WeightsStore[7][307]<=0;WeightsStore[7][308]<=0;WeightsStore[7][309]<=0;WeightsStore[7][310]<=0;WeightsStore[7][311]<=0;WeightsStore[7][312]<=0;WeightsStore[7][313]<=0;WeightsStore[7][314]<=0;WeightsStore[7][315]<=0;WeightsStore[7][316]<=0;WeightsStore[7][317]<=0;WeightsStore[7][318]<=0;WeightsStore[7][319]<=0;WeightsStore[7][320]<=0;WeightsStore[7][321]<=0;WeightsStore[7][322]<=0;WeightsStore[7][323]<=0;WeightsStore[7][324]<=0;WeightsStore[7][325]<=0;WeightsStore[7][326]<=0;WeightsStore[7][327]<=0;WeightsStore[7][328]<=0;WeightsStore[7][329]<=0;WeightsStore[7][330]<=0;WeightsStore[7][331]<=0;WeightsStore[7][332]<=0;WeightsStore[7][333]<=0;WeightsStore[7][334]<=0;WeightsStore[7][335]<=0;WeightsStore[7][336]<=0;WeightsStore[7][337]<=0;WeightsStore[7][338]<=0;WeightsStore[7][339]<=0;WeightsStore[7][340]<=0;WeightsStore[7][341]<=0;WeightsStore[7][342]<=0;WeightsStore[7][343]<=0;WeightsStore[7][344]<=0;WeightsStore[7][345]<=0;WeightsStore[7][346]<=0;WeightsStore[7][347]<=0;WeightsStore[7][348]<=0;WeightsStore[7][349]<=0;WeightsStore[7][350]<=0;WeightsStore[7][351]<=0;WeightsStore[7][352]<=0;WeightsStore[7][353]<=0;WeightsStore[7][354]<=0;WeightsStore[7][355]<=0;WeightsStore[7][356]<=0;WeightsStore[7][357]<=0;WeightsStore[7][358]<=0;WeightsStore[7][359]<=0;WeightsStore[7][360]<=0;WeightsStore[7][361]<=0;WeightsStore[7][362]<=0;WeightsStore[7][363]<=0;WeightsStore[7][364]<=0;WeightsStore[7][365]<=0;WeightsStore[7][366]<=0;WeightsStore[7][367]<=0;WeightsStore[7][368]<=0;WeightsStore[7][369]<=0;WeightsStore[7][370]<=0;WeightsStore[7][371]<=0;WeightsStore[7][372]<=0;WeightsStore[7][373]<=0;WeightsStore[7][374]<=0;WeightsStore[7][375]<=0;WeightsStore[7][376]<=0;WeightsStore[7][377]<=0;WeightsStore[7][378]<=0;WeightsStore[7][379]<=0;WeightsStore[7][380]<=0;WeightsStore[7][381]<=0;WeightsStore[7][382]<=0;WeightsStore[7][383]<=0;WeightsStore[7][384]<=0;WeightsStore[7][385]<=0;WeightsStore[7][386]<=0;WeightsStore[7][387]<=0;WeightsStore[7][388]<=0;WeightsStore[7][389]<=0;WeightsStore[7][390]<=0;WeightsStore[7][391]<=0;WeightsStore[7][392]<=0;WeightsStore[7][393]<=0;WeightsStore[7][394]<=0;WeightsStore[7][395]<=0;WeightsStore[7][396]<=0;WeightsStore[7][397]<=0;WeightsStore[7][398]<=0;WeightsStore[7][399]<=0;WeightsStore[7][400]<=0;WeightsStore[7][401]<=0;WeightsStore[7][402]<=0;WeightsStore[7][403]<=0;WeightsStore[7][404]<=0;WeightsStore[7][405]<=0;WeightsStore[7][406]<=0;WeightsStore[7][407]<=0;WeightsStore[7][408]<=0;WeightsStore[7][409]<=0;WeightsStore[7][410]<=0;WeightsStore[7][411]<=0;WeightsStore[7][412]<=0;WeightsStore[7][413]<=0;WeightsStore[7][414]<=0;WeightsStore[7][415]<=0;WeightsStore[7][416]<=0;WeightsStore[7][417]<=0;WeightsStore[7][418]<=0;WeightsStore[7][419]<=0;WeightsStore[7][420]<=0;WeightsStore[7][421]<=0;WeightsStore[7][422]<=0;WeightsStore[7][423]<=0;WeightsStore[7][424]<=0;WeightsStore[7][425]<=0;WeightsStore[7][426]<=0;WeightsStore[7][427]<=0;WeightsStore[7][428]<=0;WeightsStore[7][429]<=0;WeightsStore[7][430]<=0;WeightsStore[7][431]<=0;WeightsStore[7][432]<=0;WeightsStore[7][433]<=0;WeightsStore[7][434]<=0;WeightsStore[7][435]<=0;WeightsStore[7][436]<=0;WeightsStore[7][437]<=0;WeightsStore[7][438]<=0;WeightsStore[7][439]<=0;WeightsStore[7][440]<=0;WeightsStore[7][441]<=0;WeightsStore[7][442]<=0;WeightsStore[7][443]<=0;WeightsStore[7][444]<=0;WeightsStore[7][445]<=0;WeightsStore[7][446]<=0;WeightsStore[7][447]<=0;WeightsStore[7][448]<=0;WeightsStore[7][449]<=0;WeightsStore[7][450]<=0;WeightsStore[7][451]<=0;WeightsStore[7][452]<=0;WeightsStore[7][453]<=0;WeightsStore[7][454]<=0;WeightsStore[7][455]<=0;WeightsStore[7][456]<=0;WeightsStore[7][457]<=0;WeightsStore[7][458]<=0;WeightsStore[7][459]<=0;WeightsStore[7][460]<=0;WeightsStore[7][461]<=0;WeightsStore[7][462]<=0;WeightsStore[7][463]<=0;WeightsStore[7][464]<=0;WeightsStore[7][465]<=0;WeightsStore[7][466]<=0;WeightsStore[7][467]<=0;WeightsStore[7][468]<=0;WeightsStore[7][469]<=0;WeightsStore[7][470]<=0;WeightsStore[7][471]<=0;WeightsStore[7][472]<=0;WeightsStore[7][473]<=0;WeightsStore[7][474]<=0;WeightsStore[7][475]<=0;WeightsStore[7][476]<=0;WeightsStore[7][477]<=0;WeightsStore[7][478]<=0;WeightsStore[7][479]<=0;WeightsStore[7][480]<=0;WeightsStore[7][481]<=0;WeightsStore[7][482]<=0;WeightsStore[7][483]<=0;WeightsStore[7][484]<=0;WeightsStore[7][485]<=0;WeightsStore[7][486]<=0;WeightsStore[7][487]<=0;WeightsStore[7][488]<=0;WeightsStore[7][489]<=0;WeightsStore[7][490]<=0;WeightsStore[7][491]<=0;WeightsStore[7][492]<=0;WeightsStore[7][493]<=0;WeightsStore[7][494]<=0;WeightsStore[7][495]<=0;WeightsStore[7][496]<=0;WeightsStore[7][497]<=0;WeightsStore[7][498]<=0;WeightsStore[7][499]<=0;WeightsStore[7][500]<=0;WeightsStore[7][501]<=0;WeightsStore[7][502]<=0;WeightsStore[7][503]<=0;WeightsStore[7][504]<=0;WeightsStore[7][505]<=0;WeightsStore[7][506]<=0;WeightsStore[7][507]<=0;WeightsStore[7][508]<=0;WeightsStore[7][509]<=0;WeightsStore[7][510]<=0;WeightsStore[7][511]<=0;WeightsStore[7][512]<=0;WeightsStore[7][513]<=0;WeightsStore[7][514]<=0;WeightsStore[7][515]<=0;WeightsStore[7][516]<=0;WeightsStore[7][517]<=0;WeightsStore[7][518]<=0;WeightsStore[7][519]<=0;WeightsStore[7][520]<=0;WeightsStore[7][521]<=0;WeightsStore[7][522]<=0;WeightsStore[7][523]<=0;WeightsStore[7][524]<=0;WeightsStore[7][525]<=0;WeightsStore[7][526]<=0;WeightsStore[7][527]<=0;WeightsStore[7][528]<=0;WeightsStore[7][529]<=0;WeightsStore[7][530]<=0;WeightsStore[7][531]<=0;WeightsStore[7][532]<=0;WeightsStore[7][533]<=0;WeightsStore[7][534]<=0;WeightsStore[7][535]<=0;WeightsStore[7][536]<=0;WeightsStore[7][537]<=0;WeightsStore[7][538]<=0;WeightsStore[7][539]<=0;WeightsStore[7][540]<=0;WeightsStore[7][541]<=0;WeightsStore[7][542]<=0;WeightsStore[7][543]<=0;WeightsStore[7][544]<=0;WeightsStore[7][545]<=0;WeightsStore[7][546]<=0;WeightsStore[7][547]<=0;WeightsStore[7][548]<=0;WeightsStore[7][549]<=0;WeightsStore[7][550]<=0;WeightsStore[7][551]<=0;WeightsStore[7][552]<=0;WeightsStore[7][553]<=0;WeightsStore[7][554]<=0;WeightsStore[7][555]<=0;WeightsStore[7][556]<=0;WeightsStore[7][557]<=0;WeightsStore[7][558]<=0;WeightsStore[7][559]<=0;WeightsStore[7][560]<=0;WeightsStore[7][561]<=0;WeightsStore[7][562]<=0;WeightsStore[7][563]<=0;WeightsStore[7][564]<=0;WeightsStore[7][565]<=0;WeightsStore[7][566]<=0;WeightsStore[7][567]<=0;WeightsStore[7][568]<=0;WeightsStore[7][569]<=0;WeightsStore[7][570]<=0;WeightsStore[7][571]<=0;WeightsStore[7][572]<=0;WeightsStore[7][573]<=0;WeightsStore[7][574]<=0;WeightsStore[7][575]<=0;WeightsStore[7][576]<=0;WeightsStore[7][577]<=0;WeightsStore[7][578]<=0;WeightsStore[7][579]<=0;WeightsStore[7][580]<=0;WeightsStore[7][581]<=0;WeightsStore[7][582]<=0;WeightsStore[7][583]<=0;WeightsStore[7][584]<=0;WeightsStore[7][585]<=0;WeightsStore[7][586]<=0;WeightsStore[7][587]<=0;WeightsStore[7][588]<=0;WeightsStore[7][589]<=0;WeightsStore[7][590]<=0;WeightsStore[7][591]<=0;WeightsStore[7][592]<=0;WeightsStore[7][593]<=0;WeightsStore[7][594]<=0;WeightsStore[7][595]<=0;WeightsStore[7][596]<=0;WeightsStore[7][597]<=0;WeightsStore[7][598]<=0;WeightsStore[7][599]<=0;WeightsStore[7][600]<=0;WeightsStore[7][601]<=0;WeightsStore[7][602]<=0;WeightsStore[7][603]<=0;WeightsStore[7][604]<=0;WeightsStore[7][605]<=0;WeightsStore[7][606]<=0;WeightsStore[7][607]<=0;WeightsStore[7][608]<=0;WeightsStore[7][609]<=0;WeightsStore[7][610]<=0;WeightsStore[7][611]<=0;WeightsStore[7][612]<=0;WeightsStore[7][613]<=0;WeightsStore[7][614]<=0;WeightsStore[7][615]<=0;WeightsStore[7][616]<=0;WeightsStore[7][617]<=0;WeightsStore[7][618]<=0;WeightsStore[7][619]<=0;WeightsStore[7][620]<=0;WeightsStore[7][621]<=0;WeightsStore[7][622]<=0;WeightsStore[7][623]<=0;WeightsStore[7][624]<=0;WeightsStore[7][625]<=0;WeightsStore[7][626]<=0;WeightsStore[7][627]<=0;WeightsStore[7][628]<=0;WeightsStore[7][629]<=0;WeightsStore[7][630]<=0;WeightsStore[7][631]<=0;WeightsStore[7][632]<=0;WeightsStore[7][633]<=0;WeightsStore[7][634]<=0;WeightsStore[7][635]<=0;WeightsStore[7][636]<=0;WeightsStore[7][637]<=0;WeightsStore[7][638]<=0;WeightsStore[7][639]<=0;WeightsStore[7][640]<=0;WeightsStore[7][641]<=0;WeightsStore[7][642]<=0;WeightsStore[7][643]<=0;WeightsStore[7][644]<=0;WeightsStore[7][645]<=0;WeightsStore[7][646]<=0;WeightsStore[7][647]<=0;WeightsStore[7][648]<=0;WeightsStore[7][649]<=0;WeightsStore[7][650]<=0;WeightsStore[7][651]<=0;WeightsStore[7][652]<=0;WeightsStore[7][653]<=0;WeightsStore[7][654]<=0;WeightsStore[7][655]<=0;WeightsStore[7][656]<=0;WeightsStore[7][657]<=0;WeightsStore[7][658]<=0;WeightsStore[7][659]<=0;WeightsStore[7][660]<=0;WeightsStore[7][661]<=0;WeightsStore[7][662]<=0;WeightsStore[7][663]<=0;WeightsStore[7][664]<=0;WeightsStore[7][665]<=0;WeightsStore[7][666]<=0;WeightsStore[7][667]<=0;WeightsStore[7][668]<=0;WeightsStore[7][669]<=0;WeightsStore[7][670]<=0;WeightsStore[7][671]<=0;WeightsStore[7][672]<=0;WeightsStore[7][673]<=0;WeightsStore[7][674]<=0;WeightsStore[7][675]<=0;WeightsStore[7][676]<=0;WeightsStore[7][677]<=0;WeightsStore[7][678]<=0;WeightsStore[7][679]<=0;WeightsStore[7][680]<=0;WeightsStore[7][681]<=0;WeightsStore[7][682]<=0;WeightsStore[7][683]<=0;WeightsStore[7][684]<=0;WeightsStore[7][685]<=0;WeightsStore[7][686]<=0;WeightsStore[7][687]<=0;WeightsStore[7][688]<=0;WeightsStore[7][689]<=0;WeightsStore[7][690]<=0;WeightsStore[7][691]<=0;WeightsStore[7][692]<=0;WeightsStore[7][693]<=0;WeightsStore[7][694]<=0;WeightsStore[7][695]<=0;WeightsStore[7][696]<=0;WeightsStore[7][697]<=0;WeightsStore[7][698]<=0;WeightsStore[7][699]<=0;WeightsStore[7][700]<=0;WeightsStore[7][701]<=0;WeightsStore[7][702]<=0;WeightsStore[7][703]<=0;WeightsStore[7][704]<=0;WeightsStore[7][705]<=0;WeightsStore[7][706]<=0;WeightsStore[7][707]<=0;WeightsStore[7][708]<=0;WeightsStore[7][709]<=0;WeightsStore[7][710]<=0;WeightsStore[7][711]<=0;WeightsStore[7][712]<=0;WeightsStore[7][713]<=0;WeightsStore[7][714]<=0;WeightsStore[7][715]<=0;WeightsStore[7][716]<=0;WeightsStore[7][717]<=0;WeightsStore[7][718]<=0;WeightsStore[7][719]<=0;WeightsStore[7][720]<=0;WeightsStore[7][721]<=0;WeightsStore[7][722]<=0;WeightsStore[7][723]<=0;WeightsStore[7][724]<=0;WeightsStore[7][725]<=0;WeightsStore[7][726]<=0;WeightsStore[7][727]<=0;WeightsStore[7][728]<=0;WeightsStore[7][729]<=0;WeightsStore[7][730]<=0;WeightsStore[7][731]<=0;WeightsStore[7][732]<=0;WeightsStore[7][733]<=0;WeightsStore[7][734]<=0;WeightsStore[7][735]<=0;WeightsStore[7][736]<=0;WeightsStore[7][737]<=0;WeightsStore[7][738]<=0;WeightsStore[7][739]<=0;WeightsStore[7][740]<=0;WeightsStore[7][741]<=0;WeightsStore[7][742]<=0;WeightsStore[7][743]<=0;WeightsStore[7][744]<=0;WeightsStore[7][745]<=0;WeightsStore[7][746]<=0;WeightsStore[7][747]<=0;WeightsStore[7][748]<=0;WeightsStore[7][749]<=0;WeightsStore[7][750]<=0;WeightsStore[7][751]<=0;WeightsStore[7][752]<=0;WeightsStore[7][753]<=0;WeightsStore[7][754]<=0;WeightsStore[7][755]<=0;WeightsStore[7][756]<=0;WeightsStore[7][757]<=0;WeightsStore[7][758]<=0;WeightsStore[7][759]<=0;WeightsStore[7][760]<=0;WeightsStore[7][761]<=0;WeightsStore[7][762]<=0;WeightsStore[7][763]<=0;WeightsStore[7][764]<=0;WeightsStore[7][765]<=0;WeightsStore[7][766]<=0;WeightsStore[7][767]<=0;WeightsStore[7][768]<=0;WeightsStore[7][769]<=0;WeightsStore[7][770]<=0;WeightsStore[7][771]<=0;WeightsStore[7][772]<=0;WeightsStore[7][773]<=0;WeightsStore[7][774]<=0;WeightsStore[7][775]<=0;WeightsStore[7][776]<=0;WeightsStore[7][777]<=0;WeightsStore[7][778]<=0;WeightsStore[7][779]<=0;WeightsStore[7][780]<=0;WeightsStore[7][781]<=0;WeightsStore[7][782]<=0;WeightsStore[7][783]<=0;WeightsStore[7][784]<=0;WeightsStore[8][0]<=0;WeightsStore[8][1]<=0;WeightsStore[8][2]<=0;WeightsStore[8][3]<=0;WeightsStore[8][4]<=0;WeightsStore[8][5]<=0;WeightsStore[8][6]<=0;WeightsStore[8][7]<=0;WeightsStore[8][8]<=0;WeightsStore[8][9]<=0;WeightsStore[8][10]<=0;WeightsStore[8][11]<=0;WeightsStore[8][12]<=0;WeightsStore[8][13]<=0;WeightsStore[8][14]<=0;WeightsStore[8][15]<=0;WeightsStore[8][16]<=0;WeightsStore[8][17]<=0;WeightsStore[8][18]<=0;WeightsStore[8][19]<=0;WeightsStore[8][20]<=0;WeightsStore[8][21]<=0;WeightsStore[8][22]<=0;WeightsStore[8][23]<=0;WeightsStore[8][24]<=0;WeightsStore[8][25]<=0;WeightsStore[8][26]<=0;WeightsStore[8][27]<=0;WeightsStore[8][28]<=0;WeightsStore[8][29]<=0;WeightsStore[8][30]<=0;WeightsStore[8][31]<=0;WeightsStore[8][32]<=0;WeightsStore[8][33]<=0;WeightsStore[8][34]<=0;WeightsStore[8][35]<=0;WeightsStore[8][36]<=0;WeightsStore[8][37]<=0;WeightsStore[8][38]<=0;WeightsStore[8][39]<=0;WeightsStore[8][40]<=0;WeightsStore[8][41]<=0;WeightsStore[8][42]<=0;WeightsStore[8][43]<=0;WeightsStore[8][44]<=0;WeightsStore[8][45]<=0;WeightsStore[8][46]<=0;WeightsStore[8][47]<=0;WeightsStore[8][48]<=0;WeightsStore[8][49]<=0;WeightsStore[8][50]<=0;WeightsStore[8][51]<=0;WeightsStore[8][52]<=0;WeightsStore[8][53]<=0;WeightsStore[8][54]<=0;WeightsStore[8][55]<=0;WeightsStore[8][56]<=0;WeightsStore[8][57]<=0;WeightsStore[8][58]<=0;WeightsStore[8][59]<=0;WeightsStore[8][60]<=0;WeightsStore[8][61]<=0;WeightsStore[8][62]<=0;WeightsStore[8][63]<=0;WeightsStore[8][64]<=0;WeightsStore[8][65]<=0;WeightsStore[8][66]<=0;WeightsStore[8][67]<=0;WeightsStore[8][68]<=0;WeightsStore[8][69]<=0;WeightsStore[8][70]<=0;WeightsStore[8][71]<=0;WeightsStore[8][72]<=0;WeightsStore[8][73]<=0;WeightsStore[8][74]<=0;WeightsStore[8][75]<=0;WeightsStore[8][76]<=0;WeightsStore[8][77]<=0;WeightsStore[8][78]<=0;WeightsStore[8][79]<=0;WeightsStore[8][80]<=0;WeightsStore[8][81]<=0;WeightsStore[8][82]<=0;WeightsStore[8][83]<=0;WeightsStore[8][84]<=0;WeightsStore[8][85]<=0;WeightsStore[8][86]<=0;WeightsStore[8][87]<=0;WeightsStore[8][88]<=0;WeightsStore[8][89]<=0;WeightsStore[8][90]<=0;WeightsStore[8][91]<=0;WeightsStore[8][92]<=0;WeightsStore[8][93]<=0;WeightsStore[8][94]<=0;WeightsStore[8][95]<=0;WeightsStore[8][96]<=0;WeightsStore[8][97]<=0;WeightsStore[8][98]<=0;WeightsStore[8][99]<=0;WeightsStore[8][100]<=0;WeightsStore[8][101]<=0;WeightsStore[8][102]<=0;WeightsStore[8][103]<=0;WeightsStore[8][104]<=0;WeightsStore[8][105]<=0;WeightsStore[8][106]<=0;WeightsStore[8][107]<=0;WeightsStore[8][108]<=0;WeightsStore[8][109]<=0;WeightsStore[8][110]<=0;WeightsStore[8][111]<=0;WeightsStore[8][112]<=0;WeightsStore[8][113]<=0;WeightsStore[8][114]<=0;WeightsStore[8][115]<=0;WeightsStore[8][116]<=0;WeightsStore[8][117]<=0;WeightsStore[8][118]<=0;WeightsStore[8][119]<=0;WeightsStore[8][120]<=0;WeightsStore[8][121]<=0;WeightsStore[8][122]<=0;WeightsStore[8][123]<=0;WeightsStore[8][124]<=0;WeightsStore[8][125]<=0;WeightsStore[8][126]<=0;WeightsStore[8][127]<=0;WeightsStore[8][128]<=0;WeightsStore[8][129]<=0;WeightsStore[8][130]<=0;WeightsStore[8][131]<=0;WeightsStore[8][132]<=0;WeightsStore[8][133]<=0;WeightsStore[8][134]<=0;WeightsStore[8][135]<=0;WeightsStore[8][136]<=0;WeightsStore[8][137]<=0;WeightsStore[8][138]<=0;WeightsStore[8][139]<=0;WeightsStore[8][140]<=0;WeightsStore[8][141]<=0;WeightsStore[8][142]<=0;WeightsStore[8][143]<=0;WeightsStore[8][144]<=0;WeightsStore[8][145]<=0;WeightsStore[8][146]<=0;WeightsStore[8][147]<=0;WeightsStore[8][148]<=0;WeightsStore[8][149]<=0;WeightsStore[8][150]<=0;WeightsStore[8][151]<=0;WeightsStore[8][152]<=0;WeightsStore[8][153]<=0;WeightsStore[8][154]<=0;WeightsStore[8][155]<=0;WeightsStore[8][156]<=0;WeightsStore[8][157]<=0;WeightsStore[8][158]<=0;WeightsStore[8][159]<=0;WeightsStore[8][160]<=0;WeightsStore[8][161]<=0;WeightsStore[8][162]<=0;WeightsStore[8][163]<=0;WeightsStore[8][164]<=0;WeightsStore[8][165]<=0;WeightsStore[8][166]<=0;WeightsStore[8][167]<=0;WeightsStore[8][168]<=0;WeightsStore[8][169]<=0;WeightsStore[8][170]<=0;WeightsStore[8][171]<=0;WeightsStore[8][172]<=0;WeightsStore[8][173]<=0;WeightsStore[8][174]<=0;WeightsStore[8][175]<=0;WeightsStore[8][176]<=0;WeightsStore[8][177]<=0;WeightsStore[8][178]<=0;WeightsStore[8][179]<=0;WeightsStore[8][180]<=0;WeightsStore[8][181]<=0;WeightsStore[8][182]<=0;WeightsStore[8][183]<=0;WeightsStore[8][184]<=0;WeightsStore[8][185]<=0;WeightsStore[8][186]<=0;WeightsStore[8][187]<=0;WeightsStore[8][188]<=0;WeightsStore[8][189]<=0;WeightsStore[8][190]<=0;WeightsStore[8][191]<=0;WeightsStore[8][192]<=0;WeightsStore[8][193]<=0;WeightsStore[8][194]<=0;WeightsStore[8][195]<=0;WeightsStore[8][196]<=0;WeightsStore[8][197]<=0;WeightsStore[8][198]<=0;WeightsStore[8][199]<=0;WeightsStore[8][200]<=0;WeightsStore[8][201]<=0;WeightsStore[8][202]<=0;WeightsStore[8][203]<=0;WeightsStore[8][204]<=0;WeightsStore[8][205]<=0;WeightsStore[8][206]<=0;WeightsStore[8][207]<=0;WeightsStore[8][208]<=0;WeightsStore[8][209]<=0;WeightsStore[8][210]<=0;WeightsStore[8][211]<=0;WeightsStore[8][212]<=0;WeightsStore[8][213]<=0;WeightsStore[8][214]<=0;WeightsStore[8][215]<=0;WeightsStore[8][216]<=0;WeightsStore[8][217]<=0;WeightsStore[8][218]<=0;WeightsStore[8][219]<=0;WeightsStore[8][220]<=0;WeightsStore[8][221]<=0;WeightsStore[8][222]<=0;WeightsStore[8][223]<=0;WeightsStore[8][224]<=0;WeightsStore[8][225]<=0;WeightsStore[8][226]<=0;WeightsStore[8][227]<=0;WeightsStore[8][228]<=0;WeightsStore[8][229]<=0;WeightsStore[8][230]<=0;WeightsStore[8][231]<=0;WeightsStore[8][232]<=0;WeightsStore[8][233]<=0;WeightsStore[8][234]<=0;WeightsStore[8][235]<=0;WeightsStore[8][236]<=0;WeightsStore[8][237]<=0;WeightsStore[8][238]<=0;WeightsStore[8][239]<=0;WeightsStore[8][240]<=0;WeightsStore[8][241]<=0;WeightsStore[8][242]<=0;WeightsStore[8][243]<=0;WeightsStore[8][244]<=0;WeightsStore[8][245]<=0;WeightsStore[8][246]<=0;WeightsStore[8][247]<=0;WeightsStore[8][248]<=0;WeightsStore[8][249]<=0;WeightsStore[8][250]<=0;WeightsStore[8][251]<=0;WeightsStore[8][252]<=0;WeightsStore[8][253]<=0;WeightsStore[8][254]<=0;WeightsStore[8][255]<=0;WeightsStore[8][256]<=0;WeightsStore[8][257]<=0;WeightsStore[8][258]<=0;WeightsStore[8][259]<=0;WeightsStore[8][260]<=0;WeightsStore[8][261]<=0;WeightsStore[8][262]<=0;WeightsStore[8][263]<=0;WeightsStore[8][264]<=0;WeightsStore[8][265]<=0;WeightsStore[8][266]<=0;WeightsStore[8][267]<=0;WeightsStore[8][268]<=0;WeightsStore[8][269]<=0;WeightsStore[8][270]<=0;WeightsStore[8][271]<=0;WeightsStore[8][272]<=0;WeightsStore[8][273]<=0;WeightsStore[8][274]<=0;WeightsStore[8][275]<=0;WeightsStore[8][276]<=0;WeightsStore[8][277]<=0;WeightsStore[8][278]<=0;WeightsStore[8][279]<=0;WeightsStore[8][280]<=0;WeightsStore[8][281]<=0;WeightsStore[8][282]<=0;WeightsStore[8][283]<=0;WeightsStore[8][284]<=0;WeightsStore[8][285]<=0;WeightsStore[8][286]<=0;WeightsStore[8][287]<=0;WeightsStore[8][288]<=0;WeightsStore[8][289]<=0;WeightsStore[8][290]<=0;WeightsStore[8][291]<=0;WeightsStore[8][292]<=0;WeightsStore[8][293]<=0;WeightsStore[8][294]<=0;WeightsStore[8][295]<=0;WeightsStore[8][296]<=0;WeightsStore[8][297]<=0;WeightsStore[8][298]<=0;WeightsStore[8][299]<=0;WeightsStore[8][300]<=0;WeightsStore[8][301]<=0;WeightsStore[8][302]<=0;WeightsStore[8][303]<=0;WeightsStore[8][304]<=0;WeightsStore[8][305]<=0;WeightsStore[8][306]<=0;WeightsStore[8][307]<=0;WeightsStore[8][308]<=0;WeightsStore[8][309]<=0;WeightsStore[8][310]<=0;WeightsStore[8][311]<=0;WeightsStore[8][312]<=0;WeightsStore[8][313]<=0;WeightsStore[8][314]<=0;WeightsStore[8][315]<=0;WeightsStore[8][316]<=0;WeightsStore[8][317]<=0;WeightsStore[8][318]<=0;WeightsStore[8][319]<=0;WeightsStore[8][320]<=0;WeightsStore[8][321]<=0;WeightsStore[8][322]<=0;WeightsStore[8][323]<=0;WeightsStore[8][324]<=0;WeightsStore[8][325]<=0;WeightsStore[8][326]<=0;WeightsStore[8][327]<=0;WeightsStore[8][328]<=0;WeightsStore[8][329]<=0;WeightsStore[8][330]<=0;WeightsStore[8][331]<=0;WeightsStore[8][332]<=0;WeightsStore[8][333]<=0;WeightsStore[8][334]<=0;WeightsStore[8][335]<=0;WeightsStore[8][336]<=0;WeightsStore[8][337]<=0;WeightsStore[8][338]<=0;WeightsStore[8][339]<=0;WeightsStore[8][340]<=0;WeightsStore[8][341]<=0;WeightsStore[8][342]<=0;WeightsStore[8][343]<=0;WeightsStore[8][344]<=0;WeightsStore[8][345]<=0;WeightsStore[8][346]<=0;WeightsStore[8][347]<=0;WeightsStore[8][348]<=0;WeightsStore[8][349]<=0;WeightsStore[8][350]<=0;WeightsStore[8][351]<=0;WeightsStore[8][352]<=0;WeightsStore[8][353]<=0;WeightsStore[8][354]<=0;WeightsStore[8][355]<=0;WeightsStore[8][356]<=0;WeightsStore[8][357]<=0;WeightsStore[8][358]<=0;WeightsStore[8][359]<=0;WeightsStore[8][360]<=0;WeightsStore[8][361]<=0;WeightsStore[8][362]<=0;WeightsStore[8][363]<=0;WeightsStore[8][364]<=0;WeightsStore[8][365]<=0;WeightsStore[8][366]<=0;WeightsStore[8][367]<=0;WeightsStore[8][368]<=0;WeightsStore[8][369]<=0;WeightsStore[8][370]<=0;WeightsStore[8][371]<=0;WeightsStore[8][372]<=0;WeightsStore[8][373]<=0;WeightsStore[8][374]<=0;WeightsStore[8][375]<=0;WeightsStore[8][376]<=0;WeightsStore[8][377]<=0;WeightsStore[8][378]<=0;WeightsStore[8][379]<=0;WeightsStore[8][380]<=0;WeightsStore[8][381]<=0;WeightsStore[8][382]<=0;WeightsStore[8][383]<=0;WeightsStore[8][384]<=0;WeightsStore[8][385]<=0;WeightsStore[8][386]<=0;WeightsStore[8][387]<=0;WeightsStore[8][388]<=0;WeightsStore[8][389]<=0;WeightsStore[8][390]<=0;WeightsStore[8][391]<=0;WeightsStore[8][392]<=0;WeightsStore[8][393]<=0;WeightsStore[8][394]<=0;WeightsStore[8][395]<=0;WeightsStore[8][396]<=0;WeightsStore[8][397]<=0;WeightsStore[8][398]<=0;WeightsStore[8][399]<=0;WeightsStore[8][400]<=0;WeightsStore[8][401]<=0;WeightsStore[8][402]<=0;WeightsStore[8][403]<=0;WeightsStore[8][404]<=0;WeightsStore[8][405]<=0;WeightsStore[8][406]<=0;WeightsStore[8][407]<=0;WeightsStore[8][408]<=0;WeightsStore[8][409]<=0;WeightsStore[8][410]<=0;WeightsStore[8][411]<=0;WeightsStore[8][412]<=0;WeightsStore[8][413]<=0;WeightsStore[8][414]<=0;WeightsStore[8][415]<=0;WeightsStore[8][416]<=0;WeightsStore[8][417]<=0;WeightsStore[8][418]<=0;WeightsStore[8][419]<=0;WeightsStore[8][420]<=0;WeightsStore[8][421]<=0;WeightsStore[8][422]<=0;WeightsStore[8][423]<=0;WeightsStore[8][424]<=0;WeightsStore[8][425]<=0;WeightsStore[8][426]<=0;WeightsStore[8][427]<=0;WeightsStore[8][428]<=0;WeightsStore[8][429]<=0;WeightsStore[8][430]<=0;WeightsStore[8][431]<=0;WeightsStore[8][432]<=0;WeightsStore[8][433]<=0;WeightsStore[8][434]<=0;WeightsStore[8][435]<=0;WeightsStore[8][436]<=0;WeightsStore[8][437]<=0;WeightsStore[8][438]<=0;WeightsStore[8][439]<=0;WeightsStore[8][440]<=0;WeightsStore[8][441]<=0;WeightsStore[8][442]<=0;WeightsStore[8][443]<=0;WeightsStore[8][444]<=0;WeightsStore[8][445]<=0;WeightsStore[8][446]<=0;WeightsStore[8][447]<=0;WeightsStore[8][448]<=0;WeightsStore[8][449]<=0;WeightsStore[8][450]<=0;WeightsStore[8][451]<=0;WeightsStore[8][452]<=0;WeightsStore[8][453]<=0;WeightsStore[8][454]<=0;WeightsStore[8][455]<=0;WeightsStore[8][456]<=0;WeightsStore[8][457]<=0;WeightsStore[8][458]<=0;WeightsStore[8][459]<=0;WeightsStore[8][460]<=0;WeightsStore[8][461]<=0;WeightsStore[8][462]<=0;WeightsStore[8][463]<=0;WeightsStore[8][464]<=0;WeightsStore[8][465]<=0;WeightsStore[8][466]<=0;WeightsStore[8][467]<=0;WeightsStore[8][468]<=0;WeightsStore[8][469]<=0;WeightsStore[8][470]<=0;WeightsStore[8][471]<=0;WeightsStore[8][472]<=0;WeightsStore[8][473]<=0;WeightsStore[8][474]<=0;WeightsStore[8][475]<=0;WeightsStore[8][476]<=0;WeightsStore[8][477]<=0;WeightsStore[8][478]<=0;WeightsStore[8][479]<=0;WeightsStore[8][480]<=0;WeightsStore[8][481]<=0;WeightsStore[8][482]<=0;WeightsStore[8][483]<=0;WeightsStore[8][484]<=0;WeightsStore[8][485]<=0;WeightsStore[8][486]<=0;WeightsStore[8][487]<=0;WeightsStore[8][488]<=0;WeightsStore[8][489]<=0;WeightsStore[8][490]<=0;WeightsStore[8][491]<=0;WeightsStore[8][492]<=0;WeightsStore[8][493]<=0;WeightsStore[8][494]<=0;WeightsStore[8][495]<=0;WeightsStore[8][496]<=0;WeightsStore[8][497]<=0;WeightsStore[8][498]<=0;WeightsStore[8][499]<=0;WeightsStore[8][500]<=0;WeightsStore[8][501]<=0;WeightsStore[8][502]<=0;WeightsStore[8][503]<=0;WeightsStore[8][504]<=0;WeightsStore[8][505]<=0;WeightsStore[8][506]<=0;WeightsStore[8][507]<=0;WeightsStore[8][508]<=0;WeightsStore[8][509]<=0;WeightsStore[8][510]<=0;WeightsStore[8][511]<=0;WeightsStore[8][512]<=0;WeightsStore[8][513]<=0;WeightsStore[8][514]<=0;WeightsStore[8][515]<=0;WeightsStore[8][516]<=0;WeightsStore[8][517]<=0;WeightsStore[8][518]<=0;WeightsStore[8][519]<=0;WeightsStore[8][520]<=0;WeightsStore[8][521]<=0;WeightsStore[8][522]<=0;WeightsStore[8][523]<=0;WeightsStore[8][524]<=0;WeightsStore[8][525]<=0;WeightsStore[8][526]<=0;WeightsStore[8][527]<=0;WeightsStore[8][528]<=0;WeightsStore[8][529]<=0;WeightsStore[8][530]<=0;WeightsStore[8][531]<=0;WeightsStore[8][532]<=0;WeightsStore[8][533]<=0;WeightsStore[8][534]<=0;WeightsStore[8][535]<=0;WeightsStore[8][536]<=0;WeightsStore[8][537]<=0;WeightsStore[8][538]<=0;WeightsStore[8][539]<=0;WeightsStore[8][540]<=0;WeightsStore[8][541]<=0;WeightsStore[8][542]<=0;WeightsStore[8][543]<=0;WeightsStore[8][544]<=0;WeightsStore[8][545]<=0;WeightsStore[8][546]<=0;WeightsStore[8][547]<=0;WeightsStore[8][548]<=0;WeightsStore[8][549]<=0;WeightsStore[8][550]<=0;WeightsStore[8][551]<=0;WeightsStore[8][552]<=0;WeightsStore[8][553]<=0;WeightsStore[8][554]<=0;WeightsStore[8][555]<=0;WeightsStore[8][556]<=0;WeightsStore[8][557]<=0;WeightsStore[8][558]<=0;WeightsStore[8][559]<=0;WeightsStore[8][560]<=0;WeightsStore[8][561]<=0;WeightsStore[8][562]<=0;WeightsStore[8][563]<=0;WeightsStore[8][564]<=0;WeightsStore[8][565]<=0;WeightsStore[8][566]<=0;WeightsStore[8][567]<=0;WeightsStore[8][568]<=0;WeightsStore[8][569]<=0;WeightsStore[8][570]<=0;WeightsStore[8][571]<=0;WeightsStore[8][572]<=0;WeightsStore[8][573]<=0;WeightsStore[8][574]<=0;WeightsStore[8][575]<=0;WeightsStore[8][576]<=0;WeightsStore[8][577]<=0;WeightsStore[8][578]<=0;WeightsStore[8][579]<=0;WeightsStore[8][580]<=0;WeightsStore[8][581]<=0;WeightsStore[8][582]<=0;WeightsStore[8][583]<=0;WeightsStore[8][584]<=0;WeightsStore[8][585]<=0;WeightsStore[8][586]<=0;WeightsStore[8][587]<=0;WeightsStore[8][588]<=0;WeightsStore[8][589]<=0;WeightsStore[8][590]<=0;WeightsStore[8][591]<=0;WeightsStore[8][592]<=0;WeightsStore[8][593]<=0;WeightsStore[8][594]<=0;WeightsStore[8][595]<=0;WeightsStore[8][596]<=0;WeightsStore[8][597]<=0;WeightsStore[8][598]<=0;WeightsStore[8][599]<=0;WeightsStore[8][600]<=0;WeightsStore[8][601]<=0;WeightsStore[8][602]<=0;WeightsStore[8][603]<=0;WeightsStore[8][604]<=0;WeightsStore[8][605]<=0;WeightsStore[8][606]<=0;WeightsStore[8][607]<=0;WeightsStore[8][608]<=0;WeightsStore[8][609]<=0;WeightsStore[8][610]<=0;WeightsStore[8][611]<=0;WeightsStore[8][612]<=0;WeightsStore[8][613]<=0;WeightsStore[8][614]<=0;WeightsStore[8][615]<=0;WeightsStore[8][616]<=0;WeightsStore[8][617]<=0;WeightsStore[8][618]<=0;WeightsStore[8][619]<=0;WeightsStore[8][620]<=0;WeightsStore[8][621]<=0;WeightsStore[8][622]<=0;WeightsStore[8][623]<=0;WeightsStore[8][624]<=0;WeightsStore[8][625]<=0;WeightsStore[8][626]<=0;WeightsStore[8][627]<=0;WeightsStore[8][628]<=0;WeightsStore[8][629]<=0;WeightsStore[8][630]<=0;WeightsStore[8][631]<=0;WeightsStore[8][632]<=0;WeightsStore[8][633]<=0;WeightsStore[8][634]<=0;WeightsStore[8][635]<=0;WeightsStore[8][636]<=0;WeightsStore[8][637]<=0;WeightsStore[8][638]<=0;WeightsStore[8][639]<=0;WeightsStore[8][640]<=0;WeightsStore[8][641]<=0;WeightsStore[8][642]<=0;WeightsStore[8][643]<=0;WeightsStore[8][644]<=0;WeightsStore[8][645]<=0;WeightsStore[8][646]<=0;WeightsStore[8][647]<=0;WeightsStore[8][648]<=0;WeightsStore[8][649]<=0;WeightsStore[8][650]<=0;WeightsStore[8][651]<=0;WeightsStore[8][652]<=0;WeightsStore[8][653]<=0;WeightsStore[8][654]<=0;WeightsStore[8][655]<=0;WeightsStore[8][656]<=0;WeightsStore[8][657]<=0;WeightsStore[8][658]<=0;WeightsStore[8][659]<=0;WeightsStore[8][660]<=0;WeightsStore[8][661]<=0;WeightsStore[8][662]<=0;WeightsStore[8][663]<=0;WeightsStore[8][664]<=0;WeightsStore[8][665]<=0;WeightsStore[8][666]<=0;WeightsStore[8][667]<=0;WeightsStore[8][668]<=0;WeightsStore[8][669]<=0;WeightsStore[8][670]<=0;WeightsStore[8][671]<=0;WeightsStore[8][672]<=0;WeightsStore[8][673]<=0;WeightsStore[8][674]<=0;WeightsStore[8][675]<=0;WeightsStore[8][676]<=0;WeightsStore[8][677]<=0;WeightsStore[8][678]<=0;WeightsStore[8][679]<=0;WeightsStore[8][680]<=0;WeightsStore[8][681]<=0;WeightsStore[8][682]<=0;WeightsStore[8][683]<=0;WeightsStore[8][684]<=0;WeightsStore[8][685]<=0;WeightsStore[8][686]<=0;WeightsStore[8][687]<=0;WeightsStore[8][688]<=0;WeightsStore[8][689]<=0;WeightsStore[8][690]<=0;WeightsStore[8][691]<=0;WeightsStore[8][692]<=0;WeightsStore[8][693]<=0;WeightsStore[8][694]<=0;WeightsStore[8][695]<=0;WeightsStore[8][696]<=0;WeightsStore[8][697]<=0;WeightsStore[8][698]<=0;WeightsStore[8][699]<=0;WeightsStore[8][700]<=0;WeightsStore[8][701]<=0;WeightsStore[8][702]<=0;WeightsStore[8][703]<=0;WeightsStore[8][704]<=0;WeightsStore[8][705]<=0;WeightsStore[8][706]<=0;WeightsStore[8][707]<=0;WeightsStore[8][708]<=0;WeightsStore[8][709]<=0;WeightsStore[8][710]<=0;WeightsStore[8][711]<=0;WeightsStore[8][712]<=0;WeightsStore[8][713]<=0;WeightsStore[8][714]<=0;WeightsStore[8][715]<=0;WeightsStore[8][716]<=0;WeightsStore[8][717]<=0;WeightsStore[8][718]<=0;WeightsStore[8][719]<=0;WeightsStore[8][720]<=0;WeightsStore[8][721]<=0;WeightsStore[8][722]<=0;WeightsStore[8][723]<=0;WeightsStore[8][724]<=0;WeightsStore[8][725]<=0;WeightsStore[8][726]<=0;WeightsStore[8][727]<=0;WeightsStore[8][728]<=0;WeightsStore[8][729]<=0;WeightsStore[8][730]<=0;WeightsStore[8][731]<=0;WeightsStore[8][732]<=0;WeightsStore[8][733]<=0;WeightsStore[8][734]<=0;WeightsStore[8][735]<=0;WeightsStore[8][736]<=0;WeightsStore[8][737]<=0;WeightsStore[8][738]<=0;WeightsStore[8][739]<=0;WeightsStore[8][740]<=0;WeightsStore[8][741]<=0;WeightsStore[8][742]<=0;WeightsStore[8][743]<=0;WeightsStore[8][744]<=0;WeightsStore[8][745]<=0;WeightsStore[8][746]<=0;WeightsStore[8][747]<=0;WeightsStore[8][748]<=0;WeightsStore[8][749]<=0;WeightsStore[8][750]<=0;WeightsStore[8][751]<=0;WeightsStore[8][752]<=0;WeightsStore[8][753]<=0;WeightsStore[8][754]<=0;WeightsStore[8][755]<=0;WeightsStore[8][756]<=0;WeightsStore[8][757]<=0;WeightsStore[8][758]<=0;WeightsStore[8][759]<=0;WeightsStore[8][760]<=0;WeightsStore[8][761]<=0;WeightsStore[8][762]<=0;WeightsStore[8][763]<=0;WeightsStore[8][764]<=0;WeightsStore[8][765]<=0;WeightsStore[8][766]<=0;WeightsStore[8][767]<=0;WeightsStore[8][768]<=0;WeightsStore[8][769]<=0;WeightsStore[8][770]<=0;WeightsStore[8][771]<=0;WeightsStore[8][772]<=0;WeightsStore[8][773]<=0;WeightsStore[8][774]<=0;WeightsStore[8][775]<=0;WeightsStore[8][776]<=0;WeightsStore[8][777]<=0;WeightsStore[8][778]<=0;WeightsStore[8][779]<=0;WeightsStore[8][780]<=0;WeightsStore[8][781]<=0;WeightsStore[8][782]<=0;WeightsStore[8][783]<=0;WeightsStore[8][784]<=0;WeightsStore[9][0]<=0;WeightsStore[9][1]<=0;WeightsStore[9][2]<=0;WeightsStore[9][3]<=0;WeightsStore[9][4]<=0;WeightsStore[9][5]<=0;WeightsStore[9][6]<=0;WeightsStore[9][7]<=0;WeightsStore[9][8]<=0;WeightsStore[9][9]<=0;WeightsStore[9][10]<=0;WeightsStore[9][11]<=0;WeightsStore[9][12]<=0;WeightsStore[9][13]<=0;WeightsStore[9][14]<=0;WeightsStore[9][15]<=0;WeightsStore[9][16]<=0;WeightsStore[9][17]<=0;WeightsStore[9][18]<=0;WeightsStore[9][19]<=0;WeightsStore[9][20]<=0;WeightsStore[9][21]<=0;WeightsStore[9][22]<=0;WeightsStore[9][23]<=0;WeightsStore[9][24]<=0;WeightsStore[9][25]<=0;WeightsStore[9][26]<=0;WeightsStore[9][27]<=0;WeightsStore[9][28]<=0;WeightsStore[9][29]<=0;WeightsStore[9][30]<=0;WeightsStore[9][31]<=0;WeightsStore[9][32]<=0;WeightsStore[9][33]<=0;WeightsStore[9][34]<=0;WeightsStore[9][35]<=0;WeightsStore[9][36]<=0;WeightsStore[9][37]<=0;WeightsStore[9][38]<=0;WeightsStore[9][39]<=0;WeightsStore[9][40]<=0;WeightsStore[9][41]<=0;WeightsStore[9][42]<=0;WeightsStore[9][43]<=0;WeightsStore[9][44]<=0;WeightsStore[9][45]<=0;WeightsStore[9][46]<=0;WeightsStore[9][47]<=0;WeightsStore[9][48]<=0;WeightsStore[9][49]<=0;WeightsStore[9][50]<=0;WeightsStore[9][51]<=0;WeightsStore[9][52]<=0;WeightsStore[9][53]<=0;WeightsStore[9][54]<=0;WeightsStore[9][55]<=0;WeightsStore[9][56]<=0;WeightsStore[9][57]<=0;WeightsStore[9][58]<=0;WeightsStore[9][59]<=0;WeightsStore[9][60]<=0;WeightsStore[9][61]<=0;WeightsStore[9][62]<=0;WeightsStore[9][63]<=0;WeightsStore[9][64]<=0;WeightsStore[9][65]<=0;WeightsStore[9][66]<=0;WeightsStore[9][67]<=0;WeightsStore[9][68]<=0;WeightsStore[9][69]<=0;WeightsStore[9][70]<=0;WeightsStore[9][71]<=0;WeightsStore[9][72]<=0;WeightsStore[9][73]<=0;WeightsStore[9][74]<=0;WeightsStore[9][75]<=0;WeightsStore[9][76]<=0;WeightsStore[9][77]<=0;WeightsStore[9][78]<=0;WeightsStore[9][79]<=0;WeightsStore[9][80]<=0;WeightsStore[9][81]<=0;WeightsStore[9][82]<=0;WeightsStore[9][83]<=0;WeightsStore[9][84]<=0;WeightsStore[9][85]<=0;WeightsStore[9][86]<=0;WeightsStore[9][87]<=0;WeightsStore[9][88]<=0;WeightsStore[9][89]<=0;WeightsStore[9][90]<=0;WeightsStore[9][91]<=0;WeightsStore[9][92]<=0;WeightsStore[9][93]<=0;WeightsStore[9][94]<=0;WeightsStore[9][95]<=0;WeightsStore[9][96]<=0;WeightsStore[9][97]<=0;WeightsStore[9][98]<=0;WeightsStore[9][99]<=0;WeightsStore[9][100]<=0;WeightsStore[9][101]<=0;WeightsStore[9][102]<=0;WeightsStore[9][103]<=0;WeightsStore[9][104]<=0;WeightsStore[9][105]<=0;WeightsStore[9][106]<=0;WeightsStore[9][107]<=0;WeightsStore[9][108]<=0;WeightsStore[9][109]<=0;WeightsStore[9][110]<=0;WeightsStore[9][111]<=0;WeightsStore[9][112]<=0;WeightsStore[9][113]<=0;WeightsStore[9][114]<=0;WeightsStore[9][115]<=0;WeightsStore[9][116]<=0;WeightsStore[9][117]<=0;WeightsStore[9][118]<=0;WeightsStore[9][119]<=0;WeightsStore[9][120]<=0;WeightsStore[9][121]<=0;WeightsStore[9][122]<=0;WeightsStore[9][123]<=0;WeightsStore[9][124]<=0;WeightsStore[9][125]<=0;WeightsStore[9][126]<=0;WeightsStore[9][127]<=0;WeightsStore[9][128]<=0;WeightsStore[9][129]<=0;WeightsStore[9][130]<=0;WeightsStore[9][131]<=0;WeightsStore[9][132]<=0;WeightsStore[9][133]<=0;WeightsStore[9][134]<=0;WeightsStore[9][135]<=0;WeightsStore[9][136]<=0;WeightsStore[9][137]<=0;WeightsStore[9][138]<=0;WeightsStore[9][139]<=0;WeightsStore[9][140]<=0;WeightsStore[9][141]<=0;WeightsStore[9][142]<=0;WeightsStore[9][143]<=0;WeightsStore[9][144]<=0;WeightsStore[9][145]<=0;WeightsStore[9][146]<=0;WeightsStore[9][147]<=0;WeightsStore[9][148]<=0;WeightsStore[9][149]<=0;WeightsStore[9][150]<=0;WeightsStore[9][151]<=0;WeightsStore[9][152]<=0;WeightsStore[9][153]<=0;WeightsStore[9][154]<=0;WeightsStore[9][155]<=0;WeightsStore[9][156]<=0;WeightsStore[9][157]<=0;WeightsStore[9][158]<=0;WeightsStore[9][159]<=0;WeightsStore[9][160]<=0;WeightsStore[9][161]<=0;WeightsStore[9][162]<=0;WeightsStore[9][163]<=0;WeightsStore[9][164]<=0;WeightsStore[9][165]<=0;WeightsStore[9][166]<=0;WeightsStore[9][167]<=0;WeightsStore[9][168]<=0;WeightsStore[9][169]<=0;WeightsStore[9][170]<=0;WeightsStore[9][171]<=0;WeightsStore[9][172]<=0;WeightsStore[9][173]<=0;WeightsStore[9][174]<=0;WeightsStore[9][175]<=0;WeightsStore[9][176]<=0;WeightsStore[9][177]<=0;WeightsStore[9][178]<=0;WeightsStore[9][179]<=0;WeightsStore[9][180]<=0;WeightsStore[9][181]<=0;WeightsStore[9][182]<=0;WeightsStore[9][183]<=0;WeightsStore[9][184]<=0;WeightsStore[9][185]<=0;WeightsStore[9][186]<=0;WeightsStore[9][187]<=0;WeightsStore[9][188]<=0;WeightsStore[9][189]<=0;WeightsStore[9][190]<=0;WeightsStore[9][191]<=0;WeightsStore[9][192]<=0;WeightsStore[9][193]<=0;WeightsStore[9][194]<=0;WeightsStore[9][195]<=0;WeightsStore[9][196]<=0;WeightsStore[9][197]<=0;WeightsStore[9][198]<=0;WeightsStore[9][199]<=0;WeightsStore[9][200]<=0;WeightsStore[9][201]<=0;WeightsStore[9][202]<=0;WeightsStore[9][203]<=0;WeightsStore[9][204]<=0;WeightsStore[9][205]<=0;WeightsStore[9][206]<=0;WeightsStore[9][207]<=0;WeightsStore[9][208]<=0;WeightsStore[9][209]<=0;WeightsStore[9][210]<=0;WeightsStore[9][211]<=0;WeightsStore[9][212]<=0;WeightsStore[9][213]<=0;WeightsStore[9][214]<=0;WeightsStore[9][215]<=0;WeightsStore[9][216]<=0;WeightsStore[9][217]<=0;WeightsStore[9][218]<=0;WeightsStore[9][219]<=0;WeightsStore[9][220]<=0;WeightsStore[9][221]<=0;WeightsStore[9][222]<=0;WeightsStore[9][223]<=0;WeightsStore[9][224]<=0;WeightsStore[9][225]<=0;WeightsStore[9][226]<=0;WeightsStore[9][227]<=0;WeightsStore[9][228]<=0;WeightsStore[9][229]<=0;WeightsStore[9][230]<=0;WeightsStore[9][231]<=0;WeightsStore[9][232]<=0;WeightsStore[9][233]<=0;WeightsStore[9][234]<=0;WeightsStore[9][235]<=0;WeightsStore[9][236]<=0;WeightsStore[9][237]<=0;WeightsStore[9][238]<=0;WeightsStore[9][239]<=0;WeightsStore[9][240]<=0;WeightsStore[9][241]<=0;WeightsStore[9][242]<=0;WeightsStore[9][243]<=0;WeightsStore[9][244]<=0;WeightsStore[9][245]<=0;WeightsStore[9][246]<=0;WeightsStore[9][247]<=0;WeightsStore[9][248]<=0;WeightsStore[9][249]<=0;WeightsStore[9][250]<=0;WeightsStore[9][251]<=0;WeightsStore[9][252]<=0;WeightsStore[9][253]<=0;WeightsStore[9][254]<=0;WeightsStore[9][255]<=0;WeightsStore[9][256]<=0;WeightsStore[9][257]<=0;WeightsStore[9][258]<=0;WeightsStore[9][259]<=0;WeightsStore[9][260]<=0;WeightsStore[9][261]<=0;WeightsStore[9][262]<=0;WeightsStore[9][263]<=0;WeightsStore[9][264]<=0;WeightsStore[9][265]<=0;WeightsStore[9][266]<=0;WeightsStore[9][267]<=0;WeightsStore[9][268]<=0;WeightsStore[9][269]<=0;WeightsStore[9][270]<=0;WeightsStore[9][271]<=0;WeightsStore[9][272]<=0;WeightsStore[9][273]<=0;WeightsStore[9][274]<=0;WeightsStore[9][275]<=0;WeightsStore[9][276]<=0;WeightsStore[9][277]<=0;WeightsStore[9][278]<=0;WeightsStore[9][279]<=0;WeightsStore[9][280]<=0;WeightsStore[9][281]<=0;WeightsStore[9][282]<=0;WeightsStore[9][283]<=0;WeightsStore[9][284]<=0;WeightsStore[9][285]<=0;WeightsStore[9][286]<=0;WeightsStore[9][287]<=0;WeightsStore[9][288]<=0;WeightsStore[9][289]<=0;WeightsStore[9][290]<=0;WeightsStore[9][291]<=0;WeightsStore[9][292]<=0;WeightsStore[9][293]<=0;WeightsStore[9][294]<=0;WeightsStore[9][295]<=0;WeightsStore[9][296]<=0;WeightsStore[9][297]<=0;WeightsStore[9][298]<=0;WeightsStore[9][299]<=0;WeightsStore[9][300]<=0;WeightsStore[9][301]<=0;WeightsStore[9][302]<=0;WeightsStore[9][303]<=0;WeightsStore[9][304]<=0;WeightsStore[9][305]<=0;WeightsStore[9][306]<=0;WeightsStore[9][307]<=0;WeightsStore[9][308]<=0;WeightsStore[9][309]<=0;WeightsStore[9][310]<=0;WeightsStore[9][311]<=0;WeightsStore[9][312]<=0;WeightsStore[9][313]<=0;WeightsStore[9][314]<=0;WeightsStore[9][315]<=0;WeightsStore[9][316]<=0;WeightsStore[9][317]<=0;WeightsStore[9][318]<=0;WeightsStore[9][319]<=0;WeightsStore[9][320]<=0;WeightsStore[9][321]<=0;WeightsStore[9][322]<=0;WeightsStore[9][323]<=0;WeightsStore[9][324]<=0;WeightsStore[9][325]<=0;WeightsStore[9][326]<=0;WeightsStore[9][327]<=0;WeightsStore[9][328]<=0;WeightsStore[9][329]<=0;WeightsStore[9][330]<=0;WeightsStore[9][331]<=0;WeightsStore[9][332]<=0;WeightsStore[9][333]<=0;WeightsStore[9][334]<=0;WeightsStore[9][335]<=0;WeightsStore[9][336]<=0;WeightsStore[9][337]<=0;WeightsStore[9][338]<=0;WeightsStore[9][339]<=0;WeightsStore[9][340]<=0;WeightsStore[9][341]<=0;WeightsStore[9][342]<=0;WeightsStore[9][343]<=0;WeightsStore[9][344]<=0;WeightsStore[9][345]<=0;WeightsStore[9][346]<=0;WeightsStore[9][347]<=0;WeightsStore[9][348]<=0;WeightsStore[9][349]<=0;WeightsStore[9][350]<=0;WeightsStore[9][351]<=0;WeightsStore[9][352]<=0;WeightsStore[9][353]<=0;WeightsStore[9][354]<=0;WeightsStore[9][355]<=0;WeightsStore[9][356]<=0;WeightsStore[9][357]<=0;WeightsStore[9][358]<=0;WeightsStore[9][359]<=0;WeightsStore[9][360]<=0;WeightsStore[9][361]<=0;WeightsStore[9][362]<=0;WeightsStore[9][363]<=0;WeightsStore[9][364]<=0;WeightsStore[9][365]<=0;WeightsStore[9][366]<=0;WeightsStore[9][367]<=0;WeightsStore[9][368]<=0;WeightsStore[9][369]<=0;WeightsStore[9][370]<=0;WeightsStore[9][371]<=0;WeightsStore[9][372]<=0;WeightsStore[9][373]<=0;WeightsStore[9][374]<=0;WeightsStore[9][375]<=0;WeightsStore[9][376]<=0;WeightsStore[9][377]<=0;WeightsStore[9][378]<=0;WeightsStore[9][379]<=0;WeightsStore[9][380]<=0;WeightsStore[9][381]<=0;WeightsStore[9][382]<=0;WeightsStore[9][383]<=0;WeightsStore[9][384]<=0;WeightsStore[9][385]<=0;WeightsStore[9][386]<=0;WeightsStore[9][387]<=0;WeightsStore[9][388]<=0;WeightsStore[9][389]<=0;WeightsStore[9][390]<=0;WeightsStore[9][391]<=0;WeightsStore[9][392]<=0;WeightsStore[9][393]<=0;WeightsStore[9][394]<=0;WeightsStore[9][395]<=0;WeightsStore[9][396]<=0;WeightsStore[9][397]<=0;WeightsStore[9][398]<=0;WeightsStore[9][399]<=0;WeightsStore[9][400]<=0;WeightsStore[9][401]<=0;WeightsStore[9][402]<=0;WeightsStore[9][403]<=0;WeightsStore[9][404]<=0;WeightsStore[9][405]<=0;WeightsStore[9][406]<=0;WeightsStore[9][407]<=0;WeightsStore[9][408]<=0;WeightsStore[9][409]<=0;WeightsStore[9][410]<=0;WeightsStore[9][411]<=0;WeightsStore[9][412]<=0;WeightsStore[9][413]<=0;WeightsStore[9][414]<=0;WeightsStore[9][415]<=0;WeightsStore[9][416]<=0;WeightsStore[9][417]<=0;WeightsStore[9][418]<=0;WeightsStore[9][419]<=0;WeightsStore[9][420]<=0;WeightsStore[9][421]<=0;WeightsStore[9][422]<=0;WeightsStore[9][423]<=0;WeightsStore[9][424]<=0;WeightsStore[9][425]<=0;WeightsStore[9][426]<=0;WeightsStore[9][427]<=0;WeightsStore[9][428]<=0;WeightsStore[9][429]<=0;WeightsStore[9][430]<=0;WeightsStore[9][431]<=0;WeightsStore[9][432]<=0;WeightsStore[9][433]<=0;WeightsStore[9][434]<=0;WeightsStore[9][435]<=0;WeightsStore[9][436]<=0;WeightsStore[9][437]<=0;WeightsStore[9][438]<=0;WeightsStore[9][439]<=0;WeightsStore[9][440]<=0;WeightsStore[9][441]<=0;WeightsStore[9][442]<=0;WeightsStore[9][443]<=0;WeightsStore[9][444]<=0;WeightsStore[9][445]<=0;WeightsStore[9][446]<=0;WeightsStore[9][447]<=0;WeightsStore[9][448]<=0;WeightsStore[9][449]<=0;WeightsStore[9][450]<=0;WeightsStore[9][451]<=0;WeightsStore[9][452]<=0;WeightsStore[9][453]<=0;WeightsStore[9][454]<=0;WeightsStore[9][455]<=0;WeightsStore[9][456]<=0;WeightsStore[9][457]<=0;WeightsStore[9][458]<=0;WeightsStore[9][459]<=0;WeightsStore[9][460]<=0;WeightsStore[9][461]<=0;WeightsStore[9][462]<=0;WeightsStore[9][463]<=0;WeightsStore[9][464]<=0;WeightsStore[9][465]<=0;WeightsStore[9][466]<=0;WeightsStore[9][467]<=0;WeightsStore[9][468]<=0;WeightsStore[9][469]<=0;WeightsStore[9][470]<=0;WeightsStore[9][471]<=0;WeightsStore[9][472]<=0;WeightsStore[9][473]<=0;WeightsStore[9][474]<=0;WeightsStore[9][475]<=0;WeightsStore[9][476]<=0;WeightsStore[9][477]<=0;WeightsStore[9][478]<=0;WeightsStore[9][479]<=0;WeightsStore[9][480]<=0;WeightsStore[9][481]<=0;WeightsStore[9][482]<=0;WeightsStore[9][483]<=0;WeightsStore[9][484]<=0;WeightsStore[9][485]<=0;WeightsStore[9][486]<=0;WeightsStore[9][487]<=0;WeightsStore[9][488]<=0;WeightsStore[9][489]<=0;WeightsStore[9][490]<=0;WeightsStore[9][491]<=0;WeightsStore[9][492]<=0;WeightsStore[9][493]<=0;WeightsStore[9][494]<=0;WeightsStore[9][495]<=0;WeightsStore[9][496]<=0;WeightsStore[9][497]<=0;WeightsStore[9][498]<=0;WeightsStore[9][499]<=0;WeightsStore[9][500]<=0;WeightsStore[9][501]<=0;WeightsStore[9][502]<=0;WeightsStore[9][503]<=0;WeightsStore[9][504]<=0;WeightsStore[9][505]<=0;WeightsStore[9][506]<=0;WeightsStore[9][507]<=0;WeightsStore[9][508]<=0;WeightsStore[9][509]<=0;WeightsStore[9][510]<=0;WeightsStore[9][511]<=0;WeightsStore[9][512]<=0;WeightsStore[9][513]<=0;WeightsStore[9][514]<=0;WeightsStore[9][515]<=0;WeightsStore[9][516]<=0;WeightsStore[9][517]<=0;WeightsStore[9][518]<=0;WeightsStore[9][519]<=0;WeightsStore[9][520]<=0;WeightsStore[9][521]<=0;WeightsStore[9][522]<=0;WeightsStore[9][523]<=0;WeightsStore[9][524]<=0;WeightsStore[9][525]<=0;WeightsStore[9][526]<=0;WeightsStore[9][527]<=0;WeightsStore[9][528]<=0;WeightsStore[9][529]<=0;WeightsStore[9][530]<=0;WeightsStore[9][531]<=0;WeightsStore[9][532]<=0;WeightsStore[9][533]<=0;WeightsStore[9][534]<=0;WeightsStore[9][535]<=0;WeightsStore[9][536]<=0;WeightsStore[9][537]<=0;WeightsStore[9][538]<=0;WeightsStore[9][539]<=0;WeightsStore[9][540]<=0;WeightsStore[9][541]<=0;WeightsStore[9][542]<=0;WeightsStore[9][543]<=0;WeightsStore[9][544]<=0;WeightsStore[9][545]<=0;WeightsStore[9][546]<=0;WeightsStore[9][547]<=0;WeightsStore[9][548]<=0;WeightsStore[9][549]<=0;WeightsStore[9][550]<=0;WeightsStore[9][551]<=0;WeightsStore[9][552]<=0;WeightsStore[9][553]<=0;WeightsStore[9][554]<=0;WeightsStore[9][555]<=0;WeightsStore[9][556]<=0;WeightsStore[9][557]<=0;WeightsStore[9][558]<=0;WeightsStore[9][559]<=0;WeightsStore[9][560]<=0;WeightsStore[9][561]<=0;WeightsStore[9][562]<=0;WeightsStore[9][563]<=0;WeightsStore[9][564]<=0;WeightsStore[9][565]<=0;WeightsStore[9][566]<=0;WeightsStore[9][567]<=0;WeightsStore[9][568]<=0;WeightsStore[9][569]<=0;WeightsStore[9][570]<=0;WeightsStore[9][571]<=0;WeightsStore[9][572]<=0;WeightsStore[9][573]<=0;WeightsStore[9][574]<=0;WeightsStore[9][575]<=0;WeightsStore[9][576]<=0;WeightsStore[9][577]<=0;WeightsStore[9][578]<=0;WeightsStore[9][579]<=0;WeightsStore[9][580]<=0;WeightsStore[9][581]<=0;WeightsStore[9][582]<=0;WeightsStore[9][583]<=0;WeightsStore[9][584]<=0;WeightsStore[9][585]<=0;WeightsStore[9][586]<=0;WeightsStore[9][587]<=0;WeightsStore[9][588]<=0;WeightsStore[9][589]<=0;WeightsStore[9][590]<=0;WeightsStore[9][591]<=0;WeightsStore[9][592]<=0;WeightsStore[9][593]<=0;WeightsStore[9][594]<=0;WeightsStore[9][595]<=0;WeightsStore[9][596]<=0;WeightsStore[9][597]<=0;WeightsStore[9][598]<=0;WeightsStore[9][599]<=0;WeightsStore[9][600]<=0;WeightsStore[9][601]<=0;WeightsStore[9][602]<=0;WeightsStore[9][603]<=0;WeightsStore[9][604]<=0;WeightsStore[9][605]<=0;WeightsStore[9][606]<=0;WeightsStore[9][607]<=0;WeightsStore[9][608]<=0;WeightsStore[9][609]<=0;WeightsStore[9][610]<=0;WeightsStore[9][611]<=0;WeightsStore[9][612]<=0;WeightsStore[9][613]<=0;WeightsStore[9][614]<=0;WeightsStore[9][615]<=0;WeightsStore[9][616]<=0;WeightsStore[9][617]<=0;WeightsStore[9][618]<=0;WeightsStore[9][619]<=0;WeightsStore[9][620]<=0;WeightsStore[9][621]<=0;WeightsStore[9][622]<=0;WeightsStore[9][623]<=0;WeightsStore[9][624]<=0;WeightsStore[9][625]<=0;WeightsStore[9][626]<=0;WeightsStore[9][627]<=0;WeightsStore[9][628]<=0;WeightsStore[9][629]<=0;WeightsStore[9][630]<=0;WeightsStore[9][631]<=0;WeightsStore[9][632]<=0;WeightsStore[9][633]<=0;WeightsStore[9][634]<=0;WeightsStore[9][635]<=0;WeightsStore[9][636]<=0;WeightsStore[9][637]<=0;WeightsStore[9][638]<=0;WeightsStore[9][639]<=0;WeightsStore[9][640]<=0;WeightsStore[9][641]<=0;WeightsStore[9][642]<=0;WeightsStore[9][643]<=0;WeightsStore[9][644]<=0;WeightsStore[9][645]<=0;WeightsStore[9][646]<=0;WeightsStore[9][647]<=0;WeightsStore[9][648]<=0;WeightsStore[9][649]<=0;WeightsStore[9][650]<=0;WeightsStore[9][651]<=0;WeightsStore[9][652]<=0;WeightsStore[9][653]<=0;WeightsStore[9][654]<=0;WeightsStore[9][655]<=0;WeightsStore[9][656]<=0;WeightsStore[9][657]<=0;WeightsStore[9][658]<=0;WeightsStore[9][659]<=0;WeightsStore[9][660]<=0;WeightsStore[9][661]<=0;WeightsStore[9][662]<=0;WeightsStore[9][663]<=0;WeightsStore[9][664]<=0;WeightsStore[9][665]<=0;WeightsStore[9][666]<=0;WeightsStore[9][667]<=0;WeightsStore[9][668]<=0;WeightsStore[9][669]<=0;WeightsStore[9][670]<=0;WeightsStore[9][671]<=0;WeightsStore[9][672]<=0;WeightsStore[9][673]<=0;WeightsStore[9][674]<=0;WeightsStore[9][675]<=0;WeightsStore[9][676]<=0;WeightsStore[9][677]<=0;WeightsStore[9][678]<=0;WeightsStore[9][679]<=0;WeightsStore[9][680]<=0;WeightsStore[9][681]<=0;WeightsStore[9][682]<=0;WeightsStore[9][683]<=0;WeightsStore[9][684]<=0;WeightsStore[9][685]<=0;WeightsStore[9][686]<=0;WeightsStore[9][687]<=0;WeightsStore[9][688]<=0;WeightsStore[9][689]<=0;WeightsStore[9][690]<=0;WeightsStore[9][691]<=0;WeightsStore[9][692]<=0;WeightsStore[9][693]<=0;WeightsStore[9][694]<=0;WeightsStore[9][695]<=0;WeightsStore[9][696]<=0;WeightsStore[9][697]<=0;WeightsStore[9][698]<=0;WeightsStore[9][699]<=0;WeightsStore[9][700]<=0;WeightsStore[9][701]<=0;WeightsStore[9][702]<=0;WeightsStore[9][703]<=0;WeightsStore[9][704]<=0;WeightsStore[9][705]<=0;WeightsStore[9][706]<=0;WeightsStore[9][707]<=0;WeightsStore[9][708]<=0;WeightsStore[9][709]<=0;WeightsStore[9][710]<=0;WeightsStore[9][711]<=0;WeightsStore[9][712]<=0;WeightsStore[9][713]<=0;WeightsStore[9][714]<=0;WeightsStore[9][715]<=0;WeightsStore[9][716]<=0;WeightsStore[9][717]<=0;WeightsStore[9][718]<=0;WeightsStore[9][719]<=0;WeightsStore[9][720]<=0;WeightsStore[9][721]<=0;WeightsStore[9][722]<=0;WeightsStore[9][723]<=0;WeightsStore[9][724]<=0;WeightsStore[9][725]<=0;WeightsStore[9][726]<=0;WeightsStore[9][727]<=0;WeightsStore[9][728]<=0;WeightsStore[9][729]<=0;WeightsStore[9][730]<=0;WeightsStore[9][731]<=0;WeightsStore[9][732]<=0;WeightsStore[9][733]<=0;WeightsStore[9][734]<=0;WeightsStore[9][735]<=0;WeightsStore[9][736]<=0;WeightsStore[9][737]<=0;WeightsStore[9][738]<=0;WeightsStore[9][739]<=0;WeightsStore[9][740]<=0;WeightsStore[9][741]<=0;WeightsStore[9][742]<=0;WeightsStore[9][743]<=0;WeightsStore[9][744]<=0;WeightsStore[9][745]<=0;WeightsStore[9][746]<=0;WeightsStore[9][747]<=0;WeightsStore[9][748]<=0;WeightsStore[9][749]<=0;WeightsStore[9][750]<=0;WeightsStore[9][751]<=0;WeightsStore[9][752]<=0;WeightsStore[9][753]<=0;WeightsStore[9][754]<=0;WeightsStore[9][755]<=0;WeightsStore[9][756]<=0;WeightsStore[9][757]<=0;WeightsStore[9][758]<=0;WeightsStore[9][759]<=0;WeightsStore[9][760]<=0;WeightsStore[9][761]<=0;WeightsStore[9][762]<=0;WeightsStore[9][763]<=0;WeightsStore[9][764]<=0;WeightsStore[9][765]<=0;WeightsStore[9][766]<=0;WeightsStore[9][767]<=0;WeightsStore[9][768]<=0;WeightsStore[9][769]<=0;WeightsStore[9][770]<=0;WeightsStore[9][771]<=0;WeightsStore[9][772]<=0;WeightsStore[9][773]<=0;WeightsStore[9][774]<=0;WeightsStore[9][775]<=0;WeightsStore[9][776]<=0;WeightsStore[9][777]<=0;WeightsStore[9][778]<=0;WeightsStore[9][779]<=0;WeightsStore[9][780]<=0;WeightsStore[9][781]<=0;WeightsStore[9][782]<=0;WeightsStore[9][783]<=0;WeightsStore[9][784]<=0;
	end
	if(Input_Valid == 1'b1)begin
		switchCounter <= 32'd0;
		ready = 1'b0;
		internalReset = 1'b0;
		PixelsStore[0]<=Pix_0;PixelsStore[1]<=Pix_1;PixelsStore[2]<=Pix_2;PixelsStore[3]<=Pix_3;PixelsStore[4]<=Pix_4;PixelsStore[5]<=Pix_5;PixelsStore[6]<=Pix_6;PixelsStore[7]<=Pix_7;PixelsStore[8]<=Pix_8;PixelsStore[9]<=Pix_9;PixelsStore[10]<=Pix_10;PixelsStore[11]<=Pix_11;PixelsStore[12]<=Pix_12;PixelsStore[13]<=Pix_13;PixelsStore[14]<=Pix_14;PixelsStore[15]<=Pix_15;PixelsStore[16]<=Pix_16;PixelsStore[17]<=Pix_17;PixelsStore[18]<=Pix_18;PixelsStore[19]<=Pix_19;PixelsStore[20]<=Pix_20;PixelsStore[21]<=Pix_21;PixelsStore[22]<=Pix_22;PixelsStore[23]<=Pix_23;PixelsStore[24]<=Pix_24;PixelsStore[25]<=Pix_25;PixelsStore[26]<=Pix_26;PixelsStore[27]<=Pix_27;PixelsStore[28]<=Pix_28;PixelsStore[29]<=Pix_29;PixelsStore[30]<=Pix_30;PixelsStore[31]<=Pix_31;PixelsStore[32]<=Pix_32;PixelsStore[33]<=Pix_33;PixelsStore[34]<=Pix_34;PixelsStore[35]<=Pix_35;PixelsStore[36]<=Pix_36;PixelsStore[37]<=Pix_37;PixelsStore[38]<=Pix_38;PixelsStore[39]<=Pix_39;PixelsStore[40]<=Pix_40;PixelsStore[41]<=Pix_41;PixelsStore[42]<=Pix_42;PixelsStore[43]<=Pix_43;PixelsStore[44]<=Pix_44;PixelsStore[45]<=Pix_45;PixelsStore[46]<=Pix_46;PixelsStore[47]<=Pix_47;PixelsStore[48]<=Pix_48;PixelsStore[49]<=Pix_49;PixelsStore[50]<=Pix_50;PixelsStore[51]<=Pix_51;PixelsStore[52]<=Pix_52;PixelsStore[53]<=Pix_53;PixelsStore[54]<=Pix_54;PixelsStore[55]<=Pix_55;PixelsStore[56]<=Pix_56;PixelsStore[57]<=Pix_57;PixelsStore[58]<=Pix_58;PixelsStore[59]<=Pix_59;PixelsStore[60]<=Pix_60;PixelsStore[61]<=Pix_61;PixelsStore[62]<=Pix_62;PixelsStore[63]<=Pix_63;PixelsStore[64]<=Pix_64;PixelsStore[65]<=Pix_65;PixelsStore[66]<=Pix_66;PixelsStore[67]<=Pix_67;PixelsStore[68]<=Pix_68;PixelsStore[69]<=Pix_69;PixelsStore[70]<=Pix_70;PixelsStore[71]<=Pix_71;PixelsStore[72]<=Pix_72;PixelsStore[73]<=Pix_73;PixelsStore[74]<=Pix_74;PixelsStore[75]<=Pix_75;PixelsStore[76]<=Pix_76;PixelsStore[77]<=Pix_77;PixelsStore[78]<=Pix_78;PixelsStore[79]<=Pix_79;PixelsStore[80]<=Pix_80;PixelsStore[81]<=Pix_81;PixelsStore[82]<=Pix_82;PixelsStore[83]<=Pix_83;PixelsStore[84]<=Pix_84;PixelsStore[85]<=Pix_85;PixelsStore[86]<=Pix_86;PixelsStore[87]<=Pix_87;PixelsStore[88]<=Pix_88;PixelsStore[89]<=Pix_89;PixelsStore[90]<=Pix_90;PixelsStore[91]<=Pix_91;PixelsStore[92]<=Pix_92;PixelsStore[93]<=Pix_93;PixelsStore[94]<=Pix_94;PixelsStore[95]<=Pix_95;PixelsStore[96]<=Pix_96;PixelsStore[97]<=Pix_97;PixelsStore[98]<=Pix_98;PixelsStore[99]<=Pix_99;PixelsStore[100]<=Pix_100;PixelsStore[101]<=Pix_101;PixelsStore[102]<=Pix_102;PixelsStore[103]<=Pix_103;PixelsStore[104]<=Pix_104;PixelsStore[105]<=Pix_105;PixelsStore[106]<=Pix_106;PixelsStore[107]<=Pix_107;PixelsStore[108]<=Pix_108;PixelsStore[109]<=Pix_109;PixelsStore[110]<=Pix_110;PixelsStore[111]<=Pix_111;PixelsStore[112]<=Pix_112;PixelsStore[113]<=Pix_113;PixelsStore[114]<=Pix_114;PixelsStore[115]<=Pix_115;PixelsStore[116]<=Pix_116;PixelsStore[117]<=Pix_117;PixelsStore[118]<=Pix_118;PixelsStore[119]<=Pix_119;PixelsStore[120]<=Pix_120;PixelsStore[121]<=Pix_121;PixelsStore[122]<=Pix_122;PixelsStore[123]<=Pix_123;PixelsStore[124]<=Pix_124;PixelsStore[125]<=Pix_125;PixelsStore[126]<=Pix_126;PixelsStore[127]<=Pix_127;PixelsStore[128]<=Pix_128;PixelsStore[129]<=Pix_129;PixelsStore[130]<=Pix_130;PixelsStore[131]<=Pix_131;PixelsStore[132]<=Pix_132;PixelsStore[133]<=Pix_133;PixelsStore[134]<=Pix_134;PixelsStore[135]<=Pix_135;PixelsStore[136]<=Pix_136;PixelsStore[137]<=Pix_137;PixelsStore[138]<=Pix_138;PixelsStore[139]<=Pix_139;PixelsStore[140]<=Pix_140;PixelsStore[141]<=Pix_141;PixelsStore[142]<=Pix_142;PixelsStore[143]<=Pix_143;PixelsStore[144]<=Pix_144;PixelsStore[145]<=Pix_145;PixelsStore[146]<=Pix_146;PixelsStore[147]<=Pix_147;PixelsStore[148]<=Pix_148;PixelsStore[149]<=Pix_149;PixelsStore[150]<=Pix_150;PixelsStore[151]<=Pix_151;PixelsStore[152]<=Pix_152;PixelsStore[153]<=Pix_153;PixelsStore[154]<=Pix_154;PixelsStore[155]<=Pix_155;PixelsStore[156]<=Pix_156;PixelsStore[157]<=Pix_157;PixelsStore[158]<=Pix_158;PixelsStore[159]<=Pix_159;PixelsStore[160]<=Pix_160;PixelsStore[161]<=Pix_161;PixelsStore[162]<=Pix_162;PixelsStore[163]<=Pix_163;PixelsStore[164]<=Pix_164;PixelsStore[165]<=Pix_165;PixelsStore[166]<=Pix_166;PixelsStore[167]<=Pix_167;PixelsStore[168]<=Pix_168;PixelsStore[169]<=Pix_169;PixelsStore[170]<=Pix_170;PixelsStore[171]<=Pix_171;PixelsStore[172]<=Pix_172;PixelsStore[173]<=Pix_173;PixelsStore[174]<=Pix_174;PixelsStore[175]<=Pix_175;PixelsStore[176]<=Pix_176;PixelsStore[177]<=Pix_177;PixelsStore[178]<=Pix_178;PixelsStore[179]<=Pix_179;PixelsStore[180]<=Pix_180;PixelsStore[181]<=Pix_181;PixelsStore[182]<=Pix_182;PixelsStore[183]<=Pix_183;PixelsStore[184]<=Pix_184;PixelsStore[185]<=Pix_185;PixelsStore[186]<=Pix_186;PixelsStore[187]<=Pix_187;PixelsStore[188]<=Pix_188;PixelsStore[189]<=Pix_189;PixelsStore[190]<=Pix_190;PixelsStore[191]<=Pix_191;PixelsStore[192]<=Pix_192;PixelsStore[193]<=Pix_193;PixelsStore[194]<=Pix_194;PixelsStore[195]<=Pix_195;PixelsStore[196]<=Pix_196;PixelsStore[197]<=Pix_197;PixelsStore[198]<=Pix_198;PixelsStore[199]<=Pix_199;PixelsStore[200]<=Pix_200;PixelsStore[201]<=Pix_201;PixelsStore[202]<=Pix_202;PixelsStore[203]<=Pix_203;PixelsStore[204]<=Pix_204;PixelsStore[205]<=Pix_205;PixelsStore[206]<=Pix_206;PixelsStore[207]<=Pix_207;PixelsStore[208]<=Pix_208;PixelsStore[209]<=Pix_209;PixelsStore[210]<=Pix_210;PixelsStore[211]<=Pix_211;PixelsStore[212]<=Pix_212;PixelsStore[213]<=Pix_213;PixelsStore[214]<=Pix_214;PixelsStore[215]<=Pix_215;PixelsStore[216]<=Pix_216;PixelsStore[217]<=Pix_217;PixelsStore[218]<=Pix_218;PixelsStore[219]<=Pix_219;PixelsStore[220]<=Pix_220;PixelsStore[221]<=Pix_221;PixelsStore[222]<=Pix_222;PixelsStore[223]<=Pix_223;PixelsStore[224]<=Pix_224;PixelsStore[225]<=Pix_225;PixelsStore[226]<=Pix_226;PixelsStore[227]<=Pix_227;PixelsStore[228]<=Pix_228;PixelsStore[229]<=Pix_229;PixelsStore[230]<=Pix_230;PixelsStore[231]<=Pix_231;PixelsStore[232]<=Pix_232;PixelsStore[233]<=Pix_233;PixelsStore[234]<=Pix_234;PixelsStore[235]<=Pix_235;PixelsStore[236]<=Pix_236;PixelsStore[237]<=Pix_237;PixelsStore[238]<=Pix_238;PixelsStore[239]<=Pix_239;PixelsStore[240]<=Pix_240;PixelsStore[241]<=Pix_241;PixelsStore[242]<=Pix_242;PixelsStore[243]<=Pix_243;PixelsStore[244]<=Pix_244;PixelsStore[245]<=Pix_245;PixelsStore[246]<=Pix_246;PixelsStore[247]<=Pix_247;PixelsStore[248]<=Pix_248;PixelsStore[249]<=Pix_249;PixelsStore[250]<=Pix_250;PixelsStore[251]<=Pix_251;PixelsStore[252]<=Pix_252;PixelsStore[253]<=Pix_253;PixelsStore[254]<=Pix_254;PixelsStore[255]<=Pix_255;PixelsStore[256]<=Pix_256;PixelsStore[257]<=Pix_257;PixelsStore[258]<=Pix_258;PixelsStore[259]<=Pix_259;PixelsStore[260]<=Pix_260;PixelsStore[261]<=Pix_261;PixelsStore[262]<=Pix_262;PixelsStore[263]<=Pix_263;PixelsStore[264]<=Pix_264;PixelsStore[265]<=Pix_265;PixelsStore[266]<=Pix_266;PixelsStore[267]<=Pix_267;PixelsStore[268]<=Pix_268;PixelsStore[269]<=Pix_269;PixelsStore[270]<=Pix_270;PixelsStore[271]<=Pix_271;PixelsStore[272]<=Pix_272;PixelsStore[273]<=Pix_273;PixelsStore[274]<=Pix_274;PixelsStore[275]<=Pix_275;PixelsStore[276]<=Pix_276;PixelsStore[277]<=Pix_277;PixelsStore[278]<=Pix_278;PixelsStore[279]<=Pix_279;PixelsStore[280]<=Pix_280;PixelsStore[281]<=Pix_281;PixelsStore[282]<=Pix_282;PixelsStore[283]<=Pix_283;PixelsStore[284]<=Pix_284;PixelsStore[285]<=Pix_285;PixelsStore[286]<=Pix_286;PixelsStore[287]<=Pix_287;PixelsStore[288]<=Pix_288;PixelsStore[289]<=Pix_289;PixelsStore[290]<=Pix_290;PixelsStore[291]<=Pix_291;PixelsStore[292]<=Pix_292;PixelsStore[293]<=Pix_293;PixelsStore[294]<=Pix_294;PixelsStore[295]<=Pix_295;PixelsStore[296]<=Pix_296;PixelsStore[297]<=Pix_297;PixelsStore[298]<=Pix_298;PixelsStore[299]<=Pix_299;PixelsStore[300]<=Pix_300;PixelsStore[301]<=Pix_301;PixelsStore[302]<=Pix_302;PixelsStore[303]<=Pix_303;PixelsStore[304]<=Pix_304;PixelsStore[305]<=Pix_305;PixelsStore[306]<=Pix_306;PixelsStore[307]<=Pix_307;PixelsStore[308]<=Pix_308;PixelsStore[309]<=Pix_309;PixelsStore[310]<=Pix_310;PixelsStore[311]<=Pix_311;PixelsStore[312]<=Pix_312;PixelsStore[313]<=Pix_313;PixelsStore[314]<=Pix_314;PixelsStore[315]<=Pix_315;PixelsStore[316]<=Pix_316;PixelsStore[317]<=Pix_317;PixelsStore[318]<=Pix_318;PixelsStore[319]<=Pix_319;PixelsStore[320]<=Pix_320;PixelsStore[321]<=Pix_321;PixelsStore[322]<=Pix_322;PixelsStore[323]<=Pix_323;PixelsStore[324]<=Pix_324;PixelsStore[325]<=Pix_325;PixelsStore[326]<=Pix_326;PixelsStore[327]<=Pix_327;PixelsStore[328]<=Pix_328;PixelsStore[329]<=Pix_329;PixelsStore[330]<=Pix_330;PixelsStore[331]<=Pix_331;PixelsStore[332]<=Pix_332;PixelsStore[333]<=Pix_333;PixelsStore[334]<=Pix_334;PixelsStore[335]<=Pix_335;PixelsStore[336]<=Pix_336;PixelsStore[337]<=Pix_337;PixelsStore[338]<=Pix_338;PixelsStore[339]<=Pix_339;PixelsStore[340]<=Pix_340;PixelsStore[341]<=Pix_341;PixelsStore[342]<=Pix_342;PixelsStore[343]<=Pix_343;PixelsStore[344]<=Pix_344;PixelsStore[345]<=Pix_345;PixelsStore[346]<=Pix_346;PixelsStore[347]<=Pix_347;PixelsStore[348]<=Pix_348;PixelsStore[349]<=Pix_349;PixelsStore[350]<=Pix_350;PixelsStore[351]<=Pix_351;PixelsStore[352]<=Pix_352;PixelsStore[353]<=Pix_353;PixelsStore[354]<=Pix_354;PixelsStore[355]<=Pix_355;PixelsStore[356]<=Pix_356;PixelsStore[357]<=Pix_357;PixelsStore[358]<=Pix_358;PixelsStore[359]<=Pix_359;PixelsStore[360]<=Pix_360;PixelsStore[361]<=Pix_361;PixelsStore[362]<=Pix_362;PixelsStore[363]<=Pix_363;PixelsStore[364]<=Pix_364;PixelsStore[365]<=Pix_365;PixelsStore[366]<=Pix_366;PixelsStore[367]<=Pix_367;PixelsStore[368]<=Pix_368;PixelsStore[369]<=Pix_369;PixelsStore[370]<=Pix_370;PixelsStore[371]<=Pix_371;PixelsStore[372]<=Pix_372;PixelsStore[373]<=Pix_373;PixelsStore[374]<=Pix_374;PixelsStore[375]<=Pix_375;PixelsStore[376]<=Pix_376;PixelsStore[377]<=Pix_377;PixelsStore[378]<=Pix_378;PixelsStore[379]<=Pix_379;PixelsStore[380]<=Pix_380;PixelsStore[381]<=Pix_381;PixelsStore[382]<=Pix_382;PixelsStore[383]<=Pix_383;PixelsStore[384]<=Pix_384;PixelsStore[385]<=Pix_385;PixelsStore[386]<=Pix_386;PixelsStore[387]<=Pix_387;PixelsStore[388]<=Pix_388;PixelsStore[389]<=Pix_389;PixelsStore[390]<=Pix_390;PixelsStore[391]<=Pix_391;PixelsStore[392]<=Pix_392;PixelsStore[393]<=Pix_393;PixelsStore[394]<=Pix_394;PixelsStore[395]<=Pix_395;PixelsStore[396]<=Pix_396;PixelsStore[397]<=Pix_397;PixelsStore[398]<=Pix_398;PixelsStore[399]<=Pix_399;PixelsStore[400]<=Pix_400;PixelsStore[401]<=Pix_401;PixelsStore[402]<=Pix_402;PixelsStore[403]<=Pix_403;PixelsStore[404]<=Pix_404;PixelsStore[405]<=Pix_405;PixelsStore[406]<=Pix_406;PixelsStore[407]<=Pix_407;PixelsStore[408]<=Pix_408;PixelsStore[409]<=Pix_409;PixelsStore[410]<=Pix_410;PixelsStore[411]<=Pix_411;PixelsStore[412]<=Pix_412;PixelsStore[413]<=Pix_413;PixelsStore[414]<=Pix_414;PixelsStore[415]<=Pix_415;PixelsStore[416]<=Pix_416;PixelsStore[417]<=Pix_417;PixelsStore[418]<=Pix_418;PixelsStore[419]<=Pix_419;PixelsStore[420]<=Pix_420;PixelsStore[421]<=Pix_421;PixelsStore[422]<=Pix_422;PixelsStore[423]<=Pix_423;PixelsStore[424]<=Pix_424;PixelsStore[425]<=Pix_425;PixelsStore[426]<=Pix_426;PixelsStore[427]<=Pix_427;PixelsStore[428]<=Pix_428;PixelsStore[429]<=Pix_429;PixelsStore[430]<=Pix_430;PixelsStore[431]<=Pix_431;PixelsStore[432]<=Pix_432;PixelsStore[433]<=Pix_433;PixelsStore[434]<=Pix_434;PixelsStore[435]<=Pix_435;PixelsStore[436]<=Pix_436;PixelsStore[437]<=Pix_437;PixelsStore[438]<=Pix_438;PixelsStore[439]<=Pix_439;PixelsStore[440]<=Pix_440;PixelsStore[441]<=Pix_441;PixelsStore[442]<=Pix_442;PixelsStore[443]<=Pix_443;PixelsStore[444]<=Pix_444;PixelsStore[445]<=Pix_445;PixelsStore[446]<=Pix_446;PixelsStore[447]<=Pix_447;PixelsStore[448]<=Pix_448;PixelsStore[449]<=Pix_449;PixelsStore[450]<=Pix_450;PixelsStore[451]<=Pix_451;PixelsStore[452]<=Pix_452;PixelsStore[453]<=Pix_453;PixelsStore[454]<=Pix_454;PixelsStore[455]<=Pix_455;PixelsStore[456]<=Pix_456;PixelsStore[457]<=Pix_457;PixelsStore[458]<=Pix_458;PixelsStore[459]<=Pix_459;PixelsStore[460]<=Pix_460;PixelsStore[461]<=Pix_461;PixelsStore[462]<=Pix_462;PixelsStore[463]<=Pix_463;PixelsStore[464]<=Pix_464;PixelsStore[465]<=Pix_465;PixelsStore[466]<=Pix_466;PixelsStore[467]<=Pix_467;PixelsStore[468]<=Pix_468;PixelsStore[469]<=Pix_469;PixelsStore[470]<=Pix_470;PixelsStore[471]<=Pix_471;PixelsStore[472]<=Pix_472;PixelsStore[473]<=Pix_473;PixelsStore[474]<=Pix_474;PixelsStore[475]<=Pix_475;PixelsStore[476]<=Pix_476;PixelsStore[477]<=Pix_477;PixelsStore[478]<=Pix_478;PixelsStore[479]<=Pix_479;PixelsStore[480]<=Pix_480;PixelsStore[481]<=Pix_481;PixelsStore[482]<=Pix_482;PixelsStore[483]<=Pix_483;PixelsStore[484]<=Pix_484;PixelsStore[485]<=Pix_485;PixelsStore[486]<=Pix_486;PixelsStore[487]<=Pix_487;PixelsStore[488]<=Pix_488;PixelsStore[489]<=Pix_489;PixelsStore[490]<=Pix_490;PixelsStore[491]<=Pix_491;PixelsStore[492]<=Pix_492;PixelsStore[493]<=Pix_493;PixelsStore[494]<=Pix_494;PixelsStore[495]<=Pix_495;PixelsStore[496]<=Pix_496;PixelsStore[497]<=Pix_497;PixelsStore[498]<=Pix_498;PixelsStore[499]<=Pix_499;PixelsStore[500]<=Pix_500;PixelsStore[501]<=Pix_501;PixelsStore[502]<=Pix_502;PixelsStore[503]<=Pix_503;PixelsStore[504]<=Pix_504;PixelsStore[505]<=Pix_505;PixelsStore[506]<=Pix_506;PixelsStore[507]<=Pix_507;PixelsStore[508]<=Pix_508;PixelsStore[509]<=Pix_509;PixelsStore[510]<=Pix_510;PixelsStore[511]<=Pix_511;PixelsStore[512]<=Pix_512;PixelsStore[513]<=Pix_513;PixelsStore[514]<=Pix_514;PixelsStore[515]<=Pix_515;PixelsStore[516]<=Pix_516;PixelsStore[517]<=Pix_517;PixelsStore[518]<=Pix_518;PixelsStore[519]<=Pix_519;PixelsStore[520]<=Pix_520;PixelsStore[521]<=Pix_521;PixelsStore[522]<=Pix_522;PixelsStore[523]<=Pix_523;PixelsStore[524]<=Pix_524;PixelsStore[525]<=Pix_525;PixelsStore[526]<=Pix_526;PixelsStore[527]<=Pix_527;PixelsStore[528]<=Pix_528;PixelsStore[529]<=Pix_529;PixelsStore[530]<=Pix_530;PixelsStore[531]<=Pix_531;PixelsStore[532]<=Pix_532;PixelsStore[533]<=Pix_533;PixelsStore[534]<=Pix_534;PixelsStore[535]<=Pix_535;PixelsStore[536]<=Pix_536;PixelsStore[537]<=Pix_537;PixelsStore[538]<=Pix_538;PixelsStore[539]<=Pix_539;PixelsStore[540]<=Pix_540;PixelsStore[541]<=Pix_541;PixelsStore[542]<=Pix_542;PixelsStore[543]<=Pix_543;PixelsStore[544]<=Pix_544;PixelsStore[545]<=Pix_545;PixelsStore[546]<=Pix_546;PixelsStore[547]<=Pix_547;PixelsStore[548]<=Pix_548;PixelsStore[549]<=Pix_549;PixelsStore[550]<=Pix_550;PixelsStore[551]<=Pix_551;PixelsStore[552]<=Pix_552;PixelsStore[553]<=Pix_553;PixelsStore[554]<=Pix_554;PixelsStore[555]<=Pix_555;PixelsStore[556]<=Pix_556;PixelsStore[557]<=Pix_557;PixelsStore[558]<=Pix_558;PixelsStore[559]<=Pix_559;PixelsStore[560]<=Pix_560;PixelsStore[561]<=Pix_561;PixelsStore[562]<=Pix_562;PixelsStore[563]<=Pix_563;PixelsStore[564]<=Pix_564;PixelsStore[565]<=Pix_565;PixelsStore[566]<=Pix_566;PixelsStore[567]<=Pix_567;PixelsStore[568]<=Pix_568;PixelsStore[569]<=Pix_569;PixelsStore[570]<=Pix_570;PixelsStore[571]<=Pix_571;PixelsStore[572]<=Pix_572;PixelsStore[573]<=Pix_573;PixelsStore[574]<=Pix_574;PixelsStore[575]<=Pix_575;PixelsStore[576]<=Pix_576;PixelsStore[577]<=Pix_577;PixelsStore[578]<=Pix_578;PixelsStore[579]<=Pix_579;PixelsStore[580]<=Pix_580;PixelsStore[581]<=Pix_581;PixelsStore[582]<=Pix_582;PixelsStore[583]<=Pix_583;PixelsStore[584]<=Pix_584;PixelsStore[585]<=Pix_585;PixelsStore[586]<=Pix_586;PixelsStore[587]<=Pix_587;PixelsStore[588]<=Pix_588;PixelsStore[589]<=Pix_589;PixelsStore[590]<=Pix_590;PixelsStore[591]<=Pix_591;PixelsStore[592]<=Pix_592;PixelsStore[593]<=Pix_593;PixelsStore[594]<=Pix_594;PixelsStore[595]<=Pix_595;PixelsStore[596]<=Pix_596;PixelsStore[597]<=Pix_597;PixelsStore[598]<=Pix_598;PixelsStore[599]<=Pix_599;PixelsStore[600]<=Pix_600;PixelsStore[601]<=Pix_601;PixelsStore[602]<=Pix_602;PixelsStore[603]<=Pix_603;PixelsStore[604]<=Pix_604;PixelsStore[605]<=Pix_605;PixelsStore[606]<=Pix_606;PixelsStore[607]<=Pix_607;PixelsStore[608]<=Pix_608;PixelsStore[609]<=Pix_609;PixelsStore[610]<=Pix_610;PixelsStore[611]<=Pix_611;PixelsStore[612]<=Pix_612;PixelsStore[613]<=Pix_613;PixelsStore[614]<=Pix_614;PixelsStore[615]<=Pix_615;PixelsStore[616]<=Pix_616;PixelsStore[617]<=Pix_617;PixelsStore[618]<=Pix_618;PixelsStore[619]<=Pix_619;PixelsStore[620]<=Pix_620;PixelsStore[621]<=Pix_621;PixelsStore[622]<=Pix_622;PixelsStore[623]<=Pix_623;PixelsStore[624]<=Pix_624;PixelsStore[625]<=Pix_625;PixelsStore[626]<=Pix_626;PixelsStore[627]<=Pix_627;PixelsStore[628]<=Pix_628;PixelsStore[629]<=Pix_629;PixelsStore[630]<=Pix_630;PixelsStore[631]<=Pix_631;PixelsStore[632]<=Pix_632;PixelsStore[633]<=Pix_633;PixelsStore[634]<=Pix_634;PixelsStore[635]<=Pix_635;PixelsStore[636]<=Pix_636;PixelsStore[637]<=Pix_637;PixelsStore[638]<=Pix_638;PixelsStore[639]<=Pix_639;PixelsStore[640]<=Pix_640;PixelsStore[641]<=Pix_641;PixelsStore[642]<=Pix_642;PixelsStore[643]<=Pix_643;PixelsStore[644]<=Pix_644;PixelsStore[645]<=Pix_645;PixelsStore[646]<=Pix_646;PixelsStore[647]<=Pix_647;PixelsStore[648]<=Pix_648;PixelsStore[649]<=Pix_649;PixelsStore[650]<=Pix_650;PixelsStore[651]<=Pix_651;PixelsStore[652]<=Pix_652;PixelsStore[653]<=Pix_653;PixelsStore[654]<=Pix_654;PixelsStore[655]<=Pix_655;PixelsStore[656]<=Pix_656;PixelsStore[657]<=Pix_657;PixelsStore[658]<=Pix_658;PixelsStore[659]<=Pix_659;PixelsStore[660]<=Pix_660;PixelsStore[661]<=Pix_661;PixelsStore[662]<=Pix_662;PixelsStore[663]<=Pix_663;PixelsStore[664]<=Pix_664;PixelsStore[665]<=Pix_665;PixelsStore[666]<=Pix_666;PixelsStore[667]<=Pix_667;PixelsStore[668]<=Pix_668;PixelsStore[669]<=Pix_669;PixelsStore[670]<=Pix_670;PixelsStore[671]<=Pix_671;PixelsStore[672]<=Pix_672;PixelsStore[673]<=Pix_673;PixelsStore[674]<=Pix_674;PixelsStore[675]<=Pix_675;PixelsStore[676]<=Pix_676;PixelsStore[677]<=Pix_677;PixelsStore[678]<=Pix_678;PixelsStore[679]<=Pix_679;PixelsStore[680]<=Pix_680;PixelsStore[681]<=Pix_681;PixelsStore[682]<=Pix_682;PixelsStore[683]<=Pix_683;PixelsStore[684]<=Pix_684;PixelsStore[685]<=Pix_685;PixelsStore[686]<=Pix_686;PixelsStore[687]<=Pix_687;PixelsStore[688]<=Pix_688;PixelsStore[689]<=Pix_689;PixelsStore[690]<=Pix_690;PixelsStore[691]<=Pix_691;PixelsStore[692]<=Pix_692;PixelsStore[693]<=Pix_693;PixelsStore[694]<=Pix_694;PixelsStore[695]<=Pix_695;PixelsStore[696]<=Pix_696;PixelsStore[697]<=Pix_697;PixelsStore[698]<=Pix_698;PixelsStore[699]<=Pix_699;PixelsStore[700]<=Pix_700;PixelsStore[701]<=Pix_701;PixelsStore[702]<=Pix_702;PixelsStore[703]<=Pix_703;PixelsStore[704]<=Pix_704;PixelsStore[705]<=Pix_705;PixelsStore[706]<=Pix_706;PixelsStore[707]<=Pix_707;PixelsStore[708]<=Pix_708;PixelsStore[709]<=Pix_709;PixelsStore[710]<=Pix_710;PixelsStore[711]<=Pix_711;PixelsStore[712]<=Pix_712;PixelsStore[713]<=Pix_713;PixelsStore[714]<=Pix_714;PixelsStore[715]<=Pix_715;PixelsStore[716]<=Pix_716;PixelsStore[717]<=Pix_717;PixelsStore[718]<=Pix_718;PixelsStore[719]<=Pix_719;PixelsStore[720]<=Pix_720;PixelsStore[721]<=Pix_721;PixelsStore[722]<=Pix_722;PixelsStore[723]<=Pix_723;PixelsStore[724]<=Pix_724;PixelsStore[725]<=Pix_725;PixelsStore[726]<=Pix_726;PixelsStore[727]<=Pix_727;PixelsStore[728]<=Pix_728;PixelsStore[729]<=Pix_729;PixelsStore[730]<=Pix_730;PixelsStore[731]<=Pix_731;PixelsStore[732]<=Pix_732;PixelsStore[733]<=Pix_733;PixelsStore[734]<=Pix_734;PixelsStore[735]<=Pix_735;PixelsStore[736]<=Pix_736;PixelsStore[737]<=Pix_737;PixelsStore[738]<=Pix_738;PixelsStore[739]<=Pix_739;PixelsStore[740]<=Pix_740;PixelsStore[741]<=Pix_741;PixelsStore[742]<=Pix_742;PixelsStore[743]<=Pix_743;PixelsStore[744]<=Pix_744;PixelsStore[745]<=Pix_745;PixelsStore[746]<=Pix_746;PixelsStore[747]<=Pix_747;PixelsStore[748]<=Pix_748;PixelsStore[749]<=Pix_749;PixelsStore[750]<=Pix_750;PixelsStore[751]<=Pix_751;PixelsStore[752]<=Pix_752;PixelsStore[753]<=Pix_753;PixelsStore[754]<=Pix_754;PixelsStore[755]<=Pix_755;PixelsStore[756]<=Pix_756;PixelsStore[757]<=Pix_757;PixelsStore[758]<=Pix_758;PixelsStore[759]<=Pix_759;PixelsStore[760]<=Pix_760;PixelsStore[761]<=Pix_761;PixelsStore[762]<=Pix_762;PixelsStore[763]<=Pix_763;PixelsStore[764]<=Pix_764;PixelsStore[765]<=Pix_765;PixelsStore[766]<=Pix_766;PixelsStore[767]<=Pix_767;PixelsStore[768]<=Pix_768;PixelsStore[769]<=Pix_769;PixelsStore[770]<=Pix_770;PixelsStore[771]<=Pix_771;PixelsStore[772]<=Pix_772;PixelsStore[773]<=Pix_773;PixelsStore[774]<=Pix_774;PixelsStore[775]<=Pix_775;PixelsStore[776]<=Pix_776;PixelsStore[777]<=Pix_777;PixelsStore[778]<=Pix_778;PixelsStore[779]<=Pix_779;PixelsStore[780]<=Pix_780;PixelsStore[781]<=Pix_781;PixelsStore[782]<=Pix_782;PixelsStore[783]<=Pix_783;PixelsStore[784]<=Pix_784;
		WeightsStore[0][0]<=Wgt_0_0;WeightsStore[0][1]<=Wgt_0_1;WeightsStore[0][2]<=Wgt_0_2;WeightsStore[0][3]<=Wgt_0_3;WeightsStore[0][4]<=Wgt_0_4;WeightsStore[0][5]<=Wgt_0_5;WeightsStore[0][6]<=Wgt_0_6;WeightsStore[0][7]<=Wgt_0_7;WeightsStore[0][8]<=Wgt_0_8;WeightsStore[0][9]<=Wgt_0_9;WeightsStore[0][10]<=Wgt_0_10;WeightsStore[0][11]<=Wgt_0_11;WeightsStore[0][12]<=Wgt_0_12;WeightsStore[0][13]<=Wgt_0_13;WeightsStore[0][14]<=Wgt_0_14;WeightsStore[0][15]<=Wgt_0_15;WeightsStore[0][16]<=Wgt_0_16;WeightsStore[0][17]<=Wgt_0_17;WeightsStore[0][18]<=Wgt_0_18;WeightsStore[0][19]<=Wgt_0_19;WeightsStore[0][20]<=Wgt_0_20;WeightsStore[0][21]<=Wgt_0_21;WeightsStore[0][22]<=Wgt_0_22;WeightsStore[0][23]<=Wgt_0_23;WeightsStore[0][24]<=Wgt_0_24;WeightsStore[0][25]<=Wgt_0_25;WeightsStore[0][26]<=Wgt_0_26;WeightsStore[0][27]<=Wgt_0_27;WeightsStore[0][28]<=Wgt_0_28;WeightsStore[0][29]<=Wgt_0_29;WeightsStore[0][30]<=Wgt_0_30;WeightsStore[0][31]<=Wgt_0_31;WeightsStore[0][32]<=Wgt_0_32;WeightsStore[0][33]<=Wgt_0_33;WeightsStore[0][34]<=Wgt_0_34;WeightsStore[0][35]<=Wgt_0_35;WeightsStore[0][36]<=Wgt_0_36;WeightsStore[0][37]<=Wgt_0_37;WeightsStore[0][38]<=Wgt_0_38;WeightsStore[0][39]<=Wgt_0_39;WeightsStore[0][40]<=Wgt_0_40;WeightsStore[0][41]<=Wgt_0_41;WeightsStore[0][42]<=Wgt_0_42;WeightsStore[0][43]<=Wgt_0_43;WeightsStore[0][44]<=Wgt_0_44;WeightsStore[0][45]<=Wgt_0_45;WeightsStore[0][46]<=Wgt_0_46;WeightsStore[0][47]<=Wgt_0_47;WeightsStore[0][48]<=Wgt_0_48;WeightsStore[0][49]<=Wgt_0_49;WeightsStore[0][50]<=Wgt_0_50;WeightsStore[0][51]<=Wgt_0_51;WeightsStore[0][52]<=Wgt_0_52;WeightsStore[0][53]<=Wgt_0_53;WeightsStore[0][54]<=Wgt_0_54;WeightsStore[0][55]<=Wgt_0_55;WeightsStore[0][56]<=Wgt_0_56;WeightsStore[0][57]<=Wgt_0_57;WeightsStore[0][58]<=Wgt_0_58;WeightsStore[0][59]<=Wgt_0_59;WeightsStore[0][60]<=Wgt_0_60;WeightsStore[0][61]<=Wgt_0_61;WeightsStore[0][62]<=Wgt_0_62;WeightsStore[0][63]<=Wgt_0_63;WeightsStore[0][64]<=Wgt_0_64;WeightsStore[0][65]<=Wgt_0_65;WeightsStore[0][66]<=Wgt_0_66;WeightsStore[0][67]<=Wgt_0_67;WeightsStore[0][68]<=Wgt_0_68;WeightsStore[0][69]<=Wgt_0_69;WeightsStore[0][70]<=Wgt_0_70;WeightsStore[0][71]<=Wgt_0_71;WeightsStore[0][72]<=Wgt_0_72;WeightsStore[0][73]<=Wgt_0_73;WeightsStore[0][74]<=Wgt_0_74;WeightsStore[0][75]<=Wgt_0_75;WeightsStore[0][76]<=Wgt_0_76;WeightsStore[0][77]<=Wgt_0_77;WeightsStore[0][78]<=Wgt_0_78;WeightsStore[0][79]<=Wgt_0_79;WeightsStore[0][80]<=Wgt_0_80;WeightsStore[0][81]<=Wgt_0_81;WeightsStore[0][82]<=Wgt_0_82;WeightsStore[0][83]<=Wgt_0_83;WeightsStore[0][84]<=Wgt_0_84;WeightsStore[0][85]<=Wgt_0_85;WeightsStore[0][86]<=Wgt_0_86;WeightsStore[0][87]<=Wgt_0_87;WeightsStore[0][88]<=Wgt_0_88;WeightsStore[0][89]<=Wgt_0_89;WeightsStore[0][90]<=Wgt_0_90;WeightsStore[0][91]<=Wgt_0_91;WeightsStore[0][92]<=Wgt_0_92;WeightsStore[0][93]<=Wgt_0_93;WeightsStore[0][94]<=Wgt_0_94;WeightsStore[0][95]<=Wgt_0_95;WeightsStore[0][96]<=Wgt_0_96;WeightsStore[0][97]<=Wgt_0_97;WeightsStore[0][98]<=Wgt_0_98;WeightsStore[0][99]<=Wgt_0_99;WeightsStore[0][100]<=Wgt_0_100;WeightsStore[0][101]<=Wgt_0_101;WeightsStore[0][102]<=Wgt_0_102;WeightsStore[0][103]<=Wgt_0_103;WeightsStore[0][104]<=Wgt_0_104;WeightsStore[0][105]<=Wgt_0_105;WeightsStore[0][106]<=Wgt_0_106;WeightsStore[0][107]<=Wgt_0_107;WeightsStore[0][108]<=Wgt_0_108;WeightsStore[0][109]<=Wgt_0_109;WeightsStore[0][110]<=Wgt_0_110;WeightsStore[0][111]<=Wgt_0_111;WeightsStore[0][112]<=Wgt_0_112;WeightsStore[0][113]<=Wgt_0_113;WeightsStore[0][114]<=Wgt_0_114;WeightsStore[0][115]<=Wgt_0_115;WeightsStore[0][116]<=Wgt_0_116;WeightsStore[0][117]<=Wgt_0_117;WeightsStore[0][118]<=Wgt_0_118;WeightsStore[0][119]<=Wgt_0_119;WeightsStore[0][120]<=Wgt_0_120;WeightsStore[0][121]<=Wgt_0_121;WeightsStore[0][122]<=Wgt_0_122;WeightsStore[0][123]<=Wgt_0_123;WeightsStore[0][124]<=Wgt_0_124;WeightsStore[0][125]<=Wgt_0_125;WeightsStore[0][126]<=Wgt_0_126;WeightsStore[0][127]<=Wgt_0_127;WeightsStore[0][128]<=Wgt_0_128;WeightsStore[0][129]<=Wgt_0_129;WeightsStore[0][130]<=Wgt_0_130;WeightsStore[0][131]<=Wgt_0_131;WeightsStore[0][132]<=Wgt_0_132;WeightsStore[0][133]<=Wgt_0_133;WeightsStore[0][134]<=Wgt_0_134;WeightsStore[0][135]<=Wgt_0_135;WeightsStore[0][136]<=Wgt_0_136;WeightsStore[0][137]<=Wgt_0_137;WeightsStore[0][138]<=Wgt_0_138;WeightsStore[0][139]<=Wgt_0_139;WeightsStore[0][140]<=Wgt_0_140;WeightsStore[0][141]<=Wgt_0_141;WeightsStore[0][142]<=Wgt_0_142;WeightsStore[0][143]<=Wgt_0_143;WeightsStore[0][144]<=Wgt_0_144;WeightsStore[0][145]<=Wgt_0_145;WeightsStore[0][146]<=Wgt_0_146;WeightsStore[0][147]<=Wgt_0_147;WeightsStore[0][148]<=Wgt_0_148;WeightsStore[0][149]<=Wgt_0_149;WeightsStore[0][150]<=Wgt_0_150;WeightsStore[0][151]<=Wgt_0_151;WeightsStore[0][152]<=Wgt_0_152;WeightsStore[0][153]<=Wgt_0_153;WeightsStore[0][154]<=Wgt_0_154;WeightsStore[0][155]<=Wgt_0_155;WeightsStore[0][156]<=Wgt_0_156;WeightsStore[0][157]<=Wgt_0_157;WeightsStore[0][158]<=Wgt_0_158;WeightsStore[0][159]<=Wgt_0_159;WeightsStore[0][160]<=Wgt_0_160;WeightsStore[0][161]<=Wgt_0_161;WeightsStore[0][162]<=Wgt_0_162;WeightsStore[0][163]<=Wgt_0_163;WeightsStore[0][164]<=Wgt_0_164;WeightsStore[0][165]<=Wgt_0_165;WeightsStore[0][166]<=Wgt_0_166;WeightsStore[0][167]<=Wgt_0_167;WeightsStore[0][168]<=Wgt_0_168;WeightsStore[0][169]<=Wgt_0_169;WeightsStore[0][170]<=Wgt_0_170;WeightsStore[0][171]<=Wgt_0_171;WeightsStore[0][172]<=Wgt_0_172;WeightsStore[0][173]<=Wgt_0_173;WeightsStore[0][174]<=Wgt_0_174;WeightsStore[0][175]<=Wgt_0_175;WeightsStore[0][176]<=Wgt_0_176;WeightsStore[0][177]<=Wgt_0_177;WeightsStore[0][178]<=Wgt_0_178;WeightsStore[0][179]<=Wgt_0_179;WeightsStore[0][180]<=Wgt_0_180;WeightsStore[0][181]<=Wgt_0_181;WeightsStore[0][182]<=Wgt_0_182;WeightsStore[0][183]<=Wgt_0_183;WeightsStore[0][184]<=Wgt_0_184;WeightsStore[0][185]<=Wgt_0_185;WeightsStore[0][186]<=Wgt_0_186;WeightsStore[0][187]<=Wgt_0_187;WeightsStore[0][188]<=Wgt_0_188;WeightsStore[0][189]<=Wgt_0_189;WeightsStore[0][190]<=Wgt_0_190;WeightsStore[0][191]<=Wgt_0_191;WeightsStore[0][192]<=Wgt_0_192;WeightsStore[0][193]<=Wgt_0_193;WeightsStore[0][194]<=Wgt_0_194;WeightsStore[0][195]<=Wgt_0_195;WeightsStore[0][196]<=Wgt_0_196;WeightsStore[0][197]<=Wgt_0_197;WeightsStore[0][198]<=Wgt_0_198;WeightsStore[0][199]<=Wgt_0_199;WeightsStore[0][200]<=Wgt_0_200;WeightsStore[0][201]<=Wgt_0_201;WeightsStore[0][202]<=Wgt_0_202;WeightsStore[0][203]<=Wgt_0_203;WeightsStore[0][204]<=Wgt_0_204;WeightsStore[0][205]<=Wgt_0_205;WeightsStore[0][206]<=Wgt_0_206;WeightsStore[0][207]<=Wgt_0_207;WeightsStore[0][208]<=Wgt_0_208;WeightsStore[0][209]<=Wgt_0_209;WeightsStore[0][210]<=Wgt_0_210;WeightsStore[0][211]<=Wgt_0_211;WeightsStore[0][212]<=Wgt_0_212;WeightsStore[0][213]<=Wgt_0_213;WeightsStore[0][214]<=Wgt_0_214;WeightsStore[0][215]<=Wgt_0_215;WeightsStore[0][216]<=Wgt_0_216;WeightsStore[0][217]<=Wgt_0_217;WeightsStore[0][218]<=Wgt_0_218;WeightsStore[0][219]<=Wgt_0_219;WeightsStore[0][220]<=Wgt_0_220;WeightsStore[0][221]<=Wgt_0_221;WeightsStore[0][222]<=Wgt_0_222;WeightsStore[0][223]<=Wgt_0_223;WeightsStore[0][224]<=Wgt_0_224;WeightsStore[0][225]<=Wgt_0_225;WeightsStore[0][226]<=Wgt_0_226;WeightsStore[0][227]<=Wgt_0_227;WeightsStore[0][228]<=Wgt_0_228;WeightsStore[0][229]<=Wgt_0_229;WeightsStore[0][230]<=Wgt_0_230;WeightsStore[0][231]<=Wgt_0_231;WeightsStore[0][232]<=Wgt_0_232;WeightsStore[0][233]<=Wgt_0_233;WeightsStore[0][234]<=Wgt_0_234;WeightsStore[0][235]<=Wgt_0_235;WeightsStore[0][236]<=Wgt_0_236;WeightsStore[0][237]<=Wgt_0_237;WeightsStore[0][238]<=Wgt_0_238;WeightsStore[0][239]<=Wgt_0_239;WeightsStore[0][240]<=Wgt_0_240;WeightsStore[0][241]<=Wgt_0_241;WeightsStore[0][242]<=Wgt_0_242;WeightsStore[0][243]<=Wgt_0_243;WeightsStore[0][244]<=Wgt_0_244;WeightsStore[0][245]<=Wgt_0_245;WeightsStore[0][246]<=Wgt_0_246;WeightsStore[0][247]<=Wgt_0_247;WeightsStore[0][248]<=Wgt_0_248;WeightsStore[0][249]<=Wgt_0_249;WeightsStore[0][250]<=Wgt_0_250;WeightsStore[0][251]<=Wgt_0_251;WeightsStore[0][252]<=Wgt_0_252;WeightsStore[0][253]<=Wgt_0_253;WeightsStore[0][254]<=Wgt_0_254;WeightsStore[0][255]<=Wgt_0_255;WeightsStore[0][256]<=Wgt_0_256;WeightsStore[0][257]<=Wgt_0_257;WeightsStore[0][258]<=Wgt_0_258;WeightsStore[0][259]<=Wgt_0_259;WeightsStore[0][260]<=Wgt_0_260;WeightsStore[0][261]<=Wgt_0_261;WeightsStore[0][262]<=Wgt_0_262;WeightsStore[0][263]<=Wgt_0_263;WeightsStore[0][264]<=Wgt_0_264;WeightsStore[0][265]<=Wgt_0_265;WeightsStore[0][266]<=Wgt_0_266;WeightsStore[0][267]<=Wgt_0_267;WeightsStore[0][268]<=Wgt_0_268;WeightsStore[0][269]<=Wgt_0_269;WeightsStore[0][270]<=Wgt_0_270;WeightsStore[0][271]<=Wgt_0_271;WeightsStore[0][272]<=Wgt_0_272;WeightsStore[0][273]<=Wgt_0_273;WeightsStore[0][274]<=Wgt_0_274;WeightsStore[0][275]<=Wgt_0_275;WeightsStore[0][276]<=Wgt_0_276;WeightsStore[0][277]<=Wgt_0_277;WeightsStore[0][278]<=Wgt_0_278;WeightsStore[0][279]<=Wgt_0_279;WeightsStore[0][280]<=Wgt_0_280;WeightsStore[0][281]<=Wgt_0_281;WeightsStore[0][282]<=Wgt_0_282;WeightsStore[0][283]<=Wgt_0_283;WeightsStore[0][284]<=Wgt_0_284;WeightsStore[0][285]<=Wgt_0_285;WeightsStore[0][286]<=Wgt_0_286;WeightsStore[0][287]<=Wgt_0_287;WeightsStore[0][288]<=Wgt_0_288;WeightsStore[0][289]<=Wgt_0_289;WeightsStore[0][290]<=Wgt_0_290;WeightsStore[0][291]<=Wgt_0_291;WeightsStore[0][292]<=Wgt_0_292;WeightsStore[0][293]<=Wgt_0_293;WeightsStore[0][294]<=Wgt_0_294;WeightsStore[0][295]<=Wgt_0_295;WeightsStore[0][296]<=Wgt_0_296;WeightsStore[0][297]<=Wgt_0_297;WeightsStore[0][298]<=Wgt_0_298;WeightsStore[0][299]<=Wgt_0_299;WeightsStore[0][300]<=Wgt_0_300;WeightsStore[0][301]<=Wgt_0_301;WeightsStore[0][302]<=Wgt_0_302;WeightsStore[0][303]<=Wgt_0_303;WeightsStore[0][304]<=Wgt_0_304;WeightsStore[0][305]<=Wgt_0_305;WeightsStore[0][306]<=Wgt_0_306;WeightsStore[0][307]<=Wgt_0_307;WeightsStore[0][308]<=Wgt_0_308;WeightsStore[0][309]<=Wgt_0_309;WeightsStore[0][310]<=Wgt_0_310;WeightsStore[0][311]<=Wgt_0_311;WeightsStore[0][312]<=Wgt_0_312;WeightsStore[0][313]<=Wgt_0_313;WeightsStore[0][314]<=Wgt_0_314;WeightsStore[0][315]<=Wgt_0_315;WeightsStore[0][316]<=Wgt_0_316;WeightsStore[0][317]<=Wgt_0_317;WeightsStore[0][318]<=Wgt_0_318;WeightsStore[0][319]<=Wgt_0_319;WeightsStore[0][320]<=Wgt_0_320;WeightsStore[0][321]<=Wgt_0_321;WeightsStore[0][322]<=Wgt_0_322;WeightsStore[0][323]<=Wgt_0_323;WeightsStore[0][324]<=Wgt_0_324;WeightsStore[0][325]<=Wgt_0_325;WeightsStore[0][326]<=Wgt_0_326;WeightsStore[0][327]<=Wgt_0_327;WeightsStore[0][328]<=Wgt_0_328;WeightsStore[0][329]<=Wgt_0_329;WeightsStore[0][330]<=Wgt_0_330;WeightsStore[0][331]<=Wgt_0_331;WeightsStore[0][332]<=Wgt_0_332;WeightsStore[0][333]<=Wgt_0_333;WeightsStore[0][334]<=Wgt_0_334;WeightsStore[0][335]<=Wgt_0_335;WeightsStore[0][336]<=Wgt_0_336;WeightsStore[0][337]<=Wgt_0_337;WeightsStore[0][338]<=Wgt_0_338;WeightsStore[0][339]<=Wgt_0_339;WeightsStore[0][340]<=Wgt_0_340;WeightsStore[0][341]<=Wgt_0_341;WeightsStore[0][342]<=Wgt_0_342;WeightsStore[0][343]<=Wgt_0_343;WeightsStore[0][344]<=Wgt_0_344;WeightsStore[0][345]<=Wgt_0_345;WeightsStore[0][346]<=Wgt_0_346;WeightsStore[0][347]<=Wgt_0_347;WeightsStore[0][348]<=Wgt_0_348;WeightsStore[0][349]<=Wgt_0_349;WeightsStore[0][350]<=Wgt_0_350;WeightsStore[0][351]<=Wgt_0_351;WeightsStore[0][352]<=Wgt_0_352;WeightsStore[0][353]<=Wgt_0_353;WeightsStore[0][354]<=Wgt_0_354;WeightsStore[0][355]<=Wgt_0_355;WeightsStore[0][356]<=Wgt_0_356;WeightsStore[0][357]<=Wgt_0_357;WeightsStore[0][358]<=Wgt_0_358;WeightsStore[0][359]<=Wgt_0_359;WeightsStore[0][360]<=Wgt_0_360;WeightsStore[0][361]<=Wgt_0_361;WeightsStore[0][362]<=Wgt_0_362;WeightsStore[0][363]<=Wgt_0_363;WeightsStore[0][364]<=Wgt_0_364;WeightsStore[0][365]<=Wgt_0_365;WeightsStore[0][366]<=Wgt_0_366;WeightsStore[0][367]<=Wgt_0_367;WeightsStore[0][368]<=Wgt_0_368;WeightsStore[0][369]<=Wgt_0_369;WeightsStore[0][370]<=Wgt_0_370;WeightsStore[0][371]<=Wgt_0_371;WeightsStore[0][372]<=Wgt_0_372;WeightsStore[0][373]<=Wgt_0_373;WeightsStore[0][374]<=Wgt_0_374;WeightsStore[0][375]<=Wgt_0_375;WeightsStore[0][376]<=Wgt_0_376;WeightsStore[0][377]<=Wgt_0_377;WeightsStore[0][378]<=Wgt_0_378;WeightsStore[0][379]<=Wgt_0_379;WeightsStore[0][380]<=Wgt_0_380;WeightsStore[0][381]<=Wgt_0_381;WeightsStore[0][382]<=Wgt_0_382;WeightsStore[0][383]<=Wgt_0_383;WeightsStore[0][384]<=Wgt_0_384;WeightsStore[0][385]<=Wgt_0_385;WeightsStore[0][386]<=Wgt_0_386;WeightsStore[0][387]<=Wgt_0_387;WeightsStore[0][388]<=Wgt_0_388;WeightsStore[0][389]<=Wgt_0_389;WeightsStore[0][390]<=Wgt_0_390;WeightsStore[0][391]<=Wgt_0_391;WeightsStore[0][392]<=Wgt_0_392;WeightsStore[0][393]<=Wgt_0_393;WeightsStore[0][394]<=Wgt_0_394;WeightsStore[0][395]<=Wgt_0_395;WeightsStore[0][396]<=Wgt_0_396;WeightsStore[0][397]<=Wgt_0_397;WeightsStore[0][398]<=Wgt_0_398;WeightsStore[0][399]<=Wgt_0_399;WeightsStore[0][400]<=Wgt_0_400;WeightsStore[0][401]<=Wgt_0_401;WeightsStore[0][402]<=Wgt_0_402;WeightsStore[0][403]<=Wgt_0_403;WeightsStore[0][404]<=Wgt_0_404;WeightsStore[0][405]<=Wgt_0_405;WeightsStore[0][406]<=Wgt_0_406;WeightsStore[0][407]<=Wgt_0_407;WeightsStore[0][408]<=Wgt_0_408;WeightsStore[0][409]<=Wgt_0_409;WeightsStore[0][410]<=Wgt_0_410;WeightsStore[0][411]<=Wgt_0_411;WeightsStore[0][412]<=Wgt_0_412;WeightsStore[0][413]<=Wgt_0_413;WeightsStore[0][414]<=Wgt_0_414;WeightsStore[0][415]<=Wgt_0_415;WeightsStore[0][416]<=Wgt_0_416;WeightsStore[0][417]<=Wgt_0_417;WeightsStore[0][418]<=Wgt_0_418;WeightsStore[0][419]<=Wgt_0_419;WeightsStore[0][420]<=Wgt_0_420;WeightsStore[0][421]<=Wgt_0_421;WeightsStore[0][422]<=Wgt_0_422;WeightsStore[0][423]<=Wgt_0_423;WeightsStore[0][424]<=Wgt_0_424;WeightsStore[0][425]<=Wgt_0_425;WeightsStore[0][426]<=Wgt_0_426;WeightsStore[0][427]<=Wgt_0_427;WeightsStore[0][428]<=Wgt_0_428;WeightsStore[0][429]<=Wgt_0_429;WeightsStore[0][430]<=Wgt_0_430;WeightsStore[0][431]<=Wgt_0_431;WeightsStore[0][432]<=Wgt_0_432;WeightsStore[0][433]<=Wgt_0_433;WeightsStore[0][434]<=Wgt_0_434;WeightsStore[0][435]<=Wgt_0_435;WeightsStore[0][436]<=Wgt_0_436;WeightsStore[0][437]<=Wgt_0_437;WeightsStore[0][438]<=Wgt_0_438;WeightsStore[0][439]<=Wgt_0_439;WeightsStore[0][440]<=Wgt_0_440;WeightsStore[0][441]<=Wgt_0_441;WeightsStore[0][442]<=Wgt_0_442;WeightsStore[0][443]<=Wgt_0_443;WeightsStore[0][444]<=Wgt_0_444;WeightsStore[0][445]<=Wgt_0_445;WeightsStore[0][446]<=Wgt_0_446;WeightsStore[0][447]<=Wgt_0_447;WeightsStore[0][448]<=Wgt_0_448;WeightsStore[0][449]<=Wgt_0_449;WeightsStore[0][450]<=Wgt_0_450;WeightsStore[0][451]<=Wgt_0_451;WeightsStore[0][452]<=Wgt_0_452;WeightsStore[0][453]<=Wgt_0_453;WeightsStore[0][454]<=Wgt_0_454;WeightsStore[0][455]<=Wgt_0_455;WeightsStore[0][456]<=Wgt_0_456;WeightsStore[0][457]<=Wgt_0_457;WeightsStore[0][458]<=Wgt_0_458;WeightsStore[0][459]<=Wgt_0_459;WeightsStore[0][460]<=Wgt_0_460;WeightsStore[0][461]<=Wgt_0_461;WeightsStore[0][462]<=Wgt_0_462;WeightsStore[0][463]<=Wgt_0_463;WeightsStore[0][464]<=Wgt_0_464;WeightsStore[0][465]<=Wgt_0_465;WeightsStore[0][466]<=Wgt_0_466;WeightsStore[0][467]<=Wgt_0_467;WeightsStore[0][468]<=Wgt_0_468;WeightsStore[0][469]<=Wgt_0_469;WeightsStore[0][470]<=Wgt_0_470;WeightsStore[0][471]<=Wgt_0_471;WeightsStore[0][472]<=Wgt_0_472;WeightsStore[0][473]<=Wgt_0_473;WeightsStore[0][474]<=Wgt_0_474;WeightsStore[0][475]<=Wgt_0_475;WeightsStore[0][476]<=Wgt_0_476;WeightsStore[0][477]<=Wgt_0_477;WeightsStore[0][478]<=Wgt_0_478;WeightsStore[0][479]<=Wgt_0_479;WeightsStore[0][480]<=Wgt_0_480;WeightsStore[0][481]<=Wgt_0_481;WeightsStore[0][482]<=Wgt_0_482;WeightsStore[0][483]<=Wgt_0_483;WeightsStore[0][484]<=Wgt_0_484;WeightsStore[0][485]<=Wgt_0_485;WeightsStore[0][486]<=Wgt_0_486;WeightsStore[0][487]<=Wgt_0_487;WeightsStore[0][488]<=Wgt_0_488;WeightsStore[0][489]<=Wgt_0_489;WeightsStore[0][490]<=Wgt_0_490;WeightsStore[0][491]<=Wgt_0_491;WeightsStore[0][492]<=Wgt_0_492;WeightsStore[0][493]<=Wgt_0_493;WeightsStore[0][494]<=Wgt_0_494;WeightsStore[0][495]<=Wgt_0_495;WeightsStore[0][496]<=Wgt_0_496;WeightsStore[0][497]<=Wgt_0_497;WeightsStore[0][498]<=Wgt_0_498;WeightsStore[0][499]<=Wgt_0_499;WeightsStore[0][500]<=Wgt_0_500;WeightsStore[0][501]<=Wgt_0_501;WeightsStore[0][502]<=Wgt_0_502;WeightsStore[0][503]<=Wgt_0_503;WeightsStore[0][504]<=Wgt_0_504;WeightsStore[0][505]<=Wgt_0_505;WeightsStore[0][506]<=Wgt_0_506;WeightsStore[0][507]<=Wgt_0_507;WeightsStore[0][508]<=Wgt_0_508;WeightsStore[0][509]<=Wgt_0_509;WeightsStore[0][510]<=Wgt_0_510;WeightsStore[0][511]<=Wgt_0_511;WeightsStore[0][512]<=Wgt_0_512;WeightsStore[0][513]<=Wgt_0_513;WeightsStore[0][514]<=Wgt_0_514;WeightsStore[0][515]<=Wgt_0_515;WeightsStore[0][516]<=Wgt_0_516;WeightsStore[0][517]<=Wgt_0_517;WeightsStore[0][518]<=Wgt_0_518;WeightsStore[0][519]<=Wgt_0_519;WeightsStore[0][520]<=Wgt_0_520;WeightsStore[0][521]<=Wgt_0_521;WeightsStore[0][522]<=Wgt_0_522;WeightsStore[0][523]<=Wgt_0_523;WeightsStore[0][524]<=Wgt_0_524;WeightsStore[0][525]<=Wgt_0_525;WeightsStore[0][526]<=Wgt_0_526;WeightsStore[0][527]<=Wgt_0_527;WeightsStore[0][528]<=Wgt_0_528;WeightsStore[0][529]<=Wgt_0_529;WeightsStore[0][530]<=Wgt_0_530;WeightsStore[0][531]<=Wgt_0_531;WeightsStore[0][532]<=Wgt_0_532;WeightsStore[0][533]<=Wgt_0_533;WeightsStore[0][534]<=Wgt_0_534;WeightsStore[0][535]<=Wgt_0_535;WeightsStore[0][536]<=Wgt_0_536;WeightsStore[0][537]<=Wgt_0_537;WeightsStore[0][538]<=Wgt_0_538;WeightsStore[0][539]<=Wgt_0_539;WeightsStore[0][540]<=Wgt_0_540;WeightsStore[0][541]<=Wgt_0_541;WeightsStore[0][542]<=Wgt_0_542;WeightsStore[0][543]<=Wgt_0_543;WeightsStore[0][544]<=Wgt_0_544;WeightsStore[0][545]<=Wgt_0_545;WeightsStore[0][546]<=Wgt_0_546;WeightsStore[0][547]<=Wgt_0_547;WeightsStore[0][548]<=Wgt_0_548;WeightsStore[0][549]<=Wgt_0_549;WeightsStore[0][550]<=Wgt_0_550;WeightsStore[0][551]<=Wgt_0_551;WeightsStore[0][552]<=Wgt_0_552;WeightsStore[0][553]<=Wgt_0_553;WeightsStore[0][554]<=Wgt_0_554;WeightsStore[0][555]<=Wgt_0_555;WeightsStore[0][556]<=Wgt_0_556;WeightsStore[0][557]<=Wgt_0_557;WeightsStore[0][558]<=Wgt_0_558;WeightsStore[0][559]<=Wgt_0_559;WeightsStore[0][560]<=Wgt_0_560;WeightsStore[0][561]<=Wgt_0_561;WeightsStore[0][562]<=Wgt_0_562;WeightsStore[0][563]<=Wgt_0_563;WeightsStore[0][564]<=Wgt_0_564;WeightsStore[0][565]<=Wgt_0_565;WeightsStore[0][566]<=Wgt_0_566;WeightsStore[0][567]<=Wgt_0_567;WeightsStore[0][568]<=Wgt_0_568;WeightsStore[0][569]<=Wgt_0_569;WeightsStore[0][570]<=Wgt_0_570;WeightsStore[0][571]<=Wgt_0_571;WeightsStore[0][572]<=Wgt_0_572;WeightsStore[0][573]<=Wgt_0_573;WeightsStore[0][574]<=Wgt_0_574;WeightsStore[0][575]<=Wgt_0_575;WeightsStore[0][576]<=Wgt_0_576;WeightsStore[0][577]<=Wgt_0_577;WeightsStore[0][578]<=Wgt_0_578;WeightsStore[0][579]<=Wgt_0_579;WeightsStore[0][580]<=Wgt_0_580;WeightsStore[0][581]<=Wgt_0_581;WeightsStore[0][582]<=Wgt_0_582;WeightsStore[0][583]<=Wgt_0_583;WeightsStore[0][584]<=Wgt_0_584;WeightsStore[0][585]<=Wgt_0_585;WeightsStore[0][586]<=Wgt_0_586;WeightsStore[0][587]<=Wgt_0_587;WeightsStore[0][588]<=Wgt_0_588;WeightsStore[0][589]<=Wgt_0_589;WeightsStore[0][590]<=Wgt_0_590;WeightsStore[0][591]<=Wgt_0_591;WeightsStore[0][592]<=Wgt_0_592;WeightsStore[0][593]<=Wgt_0_593;WeightsStore[0][594]<=Wgt_0_594;WeightsStore[0][595]<=Wgt_0_595;WeightsStore[0][596]<=Wgt_0_596;WeightsStore[0][597]<=Wgt_0_597;WeightsStore[0][598]<=Wgt_0_598;WeightsStore[0][599]<=Wgt_0_599;WeightsStore[0][600]<=Wgt_0_600;WeightsStore[0][601]<=Wgt_0_601;WeightsStore[0][602]<=Wgt_0_602;WeightsStore[0][603]<=Wgt_0_603;WeightsStore[0][604]<=Wgt_0_604;WeightsStore[0][605]<=Wgt_0_605;WeightsStore[0][606]<=Wgt_0_606;WeightsStore[0][607]<=Wgt_0_607;WeightsStore[0][608]<=Wgt_0_608;WeightsStore[0][609]<=Wgt_0_609;WeightsStore[0][610]<=Wgt_0_610;WeightsStore[0][611]<=Wgt_0_611;WeightsStore[0][612]<=Wgt_0_612;WeightsStore[0][613]<=Wgt_0_613;WeightsStore[0][614]<=Wgt_0_614;WeightsStore[0][615]<=Wgt_0_615;WeightsStore[0][616]<=Wgt_0_616;WeightsStore[0][617]<=Wgt_0_617;WeightsStore[0][618]<=Wgt_0_618;WeightsStore[0][619]<=Wgt_0_619;WeightsStore[0][620]<=Wgt_0_620;WeightsStore[0][621]<=Wgt_0_621;WeightsStore[0][622]<=Wgt_0_622;WeightsStore[0][623]<=Wgt_0_623;WeightsStore[0][624]<=Wgt_0_624;WeightsStore[0][625]<=Wgt_0_625;WeightsStore[0][626]<=Wgt_0_626;WeightsStore[0][627]<=Wgt_0_627;WeightsStore[0][628]<=Wgt_0_628;WeightsStore[0][629]<=Wgt_0_629;WeightsStore[0][630]<=Wgt_0_630;WeightsStore[0][631]<=Wgt_0_631;WeightsStore[0][632]<=Wgt_0_632;WeightsStore[0][633]<=Wgt_0_633;WeightsStore[0][634]<=Wgt_0_634;WeightsStore[0][635]<=Wgt_0_635;WeightsStore[0][636]<=Wgt_0_636;WeightsStore[0][637]<=Wgt_0_637;WeightsStore[0][638]<=Wgt_0_638;WeightsStore[0][639]<=Wgt_0_639;WeightsStore[0][640]<=Wgt_0_640;WeightsStore[0][641]<=Wgt_0_641;WeightsStore[0][642]<=Wgt_0_642;WeightsStore[0][643]<=Wgt_0_643;WeightsStore[0][644]<=Wgt_0_644;WeightsStore[0][645]<=Wgt_0_645;WeightsStore[0][646]<=Wgt_0_646;WeightsStore[0][647]<=Wgt_0_647;WeightsStore[0][648]<=Wgt_0_648;WeightsStore[0][649]<=Wgt_0_649;WeightsStore[0][650]<=Wgt_0_650;WeightsStore[0][651]<=Wgt_0_651;WeightsStore[0][652]<=Wgt_0_652;WeightsStore[0][653]<=Wgt_0_653;WeightsStore[0][654]<=Wgt_0_654;WeightsStore[0][655]<=Wgt_0_655;WeightsStore[0][656]<=Wgt_0_656;WeightsStore[0][657]<=Wgt_0_657;WeightsStore[0][658]<=Wgt_0_658;WeightsStore[0][659]<=Wgt_0_659;WeightsStore[0][660]<=Wgt_0_660;WeightsStore[0][661]<=Wgt_0_661;WeightsStore[0][662]<=Wgt_0_662;WeightsStore[0][663]<=Wgt_0_663;WeightsStore[0][664]<=Wgt_0_664;WeightsStore[0][665]<=Wgt_0_665;WeightsStore[0][666]<=Wgt_0_666;WeightsStore[0][667]<=Wgt_0_667;WeightsStore[0][668]<=Wgt_0_668;WeightsStore[0][669]<=Wgt_0_669;WeightsStore[0][670]<=Wgt_0_670;WeightsStore[0][671]<=Wgt_0_671;WeightsStore[0][672]<=Wgt_0_672;WeightsStore[0][673]<=Wgt_0_673;WeightsStore[0][674]<=Wgt_0_674;WeightsStore[0][675]<=Wgt_0_675;WeightsStore[0][676]<=Wgt_0_676;WeightsStore[0][677]<=Wgt_0_677;WeightsStore[0][678]<=Wgt_0_678;WeightsStore[0][679]<=Wgt_0_679;WeightsStore[0][680]<=Wgt_0_680;WeightsStore[0][681]<=Wgt_0_681;WeightsStore[0][682]<=Wgt_0_682;WeightsStore[0][683]<=Wgt_0_683;WeightsStore[0][684]<=Wgt_0_684;WeightsStore[0][685]<=Wgt_0_685;WeightsStore[0][686]<=Wgt_0_686;WeightsStore[0][687]<=Wgt_0_687;WeightsStore[0][688]<=Wgt_0_688;WeightsStore[0][689]<=Wgt_0_689;WeightsStore[0][690]<=Wgt_0_690;WeightsStore[0][691]<=Wgt_0_691;WeightsStore[0][692]<=Wgt_0_692;WeightsStore[0][693]<=Wgt_0_693;WeightsStore[0][694]<=Wgt_0_694;WeightsStore[0][695]<=Wgt_0_695;WeightsStore[0][696]<=Wgt_0_696;WeightsStore[0][697]<=Wgt_0_697;WeightsStore[0][698]<=Wgt_0_698;WeightsStore[0][699]<=Wgt_0_699;WeightsStore[0][700]<=Wgt_0_700;WeightsStore[0][701]<=Wgt_0_701;WeightsStore[0][702]<=Wgt_0_702;WeightsStore[0][703]<=Wgt_0_703;WeightsStore[0][704]<=Wgt_0_704;WeightsStore[0][705]<=Wgt_0_705;WeightsStore[0][706]<=Wgt_0_706;WeightsStore[0][707]<=Wgt_0_707;WeightsStore[0][708]<=Wgt_0_708;WeightsStore[0][709]<=Wgt_0_709;WeightsStore[0][710]<=Wgt_0_710;WeightsStore[0][711]<=Wgt_0_711;WeightsStore[0][712]<=Wgt_0_712;WeightsStore[0][713]<=Wgt_0_713;WeightsStore[0][714]<=Wgt_0_714;WeightsStore[0][715]<=Wgt_0_715;WeightsStore[0][716]<=Wgt_0_716;WeightsStore[0][717]<=Wgt_0_717;WeightsStore[0][718]<=Wgt_0_718;WeightsStore[0][719]<=Wgt_0_719;WeightsStore[0][720]<=Wgt_0_720;WeightsStore[0][721]<=Wgt_0_721;WeightsStore[0][722]<=Wgt_0_722;WeightsStore[0][723]<=Wgt_0_723;WeightsStore[0][724]<=Wgt_0_724;WeightsStore[0][725]<=Wgt_0_725;WeightsStore[0][726]<=Wgt_0_726;WeightsStore[0][727]<=Wgt_0_727;WeightsStore[0][728]<=Wgt_0_728;WeightsStore[0][729]<=Wgt_0_729;WeightsStore[0][730]<=Wgt_0_730;WeightsStore[0][731]<=Wgt_0_731;WeightsStore[0][732]<=Wgt_0_732;WeightsStore[0][733]<=Wgt_0_733;WeightsStore[0][734]<=Wgt_0_734;WeightsStore[0][735]<=Wgt_0_735;WeightsStore[0][736]<=Wgt_0_736;WeightsStore[0][737]<=Wgt_0_737;WeightsStore[0][738]<=Wgt_0_738;WeightsStore[0][739]<=Wgt_0_739;WeightsStore[0][740]<=Wgt_0_740;WeightsStore[0][741]<=Wgt_0_741;WeightsStore[0][742]<=Wgt_0_742;WeightsStore[0][743]<=Wgt_0_743;WeightsStore[0][744]<=Wgt_0_744;WeightsStore[0][745]<=Wgt_0_745;WeightsStore[0][746]<=Wgt_0_746;WeightsStore[0][747]<=Wgt_0_747;WeightsStore[0][748]<=Wgt_0_748;WeightsStore[0][749]<=Wgt_0_749;WeightsStore[0][750]<=Wgt_0_750;WeightsStore[0][751]<=Wgt_0_751;WeightsStore[0][752]<=Wgt_0_752;WeightsStore[0][753]<=Wgt_0_753;WeightsStore[0][754]<=Wgt_0_754;WeightsStore[0][755]<=Wgt_0_755;WeightsStore[0][756]<=Wgt_0_756;WeightsStore[0][757]<=Wgt_0_757;WeightsStore[0][758]<=Wgt_0_758;WeightsStore[0][759]<=Wgt_0_759;WeightsStore[0][760]<=Wgt_0_760;WeightsStore[0][761]<=Wgt_0_761;WeightsStore[0][762]<=Wgt_0_762;WeightsStore[0][763]<=Wgt_0_763;WeightsStore[0][764]<=Wgt_0_764;WeightsStore[0][765]<=Wgt_0_765;WeightsStore[0][766]<=Wgt_0_766;WeightsStore[0][767]<=Wgt_0_767;WeightsStore[0][768]<=Wgt_0_768;WeightsStore[0][769]<=Wgt_0_769;WeightsStore[0][770]<=Wgt_0_770;WeightsStore[0][771]<=Wgt_0_771;WeightsStore[0][772]<=Wgt_0_772;WeightsStore[0][773]<=Wgt_0_773;WeightsStore[0][774]<=Wgt_0_774;WeightsStore[0][775]<=Wgt_0_775;WeightsStore[0][776]<=Wgt_0_776;WeightsStore[0][777]<=Wgt_0_777;WeightsStore[0][778]<=Wgt_0_778;WeightsStore[0][779]<=Wgt_0_779;WeightsStore[0][780]<=Wgt_0_780;WeightsStore[0][781]<=Wgt_0_781;WeightsStore[0][782]<=Wgt_0_782;WeightsStore[0][783]<=Wgt_0_783;WeightsStore[0][784]<=Wgt_0_784;WeightsStore[1][0]<=Wgt_1_0;WeightsStore[1][1]<=Wgt_1_1;WeightsStore[1][2]<=Wgt_1_2;WeightsStore[1][3]<=Wgt_1_3;WeightsStore[1][4]<=Wgt_1_4;WeightsStore[1][5]<=Wgt_1_5;WeightsStore[1][6]<=Wgt_1_6;WeightsStore[1][7]<=Wgt_1_7;WeightsStore[1][8]<=Wgt_1_8;WeightsStore[1][9]<=Wgt_1_9;WeightsStore[1][10]<=Wgt_1_10;WeightsStore[1][11]<=Wgt_1_11;WeightsStore[1][12]<=Wgt_1_12;WeightsStore[1][13]<=Wgt_1_13;WeightsStore[1][14]<=Wgt_1_14;WeightsStore[1][15]<=Wgt_1_15;WeightsStore[1][16]<=Wgt_1_16;WeightsStore[1][17]<=Wgt_1_17;WeightsStore[1][18]<=Wgt_1_18;WeightsStore[1][19]<=Wgt_1_19;WeightsStore[1][20]<=Wgt_1_20;WeightsStore[1][21]<=Wgt_1_21;WeightsStore[1][22]<=Wgt_1_22;WeightsStore[1][23]<=Wgt_1_23;WeightsStore[1][24]<=Wgt_1_24;WeightsStore[1][25]<=Wgt_1_25;WeightsStore[1][26]<=Wgt_1_26;WeightsStore[1][27]<=Wgt_1_27;WeightsStore[1][28]<=Wgt_1_28;WeightsStore[1][29]<=Wgt_1_29;WeightsStore[1][30]<=Wgt_1_30;WeightsStore[1][31]<=Wgt_1_31;WeightsStore[1][32]<=Wgt_1_32;WeightsStore[1][33]<=Wgt_1_33;WeightsStore[1][34]<=Wgt_1_34;WeightsStore[1][35]<=Wgt_1_35;WeightsStore[1][36]<=Wgt_1_36;WeightsStore[1][37]<=Wgt_1_37;WeightsStore[1][38]<=Wgt_1_38;WeightsStore[1][39]<=Wgt_1_39;WeightsStore[1][40]<=Wgt_1_40;WeightsStore[1][41]<=Wgt_1_41;WeightsStore[1][42]<=Wgt_1_42;WeightsStore[1][43]<=Wgt_1_43;WeightsStore[1][44]<=Wgt_1_44;WeightsStore[1][45]<=Wgt_1_45;WeightsStore[1][46]<=Wgt_1_46;WeightsStore[1][47]<=Wgt_1_47;WeightsStore[1][48]<=Wgt_1_48;WeightsStore[1][49]<=Wgt_1_49;WeightsStore[1][50]<=Wgt_1_50;WeightsStore[1][51]<=Wgt_1_51;WeightsStore[1][52]<=Wgt_1_52;WeightsStore[1][53]<=Wgt_1_53;WeightsStore[1][54]<=Wgt_1_54;WeightsStore[1][55]<=Wgt_1_55;WeightsStore[1][56]<=Wgt_1_56;WeightsStore[1][57]<=Wgt_1_57;WeightsStore[1][58]<=Wgt_1_58;WeightsStore[1][59]<=Wgt_1_59;WeightsStore[1][60]<=Wgt_1_60;WeightsStore[1][61]<=Wgt_1_61;WeightsStore[1][62]<=Wgt_1_62;WeightsStore[1][63]<=Wgt_1_63;WeightsStore[1][64]<=Wgt_1_64;WeightsStore[1][65]<=Wgt_1_65;WeightsStore[1][66]<=Wgt_1_66;WeightsStore[1][67]<=Wgt_1_67;WeightsStore[1][68]<=Wgt_1_68;WeightsStore[1][69]<=Wgt_1_69;WeightsStore[1][70]<=Wgt_1_70;WeightsStore[1][71]<=Wgt_1_71;WeightsStore[1][72]<=Wgt_1_72;WeightsStore[1][73]<=Wgt_1_73;WeightsStore[1][74]<=Wgt_1_74;WeightsStore[1][75]<=Wgt_1_75;WeightsStore[1][76]<=Wgt_1_76;WeightsStore[1][77]<=Wgt_1_77;WeightsStore[1][78]<=Wgt_1_78;WeightsStore[1][79]<=Wgt_1_79;WeightsStore[1][80]<=Wgt_1_80;WeightsStore[1][81]<=Wgt_1_81;WeightsStore[1][82]<=Wgt_1_82;WeightsStore[1][83]<=Wgt_1_83;WeightsStore[1][84]<=Wgt_1_84;WeightsStore[1][85]<=Wgt_1_85;WeightsStore[1][86]<=Wgt_1_86;WeightsStore[1][87]<=Wgt_1_87;WeightsStore[1][88]<=Wgt_1_88;WeightsStore[1][89]<=Wgt_1_89;WeightsStore[1][90]<=Wgt_1_90;WeightsStore[1][91]<=Wgt_1_91;WeightsStore[1][92]<=Wgt_1_92;WeightsStore[1][93]<=Wgt_1_93;WeightsStore[1][94]<=Wgt_1_94;WeightsStore[1][95]<=Wgt_1_95;WeightsStore[1][96]<=Wgt_1_96;WeightsStore[1][97]<=Wgt_1_97;WeightsStore[1][98]<=Wgt_1_98;WeightsStore[1][99]<=Wgt_1_99;WeightsStore[1][100]<=Wgt_1_100;WeightsStore[1][101]<=Wgt_1_101;WeightsStore[1][102]<=Wgt_1_102;WeightsStore[1][103]<=Wgt_1_103;WeightsStore[1][104]<=Wgt_1_104;WeightsStore[1][105]<=Wgt_1_105;WeightsStore[1][106]<=Wgt_1_106;WeightsStore[1][107]<=Wgt_1_107;WeightsStore[1][108]<=Wgt_1_108;WeightsStore[1][109]<=Wgt_1_109;WeightsStore[1][110]<=Wgt_1_110;WeightsStore[1][111]<=Wgt_1_111;WeightsStore[1][112]<=Wgt_1_112;WeightsStore[1][113]<=Wgt_1_113;WeightsStore[1][114]<=Wgt_1_114;WeightsStore[1][115]<=Wgt_1_115;WeightsStore[1][116]<=Wgt_1_116;WeightsStore[1][117]<=Wgt_1_117;WeightsStore[1][118]<=Wgt_1_118;WeightsStore[1][119]<=Wgt_1_119;WeightsStore[1][120]<=Wgt_1_120;WeightsStore[1][121]<=Wgt_1_121;WeightsStore[1][122]<=Wgt_1_122;WeightsStore[1][123]<=Wgt_1_123;WeightsStore[1][124]<=Wgt_1_124;WeightsStore[1][125]<=Wgt_1_125;WeightsStore[1][126]<=Wgt_1_126;WeightsStore[1][127]<=Wgt_1_127;WeightsStore[1][128]<=Wgt_1_128;WeightsStore[1][129]<=Wgt_1_129;WeightsStore[1][130]<=Wgt_1_130;WeightsStore[1][131]<=Wgt_1_131;WeightsStore[1][132]<=Wgt_1_132;WeightsStore[1][133]<=Wgt_1_133;WeightsStore[1][134]<=Wgt_1_134;WeightsStore[1][135]<=Wgt_1_135;WeightsStore[1][136]<=Wgt_1_136;WeightsStore[1][137]<=Wgt_1_137;WeightsStore[1][138]<=Wgt_1_138;WeightsStore[1][139]<=Wgt_1_139;WeightsStore[1][140]<=Wgt_1_140;WeightsStore[1][141]<=Wgt_1_141;WeightsStore[1][142]<=Wgt_1_142;WeightsStore[1][143]<=Wgt_1_143;WeightsStore[1][144]<=Wgt_1_144;WeightsStore[1][145]<=Wgt_1_145;WeightsStore[1][146]<=Wgt_1_146;WeightsStore[1][147]<=Wgt_1_147;WeightsStore[1][148]<=Wgt_1_148;WeightsStore[1][149]<=Wgt_1_149;WeightsStore[1][150]<=Wgt_1_150;WeightsStore[1][151]<=Wgt_1_151;WeightsStore[1][152]<=Wgt_1_152;WeightsStore[1][153]<=Wgt_1_153;WeightsStore[1][154]<=Wgt_1_154;WeightsStore[1][155]<=Wgt_1_155;WeightsStore[1][156]<=Wgt_1_156;WeightsStore[1][157]<=Wgt_1_157;WeightsStore[1][158]<=Wgt_1_158;WeightsStore[1][159]<=Wgt_1_159;WeightsStore[1][160]<=Wgt_1_160;WeightsStore[1][161]<=Wgt_1_161;WeightsStore[1][162]<=Wgt_1_162;WeightsStore[1][163]<=Wgt_1_163;WeightsStore[1][164]<=Wgt_1_164;WeightsStore[1][165]<=Wgt_1_165;WeightsStore[1][166]<=Wgt_1_166;WeightsStore[1][167]<=Wgt_1_167;WeightsStore[1][168]<=Wgt_1_168;WeightsStore[1][169]<=Wgt_1_169;WeightsStore[1][170]<=Wgt_1_170;WeightsStore[1][171]<=Wgt_1_171;WeightsStore[1][172]<=Wgt_1_172;WeightsStore[1][173]<=Wgt_1_173;WeightsStore[1][174]<=Wgt_1_174;WeightsStore[1][175]<=Wgt_1_175;WeightsStore[1][176]<=Wgt_1_176;WeightsStore[1][177]<=Wgt_1_177;WeightsStore[1][178]<=Wgt_1_178;WeightsStore[1][179]<=Wgt_1_179;WeightsStore[1][180]<=Wgt_1_180;WeightsStore[1][181]<=Wgt_1_181;WeightsStore[1][182]<=Wgt_1_182;WeightsStore[1][183]<=Wgt_1_183;WeightsStore[1][184]<=Wgt_1_184;WeightsStore[1][185]<=Wgt_1_185;WeightsStore[1][186]<=Wgt_1_186;WeightsStore[1][187]<=Wgt_1_187;WeightsStore[1][188]<=Wgt_1_188;WeightsStore[1][189]<=Wgt_1_189;WeightsStore[1][190]<=Wgt_1_190;WeightsStore[1][191]<=Wgt_1_191;WeightsStore[1][192]<=Wgt_1_192;WeightsStore[1][193]<=Wgt_1_193;WeightsStore[1][194]<=Wgt_1_194;WeightsStore[1][195]<=Wgt_1_195;WeightsStore[1][196]<=Wgt_1_196;WeightsStore[1][197]<=Wgt_1_197;WeightsStore[1][198]<=Wgt_1_198;WeightsStore[1][199]<=Wgt_1_199;WeightsStore[1][200]<=Wgt_1_200;WeightsStore[1][201]<=Wgt_1_201;WeightsStore[1][202]<=Wgt_1_202;WeightsStore[1][203]<=Wgt_1_203;WeightsStore[1][204]<=Wgt_1_204;WeightsStore[1][205]<=Wgt_1_205;WeightsStore[1][206]<=Wgt_1_206;WeightsStore[1][207]<=Wgt_1_207;WeightsStore[1][208]<=Wgt_1_208;WeightsStore[1][209]<=Wgt_1_209;WeightsStore[1][210]<=Wgt_1_210;WeightsStore[1][211]<=Wgt_1_211;WeightsStore[1][212]<=Wgt_1_212;WeightsStore[1][213]<=Wgt_1_213;WeightsStore[1][214]<=Wgt_1_214;WeightsStore[1][215]<=Wgt_1_215;WeightsStore[1][216]<=Wgt_1_216;WeightsStore[1][217]<=Wgt_1_217;WeightsStore[1][218]<=Wgt_1_218;WeightsStore[1][219]<=Wgt_1_219;WeightsStore[1][220]<=Wgt_1_220;WeightsStore[1][221]<=Wgt_1_221;WeightsStore[1][222]<=Wgt_1_222;WeightsStore[1][223]<=Wgt_1_223;WeightsStore[1][224]<=Wgt_1_224;WeightsStore[1][225]<=Wgt_1_225;WeightsStore[1][226]<=Wgt_1_226;WeightsStore[1][227]<=Wgt_1_227;WeightsStore[1][228]<=Wgt_1_228;WeightsStore[1][229]<=Wgt_1_229;WeightsStore[1][230]<=Wgt_1_230;WeightsStore[1][231]<=Wgt_1_231;WeightsStore[1][232]<=Wgt_1_232;WeightsStore[1][233]<=Wgt_1_233;WeightsStore[1][234]<=Wgt_1_234;WeightsStore[1][235]<=Wgt_1_235;WeightsStore[1][236]<=Wgt_1_236;WeightsStore[1][237]<=Wgt_1_237;WeightsStore[1][238]<=Wgt_1_238;WeightsStore[1][239]<=Wgt_1_239;WeightsStore[1][240]<=Wgt_1_240;WeightsStore[1][241]<=Wgt_1_241;WeightsStore[1][242]<=Wgt_1_242;WeightsStore[1][243]<=Wgt_1_243;WeightsStore[1][244]<=Wgt_1_244;WeightsStore[1][245]<=Wgt_1_245;WeightsStore[1][246]<=Wgt_1_246;WeightsStore[1][247]<=Wgt_1_247;WeightsStore[1][248]<=Wgt_1_248;WeightsStore[1][249]<=Wgt_1_249;WeightsStore[1][250]<=Wgt_1_250;WeightsStore[1][251]<=Wgt_1_251;WeightsStore[1][252]<=Wgt_1_252;WeightsStore[1][253]<=Wgt_1_253;WeightsStore[1][254]<=Wgt_1_254;WeightsStore[1][255]<=Wgt_1_255;WeightsStore[1][256]<=Wgt_1_256;WeightsStore[1][257]<=Wgt_1_257;WeightsStore[1][258]<=Wgt_1_258;WeightsStore[1][259]<=Wgt_1_259;WeightsStore[1][260]<=Wgt_1_260;WeightsStore[1][261]<=Wgt_1_261;WeightsStore[1][262]<=Wgt_1_262;WeightsStore[1][263]<=Wgt_1_263;WeightsStore[1][264]<=Wgt_1_264;WeightsStore[1][265]<=Wgt_1_265;WeightsStore[1][266]<=Wgt_1_266;WeightsStore[1][267]<=Wgt_1_267;WeightsStore[1][268]<=Wgt_1_268;WeightsStore[1][269]<=Wgt_1_269;WeightsStore[1][270]<=Wgt_1_270;WeightsStore[1][271]<=Wgt_1_271;WeightsStore[1][272]<=Wgt_1_272;WeightsStore[1][273]<=Wgt_1_273;WeightsStore[1][274]<=Wgt_1_274;WeightsStore[1][275]<=Wgt_1_275;WeightsStore[1][276]<=Wgt_1_276;WeightsStore[1][277]<=Wgt_1_277;WeightsStore[1][278]<=Wgt_1_278;WeightsStore[1][279]<=Wgt_1_279;WeightsStore[1][280]<=Wgt_1_280;WeightsStore[1][281]<=Wgt_1_281;WeightsStore[1][282]<=Wgt_1_282;WeightsStore[1][283]<=Wgt_1_283;WeightsStore[1][284]<=Wgt_1_284;WeightsStore[1][285]<=Wgt_1_285;WeightsStore[1][286]<=Wgt_1_286;WeightsStore[1][287]<=Wgt_1_287;WeightsStore[1][288]<=Wgt_1_288;WeightsStore[1][289]<=Wgt_1_289;WeightsStore[1][290]<=Wgt_1_290;WeightsStore[1][291]<=Wgt_1_291;WeightsStore[1][292]<=Wgt_1_292;WeightsStore[1][293]<=Wgt_1_293;WeightsStore[1][294]<=Wgt_1_294;WeightsStore[1][295]<=Wgt_1_295;WeightsStore[1][296]<=Wgt_1_296;WeightsStore[1][297]<=Wgt_1_297;WeightsStore[1][298]<=Wgt_1_298;WeightsStore[1][299]<=Wgt_1_299;WeightsStore[1][300]<=Wgt_1_300;WeightsStore[1][301]<=Wgt_1_301;WeightsStore[1][302]<=Wgt_1_302;WeightsStore[1][303]<=Wgt_1_303;WeightsStore[1][304]<=Wgt_1_304;WeightsStore[1][305]<=Wgt_1_305;WeightsStore[1][306]<=Wgt_1_306;WeightsStore[1][307]<=Wgt_1_307;WeightsStore[1][308]<=Wgt_1_308;WeightsStore[1][309]<=Wgt_1_309;WeightsStore[1][310]<=Wgt_1_310;WeightsStore[1][311]<=Wgt_1_311;WeightsStore[1][312]<=Wgt_1_312;WeightsStore[1][313]<=Wgt_1_313;WeightsStore[1][314]<=Wgt_1_314;WeightsStore[1][315]<=Wgt_1_315;WeightsStore[1][316]<=Wgt_1_316;WeightsStore[1][317]<=Wgt_1_317;WeightsStore[1][318]<=Wgt_1_318;WeightsStore[1][319]<=Wgt_1_319;WeightsStore[1][320]<=Wgt_1_320;WeightsStore[1][321]<=Wgt_1_321;WeightsStore[1][322]<=Wgt_1_322;WeightsStore[1][323]<=Wgt_1_323;WeightsStore[1][324]<=Wgt_1_324;WeightsStore[1][325]<=Wgt_1_325;WeightsStore[1][326]<=Wgt_1_326;WeightsStore[1][327]<=Wgt_1_327;WeightsStore[1][328]<=Wgt_1_328;WeightsStore[1][329]<=Wgt_1_329;WeightsStore[1][330]<=Wgt_1_330;WeightsStore[1][331]<=Wgt_1_331;WeightsStore[1][332]<=Wgt_1_332;WeightsStore[1][333]<=Wgt_1_333;WeightsStore[1][334]<=Wgt_1_334;WeightsStore[1][335]<=Wgt_1_335;WeightsStore[1][336]<=Wgt_1_336;WeightsStore[1][337]<=Wgt_1_337;WeightsStore[1][338]<=Wgt_1_338;WeightsStore[1][339]<=Wgt_1_339;WeightsStore[1][340]<=Wgt_1_340;WeightsStore[1][341]<=Wgt_1_341;WeightsStore[1][342]<=Wgt_1_342;WeightsStore[1][343]<=Wgt_1_343;WeightsStore[1][344]<=Wgt_1_344;WeightsStore[1][345]<=Wgt_1_345;WeightsStore[1][346]<=Wgt_1_346;WeightsStore[1][347]<=Wgt_1_347;WeightsStore[1][348]<=Wgt_1_348;WeightsStore[1][349]<=Wgt_1_349;WeightsStore[1][350]<=Wgt_1_350;WeightsStore[1][351]<=Wgt_1_351;WeightsStore[1][352]<=Wgt_1_352;WeightsStore[1][353]<=Wgt_1_353;WeightsStore[1][354]<=Wgt_1_354;WeightsStore[1][355]<=Wgt_1_355;WeightsStore[1][356]<=Wgt_1_356;WeightsStore[1][357]<=Wgt_1_357;WeightsStore[1][358]<=Wgt_1_358;WeightsStore[1][359]<=Wgt_1_359;WeightsStore[1][360]<=Wgt_1_360;WeightsStore[1][361]<=Wgt_1_361;WeightsStore[1][362]<=Wgt_1_362;WeightsStore[1][363]<=Wgt_1_363;WeightsStore[1][364]<=Wgt_1_364;WeightsStore[1][365]<=Wgt_1_365;WeightsStore[1][366]<=Wgt_1_366;WeightsStore[1][367]<=Wgt_1_367;WeightsStore[1][368]<=Wgt_1_368;WeightsStore[1][369]<=Wgt_1_369;WeightsStore[1][370]<=Wgt_1_370;WeightsStore[1][371]<=Wgt_1_371;WeightsStore[1][372]<=Wgt_1_372;WeightsStore[1][373]<=Wgt_1_373;WeightsStore[1][374]<=Wgt_1_374;WeightsStore[1][375]<=Wgt_1_375;WeightsStore[1][376]<=Wgt_1_376;WeightsStore[1][377]<=Wgt_1_377;WeightsStore[1][378]<=Wgt_1_378;WeightsStore[1][379]<=Wgt_1_379;WeightsStore[1][380]<=Wgt_1_380;WeightsStore[1][381]<=Wgt_1_381;WeightsStore[1][382]<=Wgt_1_382;WeightsStore[1][383]<=Wgt_1_383;WeightsStore[1][384]<=Wgt_1_384;WeightsStore[1][385]<=Wgt_1_385;WeightsStore[1][386]<=Wgt_1_386;WeightsStore[1][387]<=Wgt_1_387;WeightsStore[1][388]<=Wgt_1_388;WeightsStore[1][389]<=Wgt_1_389;WeightsStore[1][390]<=Wgt_1_390;WeightsStore[1][391]<=Wgt_1_391;WeightsStore[1][392]<=Wgt_1_392;WeightsStore[1][393]<=Wgt_1_393;WeightsStore[1][394]<=Wgt_1_394;WeightsStore[1][395]<=Wgt_1_395;WeightsStore[1][396]<=Wgt_1_396;WeightsStore[1][397]<=Wgt_1_397;WeightsStore[1][398]<=Wgt_1_398;WeightsStore[1][399]<=Wgt_1_399;WeightsStore[1][400]<=Wgt_1_400;WeightsStore[1][401]<=Wgt_1_401;WeightsStore[1][402]<=Wgt_1_402;WeightsStore[1][403]<=Wgt_1_403;WeightsStore[1][404]<=Wgt_1_404;WeightsStore[1][405]<=Wgt_1_405;WeightsStore[1][406]<=Wgt_1_406;WeightsStore[1][407]<=Wgt_1_407;WeightsStore[1][408]<=Wgt_1_408;WeightsStore[1][409]<=Wgt_1_409;WeightsStore[1][410]<=Wgt_1_410;WeightsStore[1][411]<=Wgt_1_411;WeightsStore[1][412]<=Wgt_1_412;WeightsStore[1][413]<=Wgt_1_413;WeightsStore[1][414]<=Wgt_1_414;WeightsStore[1][415]<=Wgt_1_415;WeightsStore[1][416]<=Wgt_1_416;WeightsStore[1][417]<=Wgt_1_417;WeightsStore[1][418]<=Wgt_1_418;WeightsStore[1][419]<=Wgt_1_419;WeightsStore[1][420]<=Wgt_1_420;WeightsStore[1][421]<=Wgt_1_421;WeightsStore[1][422]<=Wgt_1_422;WeightsStore[1][423]<=Wgt_1_423;WeightsStore[1][424]<=Wgt_1_424;WeightsStore[1][425]<=Wgt_1_425;WeightsStore[1][426]<=Wgt_1_426;WeightsStore[1][427]<=Wgt_1_427;WeightsStore[1][428]<=Wgt_1_428;WeightsStore[1][429]<=Wgt_1_429;WeightsStore[1][430]<=Wgt_1_430;WeightsStore[1][431]<=Wgt_1_431;WeightsStore[1][432]<=Wgt_1_432;WeightsStore[1][433]<=Wgt_1_433;WeightsStore[1][434]<=Wgt_1_434;WeightsStore[1][435]<=Wgt_1_435;WeightsStore[1][436]<=Wgt_1_436;WeightsStore[1][437]<=Wgt_1_437;WeightsStore[1][438]<=Wgt_1_438;WeightsStore[1][439]<=Wgt_1_439;WeightsStore[1][440]<=Wgt_1_440;WeightsStore[1][441]<=Wgt_1_441;WeightsStore[1][442]<=Wgt_1_442;WeightsStore[1][443]<=Wgt_1_443;WeightsStore[1][444]<=Wgt_1_444;WeightsStore[1][445]<=Wgt_1_445;WeightsStore[1][446]<=Wgt_1_446;WeightsStore[1][447]<=Wgt_1_447;WeightsStore[1][448]<=Wgt_1_448;WeightsStore[1][449]<=Wgt_1_449;WeightsStore[1][450]<=Wgt_1_450;WeightsStore[1][451]<=Wgt_1_451;WeightsStore[1][452]<=Wgt_1_452;WeightsStore[1][453]<=Wgt_1_453;WeightsStore[1][454]<=Wgt_1_454;WeightsStore[1][455]<=Wgt_1_455;WeightsStore[1][456]<=Wgt_1_456;WeightsStore[1][457]<=Wgt_1_457;WeightsStore[1][458]<=Wgt_1_458;WeightsStore[1][459]<=Wgt_1_459;WeightsStore[1][460]<=Wgt_1_460;WeightsStore[1][461]<=Wgt_1_461;WeightsStore[1][462]<=Wgt_1_462;WeightsStore[1][463]<=Wgt_1_463;WeightsStore[1][464]<=Wgt_1_464;WeightsStore[1][465]<=Wgt_1_465;WeightsStore[1][466]<=Wgt_1_466;WeightsStore[1][467]<=Wgt_1_467;WeightsStore[1][468]<=Wgt_1_468;WeightsStore[1][469]<=Wgt_1_469;WeightsStore[1][470]<=Wgt_1_470;WeightsStore[1][471]<=Wgt_1_471;WeightsStore[1][472]<=Wgt_1_472;WeightsStore[1][473]<=Wgt_1_473;WeightsStore[1][474]<=Wgt_1_474;WeightsStore[1][475]<=Wgt_1_475;WeightsStore[1][476]<=Wgt_1_476;WeightsStore[1][477]<=Wgt_1_477;WeightsStore[1][478]<=Wgt_1_478;WeightsStore[1][479]<=Wgt_1_479;WeightsStore[1][480]<=Wgt_1_480;WeightsStore[1][481]<=Wgt_1_481;WeightsStore[1][482]<=Wgt_1_482;WeightsStore[1][483]<=Wgt_1_483;WeightsStore[1][484]<=Wgt_1_484;WeightsStore[1][485]<=Wgt_1_485;WeightsStore[1][486]<=Wgt_1_486;WeightsStore[1][487]<=Wgt_1_487;WeightsStore[1][488]<=Wgt_1_488;WeightsStore[1][489]<=Wgt_1_489;WeightsStore[1][490]<=Wgt_1_490;WeightsStore[1][491]<=Wgt_1_491;WeightsStore[1][492]<=Wgt_1_492;WeightsStore[1][493]<=Wgt_1_493;WeightsStore[1][494]<=Wgt_1_494;WeightsStore[1][495]<=Wgt_1_495;WeightsStore[1][496]<=Wgt_1_496;WeightsStore[1][497]<=Wgt_1_497;WeightsStore[1][498]<=Wgt_1_498;WeightsStore[1][499]<=Wgt_1_499;WeightsStore[1][500]<=Wgt_1_500;WeightsStore[1][501]<=Wgt_1_501;WeightsStore[1][502]<=Wgt_1_502;WeightsStore[1][503]<=Wgt_1_503;WeightsStore[1][504]<=Wgt_1_504;WeightsStore[1][505]<=Wgt_1_505;WeightsStore[1][506]<=Wgt_1_506;WeightsStore[1][507]<=Wgt_1_507;WeightsStore[1][508]<=Wgt_1_508;WeightsStore[1][509]<=Wgt_1_509;WeightsStore[1][510]<=Wgt_1_510;WeightsStore[1][511]<=Wgt_1_511;WeightsStore[1][512]<=Wgt_1_512;WeightsStore[1][513]<=Wgt_1_513;WeightsStore[1][514]<=Wgt_1_514;WeightsStore[1][515]<=Wgt_1_515;WeightsStore[1][516]<=Wgt_1_516;WeightsStore[1][517]<=Wgt_1_517;WeightsStore[1][518]<=Wgt_1_518;WeightsStore[1][519]<=Wgt_1_519;WeightsStore[1][520]<=Wgt_1_520;WeightsStore[1][521]<=Wgt_1_521;WeightsStore[1][522]<=Wgt_1_522;WeightsStore[1][523]<=Wgt_1_523;WeightsStore[1][524]<=Wgt_1_524;WeightsStore[1][525]<=Wgt_1_525;WeightsStore[1][526]<=Wgt_1_526;WeightsStore[1][527]<=Wgt_1_527;WeightsStore[1][528]<=Wgt_1_528;WeightsStore[1][529]<=Wgt_1_529;WeightsStore[1][530]<=Wgt_1_530;WeightsStore[1][531]<=Wgt_1_531;WeightsStore[1][532]<=Wgt_1_532;WeightsStore[1][533]<=Wgt_1_533;WeightsStore[1][534]<=Wgt_1_534;WeightsStore[1][535]<=Wgt_1_535;WeightsStore[1][536]<=Wgt_1_536;WeightsStore[1][537]<=Wgt_1_537;WeightsStore[1][538]<=Wgt_1_538;WeightsStore[1][539]<=Wgt_1_539;WeightsStore[1][540]<=Wgt_1_540;WeightsStore[1][541]<=Wgt_1_541;WeightsStore[1][542]<=Wgt_1_542;WeightsStore[1][543]<=Wgt_1_543;WeightsStore[1][544]<=Wgt_1_544;WeightsStore[1][545]<=Wgt_1_545;WeightsStore[1][546]<=Wgt_1_546;WeightsStore[1][547]<=Wgt_1_547;WeightsStore[1][548]<=Wgt_1_548;WeightsStore[1][549]<=Wgt_1_549;WeightsStore[1][550]<=Wgt_1_550;WeightsStore[1][551]<=Wgt_1_551;WeightsStore[1][552]<=Wgt_1_552;WeightsStore[1][553]<=Wgt_1_553;WeightsStore[1][554]<=Wgt_1_554;WeightsStore[1][555]<=Wgt_1_555;WeightsStore[1][556]<=Wgt_1_556;WeightsStore[1][557]<=Wgt_1_557;WeightsStore[1][558]<=Wgt_1_558;WeightsStore[1][559]<=Wgt_1_559;WeightsStore[1][560]<=Wgt_1_560;WeightsStore[1][561]<=Wgt_1_561;WeightsStore[1][562]<=Wgt_1_562;WeightsStore[1][563]<=Wgt_1_563;WeightsStore[1][564]<=Wgt_1_564;WeightsStore[1][565]<=Wgt_1_565;WeightsStore[1][566]<=Wgt_1_566;WeightsStore[1][567]<=Wgt_1_567;WeightsStore[1][568]<=Wgt_1_568;WeightsStore[1][569]<=Wgt_1_569;WeightsStore[1][570]<=Wgt_1_570;WeightsStore[1][571]<=Wgt_1_571;WeightsStore[1][572]<=Wgt_1_572;WeightsStore[1][573]<=Wgt_1_573;WeightsStore[1][574]<=Wgt_1_574;WeightsStore[1][575]<=Wgt_1_575;WeightsStore[1][576]<=Wgt_1_576;WeightsStore[1][577]<=Wgt_1_577;WeightsStore[1][578]<=Wgt_1_578;WeightsStore[1][579]<=Wgt_1_579;WeightsStore[1][580]<=Wgt_1_580;WeightsStore[1][581]<=Wgt_1_581;WeightsStore[1][582]<=Wgt_1_582;WeightsStore[1][583]<=Wgt_1_583;WeightsStore[1][584]<=Wgt_1_584;WeightsStore[1][585]<=Wgt_1_585;WeightsStore[1][586]<=Wgt_1_586;WeightsStore[1][587]<=Wgt_1_587;WeightsStore[1][588]<=Wgt_1_588;WeightsStore[1][589]<=Wgt_1_589;WeightsStore[1][590]<=Wgt_1_590;WeightsStore[1][591]<=Wgt_1_591;WeightsStore[1][592]<=Wgt_1_592;WeightsStore[1][593]<=Wgt_1_593;WeightsStore[1][594]<=Wgt_1_594;WeightsStore[1][595]<=Wgt_1_595;WeightsStore[1][596]<=Wgt_1_596;WeightsStore[1][597]<=Wgt_1_597;WeightsStore[1][598]<=Wgt_1_598;WeightsStore[1][599]<=Wgt_1_599;WeightsStore[1][600]<=Wgt_1_600;WeightsStore[1][601]<=Wgt_1_601;WeightsStore[1][602]<=Wgt_1_602;WeightsStore[1][603]<=Wgt_1_603;WeightsStore[1][604]<=Wgt_1_604;WeightsStore[1][605]<=Wgt_1_605;WeightsStore[1][606]<=Wgt_1_606;WeightsStore[1][607]<=Wgt_1_607;WeightsStore[1][608]<=Wgt_1_608;WeightsStore[1][609]<=Wgt_1_609;WeightsStore[1][610]<=Wgt_1_610;WeightsStore[1][611]<=Wgt_1_611;WeightsStore[1][612]<=Wgt_1_612;WeightsStore[1][613]<=Wgt_1_613;WeightsStore[1][614]<=Wgt_1_614;WeightsStore[1][615]<=Wgt_1_615;WeightsStore[1][616]<=Wgt_1_616;WeightsStore[1][617]<=Wgt_1_617;WeightsStore[1][618]<=Wgt_1_618;WeightsStore[1][619]<=Wgt_1_619;WeightsStore[1][620]<=Wgt_1_620;WeightsStore[1][621]<=Wgt_1_621;WeightsStore[1][622]<=Wgt_1_622;WeightsStore[1][623]<=Wgt_1_623;WeightsStore[1][624]<=Wgt_1_624;WeightsStore[1][625]<=Wgt_1_625;WeightsStore[1][626]<=Wgt_1_626;WeightsStore[1][627]<=Wgt_1_627;WeightsStore[1][628]<=Wgt_1_628;WeightsStore[1][629]<=Wgt_1_629;WeightsStore[1][630]<=Wgt_1_630;WeightsStore[1][631]<=Wgt_1_631;WeightsStore[1][632]<=Wgt_1_632;WeightsStore[1][633]<=Wgt_1_633;WeightsStore[1][634]<=Wgt_1_634;WeightsStore[1][635]<=Wgt_1_635;WeightsStore[1][636]<=Wgt_1_636;WeightsStore[1][637]<=Wgt_1_637;WeightsStore[1][638]<=Wgt_1_638;WeightsStore[1][639]<=Wgt_1_639;WeightsStore[1][640]<=Wgt_1_640;WeightsStore[1][641]<=Wgt_1_641;WeightsStore[1][642]<=Wgt_1_642;WeightsStore[1][643]<=Wgt_1_643;WeightsStore[1][644]<=Wgt_1_644;WeightsStore[1][645]<=Wgt_1_645;WeightsStore[1][646]<=Wgt_1_646;WeightsStore[1][647]<=Wgt_1_647;WeightsStore[1][648]<=Wgt_1_648;WeightsStore[1][649]<=Wgt_1_649;WeightsStore[1][650]<=Wgt_1_650;WeightsStore[1][651]<=Wgt_1_651;WeightsStore[1][652]<=Wgt_1_652;WeightsStore[1][653]<=Wgt_1_653;WeightsStore[1][654]<=Wgt_1_654;WeightsStore[1][655]<=Wgt_1_655;WeightsStore[1][656]<=Wgt_1_656;WeightsStore[1][657]<=Wgt_1_657;WeightsStore[1][658]<=Wgt_1_658;WeightsStore[1][659]<=Wgt_1_659;WeightsStore[1][660]<=Wgt_1_660;WeightsStore[1][661]<=Wgt_1_661;WeightsStore[1][662]<=Wgt_1_662;WeightsStore[1][663]<=Wgt_1_663;WeightsStore[1][664]<=Wgt_1_664;WeightsStore[1][665]<=Wgt_1_665;WeightsStore[1][666]<=Wgt_1_666;WeightsStore[1][667]<=Wgt_1_667;WeightsStore[1][668]<=Wgt_1_668;WeightsStore[1][669]<=Wgt_1_669;WeightsStore[1][670]<=Wgt_1_670;WeightsStore[1][671]<=Wgt_1_671;WeightsStore[1][672]<=Wgt_1_672;WeightsStore[1][673]<=Wgt_1_673;WeightsStore[1][674]<=Wgt_1_674;WeightsStore[1][675]<=Wgt_1_675;WeightsStore[1][676]<=Wgt_1_676;WeightsStore[1][677]<=Wgt_1_677;WeightsStore[1][678]<=Wgt_1_678;WeightsStore[1][679]<=Wgt_1_679;WeightsStore[1][680]<=Wgt_1_680;WeightsStore[1][681]<=Wgt_1_681;WeightsStore[1][682]<=Wgt_1_682;WeightsStore[1][683]<=Wgt_1_683;WeightsStore[1][684]<=Wgt_1_684;WeightsStore[1][685]<=Wgt_1_685;WeightsStore[1][686]<=Wgt_1_686;WeightsStore[1][687]<=Wgt_1_687;WeightsStore[1][688]<=Wgt_1_688;WeightsStore[1][689]<=Wgt_1_689;WeightsStore[1][690]<=Wgt_1_690;WeightsStore[1][691]<=Wgt_1_691;WeightsStore[1][692]<=Wgt_1_692;WeightsStore[1][693]<=Wgt_1_693;WeightsStore[1][694]<=Wgt_1_694;WeightsStore[1][695]<=Wgt_1_695;WeightsStore[1][696]<=Wgt_1_696;WeightsStore[1][697]<=Wgt_1_697;WeightsStore[1][698]<=Wgt_1_698;WeightsStore[1][699]<=Wgt_1_699;WeightsStore[1][700]<=Wgt_1_700;WeightsStore[1][701]<=Wgt_1_701;WeightsStore[1][702]<=Wgt_1_702;WeightsStore[1][703]<=Wgt_1_703;WeightsStore[1][704]<=Wgt_1_704;WeightsStore[1][705]<=Wgt_1_705;WeightsStore[1][706]<=Wgt_1_706;WeightsStore[1][707]<=Wgt_1_707;WeightsStore[1][708]<=Wgt_1_708;WeightsStore[1][709]<=Wgt_1_709;WeightsStore[1][710]<=Wgt_1_710;WeightsStore[1][711]<=Wgt_1_711;WeightsStore[1][712]<=Wgt_1_712;WeightsStore[1][713]<=Wgt_1_713;WeightsStore[1][714]<=Wgt_1_714;WeightsStore[1][715]<=Wgt_1_715;WeightsStore[1][716]<=Wgt_1_716;WeightsStore[1][717]<=Wgt_1_717;WeightsStore[1][718]<=Wgt_1_718;WeightsStore[1][719]<=Wgt_1_719;WeightsStore[1][720]<=Wgt_1_720;WeightsStore[1][721]<=Wgt_1_721;WeightsStore[1][722]<=Wgt_1_722;WeightsStore[1][723]<=Wgt_1_723;WeightsStore[1][724]<=Wgt_1_724;WeightsStore[1][725]<=Wgt_1_725;WeightsStore[1][726]<=Wgt_1_726;WeightsStore[1][727]<=Wgt_1_727;WeightsStore[1][728]<=Wgt_1_728;WeightsStore[1][729]<=Wgt_1_729;WeightsStore[1][730]<=Wgt_1_730;WeightsStore[1][731]<=Wgt_1_731;WeightsStore[1][732]<=Wgt_1_732;WeightsStore[1][733]<=Wgt_1_733;WeightsStore[1][734]<=Wgt_1_734;WeightsStore[1][735]<=Wgt_1_735;WeightsStore[1][736]<=Wgt_1_736;WeightsStore[1][737]<=Wgt_1_737;WeightsStore[1][738]<=Wgt_1_738;WeightsStore[1][739]<=Wgt_1_739;WeightsStore[1][740]<=Wgt_1_740;WeightsStore[1][741]<=Wgt_1_741;WeightsStore[1][742]<=Wgt_1_742;WeightsStore[1][743]<=Wgt_1_743;WeightsStore[1][744]<=Wgt_1_744;WeightsStore[1][745]<=Wgt_1_745;WeightsStore[1][746]<=Wgt_1_746;WeightsStore[1][747]<=Wgt_1_747;WeightsStore[1][748]<=Wgt_1_748;WeightsStore[1][749]<=Wgt_1_749;WeightsStore[1][750]<=Wgt_1_750;WeightsStore[1][751]<=Wgt_1_751;WeightsStore[1][752]<=Wgt_1_752;WeightsStore[1][753]<=Wgt_1_753;WeightsStore[1][754]<=Wgt_1_754;WeightsStore[1][755]<=Wgt_1_755;WeightsStore[1][756]<=Wgt_1_756;WeightsStore[1][757]<=Wgt_1_757;WeightsStore[1][758]<=Wgt_1_758;WeightsStore[1][759]<=Wgt_1_759;WeightsStore[1][760]<=Wgt_1_760;WeightsStore[1][761]<=Wgt_1_761;WeightsStore[1][762]<=Wgt_1_762;WeightsStore[1][763]<=Wgt_1_763;WeightsStore[1][764]<=Wgt_1_764;WeightsStore[1][765]<=Wgt_1_765;WeightsStore[1][766]<=Wgt_1_766;WeightsStore[1][767]<=Wgt_1_767;WeightsStore[1][768]<=Wgt_1_768;WeightsStore[1][769]<=Wgt_1_769;WeightsStore[1][770]<=Wgt_1_770;WeightsStore[1][771]<=Wgt_1_771;WeightsStore[1][772]<=Wgt_1_772;WeightsStore[1][773]<=Wgt_1_773;WeightsStore[1][774]<=Wgt_1_774;WeightsStore[1][775]<=Wgt_1_775;WeightsStore[1][776]<=Wgt_1_776;WeightsStore[1][777]<=Wgt_1_777;WeightsStore[1][778]<=Wgt_1_778;WeightsStore[1][779]<=Wgt_1_779;WeightsStore[1][780]<=Wgt_1_780;WeightsStore[1][781]<=Wgt_1_781;WeightsStore[1][782]<=Wgt_1_782;WeightsStore[1][783]<=Wgt_1_783;WeightsStore[1][784]<=Wgt_1_784;WeightsStore[2][0]<=Wgt_2_0;WeightsStore[2][1]<=Wgt_2_1;WeightsStore[2][2]<=Wgt_2_2;WeightsStore[2][3]<=Wgt_2_3;WeightsStore[2][4]<=Wgt_2_4;WeightsStore[2][5]<=Wgt_2_5;WeightsStore[2][6]<=Wgt_2_6;WeightsStore[2][7]<=Wgt_2_7;WeightsStore[2][8]<=Wgt_2_8;WeightsStore[2][9]<=Wgt_2_9;WeightsStore[2][10]<=Wgt_2_10;WeightsStore[2][11]<=Wgt_2_11;WeightsStore[2][12]<=Wgt_2_12;WeightsStore[2][13]<=Wgt_2_13;WeightsStore[2][14]<=Wgt_2_14;WeightsStore[2][15]<=Wgt_2_15;WeightsStore[2][16]<=Wgt_2_16;WeightsStore[2][17]<=Wgt_2_17;WeightsStore[2][18]<=Wgt_2_18;WeightsStore[2][19]<=Wgt_2_19;WeightsStore[2][20]<=Wgt_2_20;WeightsStore[2][21]<=Wgt_2_21;WeightsStore[2][22]<=Wgt_2_22;WeightsStore[2][23]<=Wgt_2_23;WeightsStore[2][24]<=Wgt_2_24;WeightsStore[2][25]<=Wgt_2_25;WeightsStore[2][26]<=Wgt_2_26;WeightsStore[2][27]<=Wgt_2_27;WeightsStore[2][28]<=Wgt_2_28;WeightsStore[2][29]<=Wgt_2_29;WeightsStore[2][30]<=Wgt_2_30;WeightsStore[2][31]<=Wgt_2_31;WeightsStore[2][32]<=Wgt_2_32;WeightsStore[2][33]<=Wgt_2_33;WeightsStore[2][34]<=Wgt_2_34;WeightsStore[2][35]<=Wgt_2_35;WeightsStore[2][36]<=Wgt_2_36;WeightsStore[2][37]<=Wgt_2_37;WeightsStore[2][38]<=Wgt_2_38;WeightsStore[2][39]<=Wgt_2_39;WeightsStore[2][40]<=Wgt_2_40;WeightsStore[2][41]<=Wgt_2_41;WeightsStore[2][42]<=Wgt_2_42;WeightsStore[2][43]<=Wgt_2_43;WeightsStore[2][44]<=Wgt_2_44;WeightsStore[2][45]<=Wgt_2_45;WeightsStore[2][46]<=Wgt_2_46;WeightsStore[2][47]<=Wgt_2_47;WeightsStore[2][48]<=Wgt_2_48;WeightsStore[2][49]<=Wgt_2_49;WeightsStore[2][50]<=Wgt_2_50;WeightsStore[2][51]<=Wgt_2_51;WeightsStore[2][52]<=Wgt_2_52;WeightsStore[2][53]<=Wgt_2_53;WeightsStore[2][54]<=Wgt_2_54;WeightsStore[2][55]<=Wgt_2_55;WeightsStore[2][56]<=Wgt_2_56;WeightsStore[2][57]<=Wgt_2_57;WeightsStore[2][58]<=Wgt_2_58;WeightsStore[2][59]<=Wgt_2_59;WeightsStore[2][60]<=Wgt_2_60;WeightsStore[2][61]<=Wgt_2_61;WeightsStore[2][62]<=Wgt_2_62;WeightsStore[2][63]<=Wgt_2_63;WeightsStore[2][64]<=Wgt_2_64;WeightsStore[2][65]<=Wgt_2_65;WeightsStore[2][66]<=Wgt_2_66;WeightsStore[2][67]<=Wgt_2_67;WeightsStore[2][68]<=Wgt_2_68;WeightsStore[2][69]<=Wgt_2_69;WeightsStore[2][70]<=Wgt_2_70;WeightsStore[2][71]<=Wgt_2_71;WeightsStore[2][72]<=Wgt_2_72;WeightsStore[2][73]<=Wgt_2_73;WeightsStore[2][74]<=Wgt_2_74;WeightsStore[2][75]<=Wgt_2_75;WeightsStore[2][76]<=Wgt_2_76;WeightsStore[2][77]<=Wgt_2_77;WeightsStore[2][78]<=Wgt_2_78;WeightsStore[2][79]<=Wgt_2_79;WeightsStore[2][80]<=Wgt_2_80;WeightsStore[2][81]<=Wgt_2_81;WeightsStore[2][82]<=Wgt_2_82;WeightsStore[2][83]<=Wgt_2_83;WeightsStore[2][84]<=Wgt_2_84;WeightsStore[2][85]<=Wgt_2_85;WeightsStore[2][86]<=Wgt_2_86;WeightsStore[2][87]<=Wgt_2_87;WeightsStore[2][88]<=Wgt_2_88;WeightsStore[2][89]<=Wgt_2_89;WeightsStore[2][90]<=Wgt_2_90;WeightsStore[2][91]<=Wgt_2_91;WeightsStore[2][92]<=Wgt_2_92;WeightsStore[2][93]<=Wgt_2_93;WeightsStore[2][94]<=Wgt_2_94;WeightsStore[2][95]<=Wgt_2_95;WeightsStore[2][96]<=Wgt_2_96;WeightsStore[2][97]<=Wgt_2_97;WeightsStore[2][98]<=Wgt_2_98;WeightsStore[2][99]<=Wgt_2_99;WeightsStore[2][100]<=Wgt_2_100;WeightsStore[2][101]<=Wgt_2_101;WeightsStore[2][102]<=Wgt_2_102;WeightsStore[2][103]<=Wgt_2_103;WeightsStore[2][104]<=Wgt_2_104;WeightsStore[2][105]<=Wgt_2_105;WeightsStore[2][106]<=Wgt_2_106;WeightsStore[2][107]<=Wgt_2_107;WeightsStore[2][108]<=Wgt_2_108;WeightsStore[2][109]<=Wgt_2_109;WeightsStore[2][110]<=Wgt_2_110;WeightsStore[2][111]<=Wgt_2_111;WeightsStore[2][112]<=Wgt_2_112;WeightsStore[2][113]<=Wgt_2_113;WeightsStore[2][114]<=Wgt_2_114;WeightsStore[2][115]<=Wgt_2_115;WeightsStore[2][116]<=Wgt_2_116;WeightsStore[2][117]<=Wgt_2_117;WeightsStore[2][118]<=Wgt_2_118;WeightsStore[2][119]<=Wgt_2_119;WeightsStore[2][120]<=Wgt_2_120;WeightsStore[2][121]<=Wgt_2_121;WeightsStore[2][122]<=Wgt_2_122;WeightsStore[2][123]<=Wgt_2_123;WeightsStore[2][124]<=Wgt_2_124;WeightsStore[2][125]<=Wgt_2_125;WeightsStore[2][126]<=Wgt_2_126;WeightsStore[2][127]<=Wgt_2_127;WeightsStore[2][128]<=Wgt_2_128;WeightsStore[2][129]<=Wgt_2_129;WeightsStore[2][130]<=Wgt_2_130;WeightsStore[2][131]<=Wgt_2_131;WeightsStore[2][132]<=Wgt_2_132;WeightsStore[2][133]<=Wgt_2_133;WeightsStore[2][134]<=Wgt_2_134;WeightsStore[2][135]<=Wgt_2_135;WeightsStore[2][136]<=Wgt_2_136;WeightsStore[2][137]<=Wgt_2_137;WeightsStore[2][138]<=Wgt_2_138;WeightsStore[2][139]<=Wgt_2_139;WeightsStore[2][140]<=Wgt_2_140;WeightsStore[2][141]<=Wgt_2_141;WeightsStore[2][142]<=Wgt_2_142;WeightsStore[2][143]<=Wgt_2_143;WeightsStore[2][144]<=Wgt_2_144;WeightsStore[2][145]<=Wgt_2_145;WeightsStore[2][146]<=Wgt_2_146;WeightsStore[2][147]<=Wgt_2_147;WeightsStore[2][148]<=Wgt_2_148;WeightsStore[2][149]<=Wgt_2_149;WeightsStore[2][150]<=Wgt_2_150;WeightsStore[2][151]<=Wgt_2_151;WeightsStore[2][152]<=Wgt_2_152;WeightsStore[2][153]<=Wgt_2_153;WeightsStore[2][154]<=Wgt_2_154;WeightsStore[2][155]<=Wgt_2_155;WeightsStore[2][156]<=Wgt_2_156;WeightsStore[2][157]<=Wgt_2_157;WeightsStore[2][158]<=Wgt_2_158;WeightsStore[2][159]<=Wgt_2_159;WeightsStore[2][160]<=Wgt_2_160;WeightsStore[2][161]<=Wgt_2_161;WeightsStore[2][162]<=Wgt_2_162;WeightsStore[2][163]<=Wgt_2_163;WeightsStore[2][164]<=Wgt_2_164;WeightsStore[2][165]<=Wgt_2_165;WeightsStore[2][166]<=Wgt_2_166;WeightsStore[2][167]<=Wgt_2_167;WeightsStore[2][168]<=Wgt_2_168;WeightsStore[2][169]<=Wgt_2_169;WeightsStore[2][170]<=Wgt_2_170;WeightsStore[2][171]<=Wgt_2_171;WeightsStore[2][172]<=Wgt_2_172;WeightsStore[2][173]<=Wgt_2_173;WeightsStore[2][174]<=Wgt_2_174;WeightsStore[2][175]<=Wgt_2_175;WeightsStore[2][176]<=Wgt_2_176;WeightsStore[2][177]<=Wgt_2_177;WeightsStore[2][178]<=Wgt_2_178;WeightsStore[2][179]<=Wgt_2_179;WeightsStore[2][180]<=Wgt_2_180;WeightsStore[2][181]<=Wgt_2_181;WeightsStore[2][182]<=Wgt_2_182;WeightsStore[2][183]<=Wgt_2_183;WeightsStore[2][184]<=Wgt_2_184;WeightsStore[2][185]<=Wgt_2_185;WeightsStore[2][186]<=Wgt_2_186;WeightsStore[2][187]<=Wgt_2_187;WeightsStore[2][188]<=Wgt_2_188;WeightsStore[2][189]<=Wgt_2_189;WeightsStore[2][190]<=Wgt_2_190;WeightsStore[2][191]<=Wgt_2_191;WeightsStore[2][192]<=Wgt_2_192;WeightsStore[2][193]<=Wgt_2_193;WeightsStore[2][194]<=Wgt_2_194;WeightsStore[2][195]<=Wgt_2_195;WeightsStore[2][196]<=Wgt_2_196;WeightsStore[2][197]<=Wgt_2_197;WeightsStore[2][198]<=Wgt_2_198;WeightsStore[2][199]<=Wgt_2_199;WeightsStore[2][200]<=Wgt_2_200;WeightsStore[2][201]<=Wgt_2_201;WeightsStore[2][202]<=Wgt_2_202;WeightsStore[2][203]<=Wgt_2_203;WeightsStore[2][204]<=Wgt_2_204;WeightsStore[2][205]<=Wgt_2_205;WeightsStore[2][206]<=Wgt_2_206;WeightsStore[2][207]<=Wgt_2_207;WeightsStore[2][208]<=Wgt_2_208;WeightsStore[2][209]<=Wgt_2_209;WeightsStore[2][210]<=Wgt_2_210;WeightsStore[2][211]<=Wgt_2_211;WeightsStore[2][212]<=Wgt_2_212;WeightsStore[2][213]<=Wgt_2_213;WeightsStore[2][214]<=Wgt_2_214;WeightsStore[2][215]<=Wgt_2_215;WeightsStore[2][216]<=Wgt_2_216;WeightsStore[2][217]<=Wgt_2_217;WeightsStore[2][218]<=Wgt_2_218;WeightsStore[2][219]<=Wgt_2_219;WeightsStore[2][220]<=Wgt_2_220;WeightsStore[2][221]<=Wgt_2_221;WeightsStore[2][222]<=Wgt_2_222;WeightsStore[2][223]<=Wgt_2_223;WeightsStore[2][224]<=Wgt_2_224;WeightsStore[2][225]<=Wgt_2_225;WeightsStore[2][226]<=Wgt_2_226;WeightsStore[2][227]<=Wgt_2_227;WeightsStore[2][228]<=Wgt_2_228;WeightsStore[2][229]<=Wgt_2_229;WeightsStore[2][230]<=Wgt_2_230;WeightsStore[2][231]<=Wgt_2_231;WeightsStore[2][232]<=Wgt_2_232;WeightsStore[2][233]<=Wgt_2_233;WeightsStore[2][234]<=Wgt_2_234;WeightsStore[2][235]<=Wgt_2_235;WeightsStore[2][236]<=Wgt_2_236;WeightsStore[2][237]<=Wgt_2_237;WeightsStore[2][238]<=Wgt_2_238;WeightsStore[2][239]<=Wgt_2_239;WeightsStore[2][240]<=Wgt_2_240;WeightsStore[2][241]<=Wgt_2_241;WeightsStore[2][242]<=Wgt_2_242;WeightsStore[2][243]<=Wgt_2_243;WeightsStore[2][244]<=Wgt_2_244;WeightsStore[2][245]<=Wgt_2_245;WeightsStore[2][246]<=Wgt_2_246;WeightsStore[2][247]<=Wgt_2_247;WeightsStore[2][248]<=Wgt_2_248;WeightsStore[2][249]<=Wgt_2_249;WeightsStore[2][250]<=Wgt_2_250;WeightsStore[2][251]<=Wgt_2_251;WeightsStore[2][252]<=Wgt_2_252;WeightsStore[2][253]<=Wgt_2_253;WeightsStore[2][254]<=Wgt_2_254;WeightsStore[2][255]<=Wgt_2_255;WeightsStore[2][256]<=Wgt_2_256;WeightsStore[2][257]<=Wgt_2_257;WeightsStore[2][258]<=Wgt_2_258;WeightsStore[2][259]<=Wgt_2_259;WeightsStore[2][260]<=Wgt_2_260;WeightsStore[2][261]<=Wgt_2_261;WeightsStore[2][262]<=Wgt_2_262;WeightsStore[2][263]<=Wgt_2_263;WeightsStore[2][264]<=Wgt_2_264;WeightsStore[2][265]<=Wgt_2_265;WeightsStore[2][266]<=Wgt_2_266;WeightsStore[2][267]<=Wgt_2_267;WeightsStore[2][268]<=Wgt_2_268;WeightsStore[2][269]<=Wgt_2_269;WeightsStore[2][270]<=Wgt_2_270;WeightsStore[2][271]<=Wgt_2_271;WeightsStore[2][272]<=Wgt_2_272;WeightsStore[2][273]<=Wgt_2_273;WeightsStore[2][274]<=Wgt_2_274;WeightsStore[2][275]<=Wgt_2_275;WeightsStore[2][276]<=Wgt_2_276;WeightsStore[2][277]<=Wgt_2_277;WeightsStore[2][278]<=Wgt_2_278;WeightsStore[2][279]<=Wgt_2_279;WeightsStore[2][280]<=Wgt_2_280;WeightsStore[2][281]<=Wgt_2_281;WeightsStore[2][282]<=Wgt_2_282;WeightsStore[2][283]<=Wgt_2_283;WeightsStore[2][284]<=Wgt_2_284;WeightsStore[2][285]<=Wgt_2_285;WeightsStore[2][286]<=Wgt_2_286;WeightsStore[2][287]<=Wgt_2_287;WeightsStore[2][288]<=Wgt_2_288;WeightsStore[2][289]<=Wgt_2_289;WeightsStore[2][290]<=Wgt_2_290;WeightsStore[2][291]<=Wgt_2_291;WeightsStore[2][292]<=Wgt_2_292;WeightsStore[2][293]<=Wgt_2_293;WeightsStore[2][294]<=Wgt_2_294;WeightsStore[2][295]<=Wgt_2_295;WeightsStore[2][296]<=Wgt_2_296;WeightsStore[2][297]<=Wgt_2_297;WeightsStore[2][298]<=Wgt_2_298;WeightsStore[2][299]<=Wgt_2_299;WeightsStore[2][300]<=Wgt_2_300;WeightsStore[2][301]<=Wgt_2_301;WeightsStore[2][302]<=Wgt_2_302;WeightsStore[2][303]<=Wgt_2_303;WeightsStore[2][304]<=Wgt_2_304;WeightsStore[2][305]<=Wgt_2_305;WeightsStore[2][306]<=Wgt_2_306;WeightsStore[2][307]<=Wgt_2_307;WeightsStore[2][308]<=Wgt_2_308;WeightsStore[2][309]<=Wgt_2_309;WeightsStore[2][310]<=Wgt_2_310;WeightsStore[2][311]<=Wgt_2_311;WeightsStore[2][312]<=Wgt_2_312;WeightsStore[2][313]<=Wgt_2_313;WeightsStore[2][314]<=Wgt_2_314;WeightsStore[2][315]<=Wgt_2_315;WeightsStore[2][316]<=Wgt_2_316;WeightsStore[2][317]<=Wgt_2_317;WeightsStore[2][318]<=Wgt_2_318;WeightsStore[2][319]<=Wgt_2_319;WeightsStore[2][320]<=Wgt_2_320;WeightsStore[2][321]<=Wgt_2_321;WeightsStore[2][322]<=Wgt_2_322;WeightsStore[2][323]<=Wgt_2_323;WeightsStore[2][324]<=Wgt_2_324;WeightsStore[2][325]<=Wgt_2_325;WeightsStore[2][326]<=Wgt_2_326;WeightsStore[2][327]<=Wgt_2_327;WeightsStore[2][328]<=Wgt_2_328;WeightsStore[2][329]<=Wgt_2_329;WeightsStore[2][330]<=Wgt_2_330;WeightsStore[2][331]<=Wgt_2_331;WeightsStore[2][332]<=Wgt_2_332;WeightsStore[2][333]<=Wgt_2_333;WeightsStore[2][334]<=Wgt_2_334;WeightsStore[2][335]<=Wgt_2_335;WeightsStore[2][336]<=Wgt_2_336;WeightsStore[2][337]<=Wgt_2_337;WeightsStore[2][338]<=Wgt_2_338;WeightsStore[2][339]<=Wgt_2_339;WeightsStore[2][340]<=Wgt_2_340;WeightsStore[2][341]<=Wgt_2_341;WeightsStore[2][342]<=Wgt_2_342;WeightsStore[2][343]<=Wgt_2_343;WeightsStore[2][344]<=Wgt_2_344;WeightsStore[2][345]<=Wgt_2_345;WeightsStore[2][346]<=Wgt_2_346;WeightsStore[2][347]<=Wgt_2_347;WeightsStore[2][348]<=Wgt_2_348;WeightsStore[2][349]<=Wgt_2_349;WeightsStore[2][350]<=Wgt_2_350;WeightsStore[2][351]<=Wgt_2_351;WeightsStore[2][352]<=Wgt_2_352;WeightsStore[2][353]<=Wgt_2_353;WeightsStore[2][354]<=Wgt_2_354;WeightsStore[2][355]<=Wgt_2_355;WeightsStore[2][356]<=Wgt_2_356;WeightsStore[2][357]<=Wgt_2_357;WeightsStore[2][358]<=Wgt_2_358;WeightsStore[2][359]<=Wgt_2_359;WeightsStore[2][360]<=Wgt_2_360;WeightsStore[2][361]<=Wgt_2_361;WeightsStore[2][362]<=Wgt_2_362;WeightsStore[2][363]<=Wgt_2_363;WeightsStore[2][364]<=Wgt_2_364;WeightsStore[2][365]<=Wgt_2_365;WeightsStore[2][366]<=Wgt_2_366;WeightsStore[2][367]<=Wgt_2_367;WeightsStore[2][368]<=Wgt_2_368;WeightsStore[2][369]<=Wgt_2_369;WeightsStore[2][370]<=Wgt_2_370;WeightsStore[2][371]<=Wgt_2_371;WeightsStore[2][372]<=Wgt_2_372;WeightsStore[2][373]<=Wgt_2_373;WeightsStore[2][374]<=Wgt_2_374;WeightsStore[2][375]<=Wgt_2_375;WeightsStore[2][376]<=Wgt_2_376;WeightsStore[2][377]<=Wgt_2_377;WeightsStore[2][378]<=Wgt_2_378;WeightsStore[2][379]<=Wgt_2_379;WeightsStore[2][380]<=Wgt_2_380;WeightsStore[2][381]<=Wgt_2_381;WeightsStore[2][382]<=Wgt_2_382;WeightsStore[2][383]<=Wgt_2_383;WeightsStore[2][384]<=Wgt_2_384;WeightsStore[2][385]<=Wgt_2_385;WeightsStore[2][386]<=Wgt_2_386;WeightsStore[2][387]<=Wgt_2_387;WeightsStore[2][388]<=Wgt_2_388;WeightsStore[2][389]<=Wgt_2_389;WeightsStore[2][390]<=Wgt_2_390;WeightsStore[2][391]<=Wgt_2_391;WeightsStore[2][392]<=Wgt_2_392;WeightsStore[2][393]<=Wgt_2_393;WeightsStore[2][394]<=Wgt_2_394;WeightsStore[2][395]<=Wgt_2_395;WeightsStore[2][396]<=Wgt_2_396;WeightsStore[2][397]<=Wgt_2_397;WeightsStore[2][398]<=Wgt_2_398;WeightsStore[2][399]<=Wgt_2_399;WeightsStore[2][400]<=Wgt_2_400;WeightsStore[2][401]<=Wgt_2_401;WeightsStore[2][402]<=Wgt_2_402;WeightsStore[2][403]<=Wgt_2_403;WeightsStore[2][404]<=Wgt_2_404;WeightsStore[2][405]<=Wgt_2_405;WeightsStore[2][406]<=Wgt_2_406;WeightsStore[2][407]<=Wgt_2_407;WeightsStore[2][408]<=Wgt_2_408;WeightsStore[2][409]<=Wgt_2_409;WeightsStore[2][410]<=Wgt_2_410;WeightsStore[2][411]<=Wgt_2_411;WeightsStore[2][412]<=Wgt_2_412;WeightsStore[2][413]<=Wgt_2_413;WeightsStore[2][414]<=Wgt_2_414;WeightsStore[2][415]<=Wgt_2_415;WeightsStore[2][416]<=Wgt_2_416;WeightsStore[2][417]<=Wgt_2_417;WeightsStore[2][418]<=Wgt_2_418;WeightsStore[2][419]<=Wgt_2_419;WeightsStore[2][420]<=Wgt_2_420;WeightsStore[2][421]<=Wgt_2_421;WeightsStore[2][422]<=Wgt_2_422;WeightsStore[2][423]<=Wgt_2_423;WeightsStore[2][424]<=Wgt_2_424;WeightsStore[2][425]<=Wgt_2_425;WeightsStore[2][426]<=Wgt_2_426;WeightsStore[2][427]<=Wgt_2_427;WeightsStore[2][428]<=Wgt_2_428;WeightsStore[2][429]<=Wgt_2_429;WeightsStore[2][430]<=Wgt_2_430;WeightsStore[2][431]<=Wgt_2_431;WeightsStore[2][432]<=Wgt_2_432;WeightsStore[2][433]<=Wgt_2_433;WeightsStore[2][434]<=Wgt_2_434;WeightsStore[2][435]<=Wgt_2_435;WeightsStore[2][436]<=Wgt_2_436;WeightsStore[2][437]<=Wgt_2_437;WeightsStore[2][438]<=Wgt_2_438;WeightsStore[2][439]<=Wgt_2_439;WeightsStore[2][440]<=Wgt_2_440;WeightsStore[2][441]<=Wgt_2_441;WeightsStore[2][442]<=Wgt_2_442;WeightsStore[2][443]<=Wgt_2_443;WeightsStore[2][444]<=Wgt_2_444;WeightsStore[2][445]<=Wgt_2_445;WeightsStore[2][446]<=Wgt_2_446;WeightsStore[2][447]<=Wgt_2_447;WeightsStore[2][448]<=Wgt_2_448;WeightsStore[2][449]<=Wgt_2_449;WeightsStore[2][450]<=Wgt_2_450;WeightsStore[2][451]<=Wgt_2_451;WeightsStore[2][452]<=Wgt_2_452;WeightsStore[2][453]<=Wgt_2_453;WeightsStore[2][454]<=Wgt_2_454;WeightsStore[2][455]<=Wgt_2_455;WeightsStore[2][456]<=Wgt_2_456;WeightsStore[2][457]<=Wgt_2_457;WeightsStore[2][458]<=Wgt_2_458;WeightsStore[2][459]<=Wgt_2_459;WeightsStore[2][460]<=Wgt_2_460;WeightsStore[2][461]<=Wgt_2_461;WeightsStore[2][462]<=Wgt_2_462;WeightsStore[2][463]<=Wgt_2_463;WeightsStore[2][464]<=Wgt_2_464;WeightsStore[2][465]<=Wgt_2_465;WeightsStore[2][466]<=Wgt_2_466;WeightsStore[2][467]<=Wgt_2_467;WeightsStore[2][468]<=Wgt_2_468;WeightsStore[2][469]<=Wgt_2_469;WeightsStore[2][470]<=Wgt_2_470;WeightsStore[2][471]<=Wgt_2_471;WeightsStore[2][472]<=Wgt_2_472;WeightsStore[2][473]<=Wgt_2_473;WeightsStore[2][474]<=Wgt_2_474;WeightsStore[2][475]<=Wgt_2_475;WeightsStore[2][476]<=Wgt_2_476;WeightsStore[2][477]<=Wgt_2_477;WeightsStore[2][478]<=Wgt_2_478;WeightsStore[2][479]<=Wgt_2_479;WeightsStore[2][480]<=Wgt_2_480;WeightsStore[2][481]<=Wgt_2_481;WeightsStore[2][482]<=Wgt_2_482;WeightsStore[2][483]<=Wgt_2_483;WeightsStore[2][484]<=Wgt_2_484;WeightsStore[2][485]<=Wgt_2_485;WeightsStore[2][486]<=Wgt_2_486;WeightsStore[2][487]<=Wgt_2_487;WeightsStore[2][488]<=Wgt_2_488;WeightsStore[2][489]<=Wgt_2_489;WeightsStore[2][490]<=Wgt_2_490;WeightsStore[2][491]<=Wgt_2_491;WeightsStore[2][492]<=Wgt_2_492;WeightsStore[2][493]<=Wgt_2_493;WeightsStore[2][494]<=Wgt_2_494;WeightsStore[2][495]<=Wgt_2_495;WeightsStore[2][496]<=Wgt_2_496;WeightsStore[2][497]<=Wgt_2_497;WeightsStore[2][498]<=Wgt_2_498;WeightsStore[2][499]<=Wgt_2_499;WeightsStore[2][500]<=Wgt_2_500;WeightsStore[2][501]<=Wgt_2_501;WeightsStore[2][502]<=Wgt_2_502;WeightsStore[2][503]<=Wgt_2_503;WeightsStore[2][504]<=Wgt_2_504;WeightsStore[2][505]<=Wgt_2_505;WeightsStore[2][506]<=Wgt_2_506;WeightsStore[2][507]<=Wgt_2_507;WeightsStore[2][508]<=Wgt_2_508;WeightsStore[2][509]<=Wgt_2_509;WeightsStore[2][510]<=Wgt_2_510;WeightsStore[2][511]<=Wgt_2_511;WeightsStore[2][512]<=Wgt_2_512;WeightsStore[2][513]<=Wgt_2_513;WeightsStore[2][514]<=Wgt_2_514;WeightsStore[2][515]<=Wgt_2_515;WeightsStore[2][516]<=Wgt_2_516;WeightsStore[2][517]<=Wgt_2_517;WeightsStore[2][518]<=Wgt_2_518;WeightsStore[2][519]<=Wgt_2_519;WeightsStore[2][520]<=Wgt_2_520;WeightsStore[2][521]<=Wgt_2_521;WeightsStore[2][522]<=Wgt_2_522;WeightsStore[2][523]<=Wgt_2_523;WeightsStore[2][524]<=Wgt_2_524;WeightsStore[2][525]<=Wgt_2_525;WeightsStore[2][526]<=Wgt_2_526;WeightsStore[2][527]<=Wgt_2_527;WeightsStore[2][528]<=Wgt_2_528;WeightsStore[2][529]<=Wgt_2_529;WeightsStore[2][530]<=Wgt_2_530;WeightsStore[2][531]<=Wgt_2_531;WeightsStore[2][532]<=Wgt_2_532;WeightsStore[2][533]<=Wgt_2_533;WeightsStore[2][534]<=Wgt_2_534;WeightsStore[2][535]<=Wgt_2_535;WeightsStore[2][536]<=Wgt_2_536;WeightsStore[2][537]<=Wgt_2_537;WeightsStore[2][538]<=Wgt_2_538;WeightsStore[2][539]<=Wgt_2_539;WeightsStore[2][540]<=Wgt_2_540;WeightsStore[2][541]<=Wgt_2_541;WeightsStore[2][542]<=Wgt_2_542;WeightsStore[2][543]<=Wgt_2_543;WeightsStore[2][544]<=Wgt_2_544;WeightsStore[2][545]<=Wgt_2_545;WeightsStore[2][546]<=Wgt_2_546;WeightsStore[2][547]<=Wgt_2_547;WeightsStore[2][548]<=Wgt_2_548;WeightsStore[2][549]<=Wgt_2_549;WeightsStore[2][550]<=Wgt_2_550;WeightsStore[2][551]<=Wgt_2_551;WeightsStore[2][552]<=Wgt_2_552;WeightsStore[2][553]<=Wgt_2_553;WeightsStore[2][554]<=Wgt_2_554;WeightsStore[2][555]<=Wgt_2_555;WeightsStore[2][556]<=Wgt_2_556;WeightsStore[2][557]<=Wgt_2_557;WeightsStore[2][558]<=Wgt_2_558;WeightsStore[2][559]<=Wgt_2_559;WeightsStore[2][560]<=Wgt_2_560;WeightsStore[2][561]<=Wgt_2_561;WeightsStore[2][562]<=Wgt_2_562;WeightsStore[2][563]<=Wgt_2_563;WeightsStore[2][564]<=Wgt_2_564;WeightsStore[2][565]<=Wgt_2_565;WeightsStore[2][566]<=Wgt_2_566;WeightsStore[2][567]<=Wgt_2_567;WeightsStore[2][568]<=Wgt_2_568;WeightsStore[2][569]<=Wgt_2_569;WeightsStore[2][570]<=Wgt_2_570;WeightsStore[2][571]<=Wgt_2_571;WeightsStore[2][572]<=Wgt_2_572;WeightsStore[2][573]<=Wgt_2_573;WeightsStore[2][574]<=Wgt_2_574;WeightsStore[2][575]<=Wgt_2_575;WeightsStore[2][576]<=Wgt_2_576;WeightsStore[2][577]<=Wgt_2_577;WeightsStore[2][578]<=Wgt_2_578;WeightsStore[2][579]<=Wgt_2_579;WeightsStore[2][580]<=Wgt_2_580;WeightsStore[2][581]<=Wgt_2_581;WeightsStore[2][582]<=Wgt_2_582;WeightsStore[2][583]<=Wgt_2_583;WeightsStore[2][584]<=Wgt_2_584;WeightsStore[2][585]<=Wgt_2_585;WeightsStore[2][586]<=Wgt_2_586;WeightsStore[2][587]<=Wgt_2_587;WeightsStore[2][588]<=Wgt_2_588;WeightsStore[2][589]<=Wgt_2_589;WeightsStore[2][590]<=Wgt_2_590;WeightsStore[2][591]<=Wgt_2_591;WeightsStore[2][592]<=Wgt_2_592;WeightsStore[2][593]<=Wgt_2_593;WeightsStore[2][594]<=Wgt_2_594;WeightsStore[2][595]<=Wgt_2_595;WeightsStore[2][596]<=Wgt_2_596;WeightsStore[2][597]<=Wgt_2_597;WeightsStore[2][598]<=Wgt_2_598;WeightsStore[2][599]<=Wgt_2_599;WeightsStore[2][600]<=Wgt_2_600;WeightsStore[2][601]<=Wgt_2_601;WeightsStore[2][602]<=Wgt_2_602;WeightsStore[2][603]<=Wgt_2_603;WeightsStore[2][604]<=Wgt_2_604;WeightsStore[2][605]<=Wgt_2_605;WeightsStore[2][606]<=Wgt_2_606;WeightsStore[2][607]<=Wgt_2_607;WeightsStore[2][608]<=Wgt_2_608;WeightsStore[2][609]<=Wgt_2_609;WeightsStore[2][610]<=Wgt_2_610;WeightsStore[2][611]<=Wgt_2_611;WeightsStore[2][612]<=Wgt_2_612;WeightsStore[2][613]<=Wgt_2_613;WeightsStore[2][614]<=Wgt_2_614;WeightsStore[2][615]<=Wgt_2_615;WeightsStore[2][616]<=Wgt_2_616;WeightsStore[2][617]<=Wgt_2_617;WeightsStore[2][618]<=Wgt_2_618;WeightsStore[2][619]<=Wgt_2_619;WeightsStore[2][620]<=Wgt_2_620;WeightsStore[2][621]<=Wgt_2_621;WeightsStore[2][622]<=Wgt_2_622;WeightsStore[2][623]<=Wgt_2_623;WeightsStore[2][624]<=Wgt_2_624;WeightsStore[2][625]<=Wgt_2_625;WeightsStore[2][626]<=Wgt_2_626;WeightsStore[2][627]<=Wgt_2_627;WeightsStore[2][628]<=Wgt_2_628;WeightsStore[2][629]<=Wgt_2_629;WeightsStore[2][630]<=Wgt_2_630;WeightsStore[2][631]<=Wgt_2_631;WeightsStore[2][632]<=Wgt_2_632;WeightsStore[2][633]<=Wgt_2_633;WeightsStore[2][634]<=Wgt_2_634;WeightsStore[2][635]<=Wgt_2_635;WeightsStore[2][636]<=Wgt_2_636;WeightsStore[2][637]<=Wgt_2_637;WeightsStore[2][638]<=Wgt_2_638;WeightsStore[2][639]<=Wgt_2_639;WeightsStore[2][640]<=Wgt_2_640;WeightsStore[2][641]<=Wgt_2_641;WeightsStore[2][642]<=Wgt_2_642;WeightsStore[2][643]<=Wgt_2_643;WeightsStore[2][644]<=Wgt_2_644;WeightsStore[2][645]<=Wgt_2_645;WeightsStore[2][646]<=Wgt_2_646;WeightsStore[2][647]<=Wgt_2_647;WeightsStore[2][648]<=Wgt_2_648;WeightsStore[2][649]<=Wgt_2_649;WeightsStore[2][650]<=Wgt_2_650;WeightsStore[2][651]<=Wgt_2_651;WeightsStore[2][652]<=Wgt_2_652;WeightsStore[2][653]<=Wgt_2_653;WeightsStore[2][654]<=Wgt_2_654;WeightsStore[2][655]<=Wgt_2_655;WeightsStore[2][656]<=Wgt_2_656;WeightsStore[2][657]<=Wgt_2_657;WeightsStore[2][658]<=Wgt_2_658;WeightsStore[2][659]<=Wgt_2_659;WeightsStore[2][660]<=Wgt_2_660;WeightsStore[2][661]<=Wgt_2_661;WeightsStore[2][662]<=Wgt_2_662;WeightsStore[2][663]<=Wgt_2_663;WeightsStore[2][664]<=Wgt_2_664;WeightsStore[2][665]<=Wgt_2_665;WeightsStore[2][666]<=Wgt_2_666;WeightsStore[2][667]<=Wgt_2_667;WeightsStore[2][668]<=Wgt_2_668;WeightsStore[2][669]<=Wgt_2_669;WeightsStore[2][670]<=Wgt_2_670;WeightsStore[2][671]<=Wgt_2_671;WeightsStore[2][672]<=Wgt_2_672;WeightsStore[2][673]<=Wgt_2_673;WeightsStore[2][674]<=Wgt_2_674;WeightsStore[2][675]<=Wgt_2_675;WeightsStore[2][676]<=Wgt_2_676;WeightsStore[2][677]<=Wgt_2_677;WeightsStore[2][678]<=Wgt_2_678;WeightsStore[2][679]<=Wgt_2_679;WeightsStore[2][680]<=Wgt_2_680;WeightsStore[2][681]<=Wgt_2_681;WeightsStore[2][682]<=Wgt_2_682;WeightsStore[2][683]<=Wgt_2_683;WeightsStore[2][684]<=Wgt_2_684;WeightsStore[2][685]<=Wgt_2_685;WeightsStore[2][686]<=Wgt_2_686;WeightsStore[2][687]<=Wgt_2_687;WeightsStore[2][688]<=Wgt_2_688;WeightsStore[2][689]<=Wgt_2_689;WeightsStore[2][690]<=Wgt_2_690;WeightsStore[2][691]<=Wgt_2_691;WeightsStore[2][692]<=Wgt_2_692;WeightsStore[2][693]<=Wgt_2_693;WeightsStore[2][694]<=Wgt_2_694;WeightsStore[2][695]<=Wgt_2_695;WeightsStore[2][696]<=Wgt_2_696;WeightsStore[2][697]<=Wgt_2_697;WeightsStore[2][698]<=Wgt_2_698;WeightsStore[2][699]<=Wgt_2_699;WeightsStore[2][700]<=Wgt_2_700;WeightsStore[2][701]<=Wgt_2_701;WeightsStore[2][702]<=Wgt_2_702;WeightsStore[2][703]<=Wgt_2_703;WeightsStore[2][704]<=Wgt_2_704;WeightsStore[2][705]<=Wgt_2_705;WeightsStore[2][706]<=Wgt_2_706;WeightsStore[2][707]<=Wgt_2_707;WeightsStore[2][708]<=Wgt_2_708;WeightsStore[2][709]<=Wgt_2_709;WeightsStore[2][710]<=Wgt_2_710;WeightsStore[2][711]<=Wgt_2_711;WeightsStore[2][712]<=Wgt_2_712;WeightsStore[2][713]<=Wgt_2_713;WeightsStore[2][714]<=Wgt_2_714;WeightsStore[2][715]<=Wgt_2_715;WeightsStore[2][716]<=Wgt_2_716;WeightsStore[2][717]<=Wgt_2_717;WeightsStore[2][718]<=Wgt_2_718;WeightsStore[2][719]<=Wgt_2_719;WeightsStore[2][720]<=Wgt_2_720;WeightsStore[2][721]<=Wgt_2_721;WeightsStore[2][722]<=Wgt_2_722;WeightsStore[2][723]<=Wgt_2_723;WeightsStore[2][724]<=Wgt_2_724;WeightsStore[2][725]<=Wgt_2_725;WeightsStore[2][726]<=Wgt_2_726;WeightsStore[2][727]<=Wgt_2_727;WeightsStore[2][728]<=Wgt_2_728;WeightsStore[2][729]<=Wgt_2_729;WeightsStore[2][730]<=Wgt_2_730;WeightsStore[2][731]<=Wgt_2_731;WeightsStore[2][732]<=Wgt_2_732;WeightsStore[2][733]<=Wgt_2_733;WeightsStore[2][734]<=Wgt_2_734;WeightsStore[2][735]<=Wgt_2_735;WeightsStore[2][736]<=Wgt_2_736;WeightsStore[2][737]<=Wgt_2_737;WeightsStore[2][738]<=Wgt_2_738;WeightsStore[2][739]<=Wgt_2_739;WeightsStore[2][740]<=Wgt_2_740;WeightsStore[2][741]<=Wgt_2_741;WeightsStore[2][742]<=Wgt_2_742;WeightsStore[2][743]<=Wgt_2_743;WeightsStore[2][744]<=Wgt_2_744;WeightsStore[2][745]<=Wgt_2_745;WeightsStore[2][746]<=Wgt_2_746;WeightsStore[2][747]<=Wgt_2_747;WeightsStore[2][748]<=Wgt_2_748;WeightsStore[2][749]<=Wgt_2_749;WeightsStore[2][750]<=Wgt_2_750;WeightsStore[2][751]<=Wgt_2_751;WeightsStore[2][752]<=Wgt_2_752;WeightsStore[2][753]<=Wgt_2_753;WeightsStore[2][754]<=Wgt_2_754;WeightsStore[2][755]<=Wgt_2_755;WeightsStore[2][756]<=Wgt_2_756;WeightsStore[2][757]<=Wgt_2_757;WeightsStore[2][758]<=Wgt_2_758;WeightsStore[2][759]<=Wgt_2_759;WeightsStore[2][760]<=Wgt_2_760;WeightsStore[2][761]<=Wgt_2_761;WeightsStore[2][762]<=Wgt_2_762;WeightsStore[2][763]<=Wgt_2_763;WeightsStore[2][764]<=Wgt_2_764;WeightsStore[2][765]<=Wgt_2_765;WeightsStore[2][766]<=Wgt_2_766;WeightsStore[2][767]<=Wgt_2_767;WeightsStore[2][768]<=Wgt_2_768;WeightsStore[2][769]<=Wgt_2_769;WeightsStore[2][770]<=Wgt_2_770;WeightsStore[2][771]<=Wgt_2_771;WeightsStore[2][772]<=Wgt_2_772;WeightsStore[2][773]<=Wgt_2_773;WeightsStore[2][774]<=Wgt_2_774;WeightsStore[2][775]<=Wgt_2_775;WeightsStore[2][776]<=Wgt_2_776;WeightsStore[2][777]<=Wgt_2_777;WeightsStore[2][778]<=Wgt_2_778;WeightsStore[2][779]<=Wgt_2_779;WeightsStore[2][780]<=Wgt_2_780;WeightsStore[2][781]<=Wgt_2_781;WeightsStore[2][782]<=Wgt_2_782;WeightsStore[2][783]<=Wgt_2_783;WeightsStore[2][784]<=Wgt_2_784;WeightsStore[3][0]<=Wgt_3_0;WeightsStore[3][1]<=Wgt_3_1;WeightsStore[3][2]<=Wgt_3_2;WeightsStore[3][3]<=Wgt_3_3;WeightsStore[3][4]<=Wgt_3_4;WeightsStore[3][5]<=Wgt_3_5;WeightsStore[3][6]<=Wgt_3_6;WeightsStore[3][7]<=Wgt_3_7;WeightsStore[3][8]<=Wgt_3_8;WeightsStore[3][9]<=Wgt_3_9;WeightsStore[3][10]<=Wgt_3_10;WeightsStore[3][11]<=Wgt_3_11;WeightsStore[3][12]<=Wgt_3_12;WeightsStore[3][13]<=Wgt_3_13;WeightsStore[3][14]<=Wgt_3_14;WeightsStore[3][15]<=Wgt_3_15;WeightsStore[3][16]<=Wgt_3_16;WeightsStore[3][17]<=Wgt_3_17;WeightsStore[3][18]<=Wgt_3_18;WeightsStore[3][19]<=Wgt_3_19;WeightsStore[3][20]<=Wgt_3_20;WeightsStore[3][21]<=Wgt_3_21;WeightsStore[3][22]<=Wgt_3_22;WeightsStore[3][23]<=Wgt_3_23;WeightsStore[3][24]<=Wgt_3_24;WeightsStore[3][25]<=Wgt_3_25;WeightsStore[3][26]<=Wgt_3_26;WeightsStore[3][27]<=Wgt_3_27;WeightsStore[3][28]<=Wgt_3_28;WeightsStore[3][29]<=Wgt_3_29;WeightsStore[3][30]<=Wgt_3_30;WeightsStore[3][31]<=Wgt_3_31;WeightsStore[3][32]<=Wgt_3_32;WeightsStore[3][33]<=Wgt_3_33;WeightsStore[3][34]<=Wgt_3_34;WeightsStore[3][35]<=Wgt_3_35;WeightsStore[3][36]<=Wgt_3_36;WeightsStore[3][37]<=Wgt_3_37;WeightsStore[3][38]<=Wgt_3_38;WeightsStore[3][39]<=Wgt_3_39;WeightsStore[3][40]<=Wgt_3_40;WeightsStore[3][41]<=Wgt_3_41;WeightsStore[3][42]<=Wgt_3_42;WeightsStore[3][43]<=Wgt_3_43;WeightsStore[3][44]<=Wgt_3_44;WeightsStore[3][45]<=Wgt_3_45;WeightsStore[3][46]<=Wgt_3_46;WeightsStore[3][47]<=Wgt_3_47;WeightsStore[3][48]<=Wgt_3_48;WeightsStore[3][49]<=Wgt_3_49;WeightsStore[3][50]<=Wgt_3_50;WeightsStore[3][51]<=Wgt_3_51;WeightsStore[3][52]<=Wgt_3_52;WeightsStore[3][53]<=Wgt_3_53;WeightsStore[3][54]<=Wgt_3_54;WeightsStore[3][55]<=Wgt_3_55;WeightsStore[3][56]<=Wgt_3_56;WeightsStore[3][57]<=Wgt_3_57;WeightsStore[3][58]<=Wgt_3_58;WeightsStore[3][59]<=Wgt_3_59;WeightsStore[3][60]<=Wgt_3_60;WeightsStore[3][61]<=Wgt_3_61;WeightsStore[3][62]<=Wgt_3_62;WeightsStore[3][63]<=Wgt_3_63;WeightsStore[3][64]<=Wgt_3_64;WeightsStore[3][65]<=Wgt_3_65;WeightsStore[3][66]<=Wgt_3_66;WeightsStore[3][67]<=Wgt_3_67;WeightsStore[3][68]<=Wgt_3_68;WeightsStore[3][69]<=Wgt_3_69;WeightsStore[3][70]<=Wgt_3_70;WeightsStore[3][71]<=Wgt_3_71;WeightsStore[3][72]<=Wgt_3_72;WeightsStore[3][73]<=Wgt_3_73;WeightsStore[3][74]<=Wgt_3_74;WeightsStore[3][75]<=Wgt_3_75;WeightsStore[3][76]<=Wgt_3_76;WeightsStore[3][77]<=Wgt_3_77;WeightsStore[3][78]<=Wgt_3_78;WeightsStore[3][79]<=Wgt_3_79;WeightsStore[3][80]<=Wgt_3_80;WeightsStore[3][81]<=Wgt_3_81;WeightsStore[3][82]<=Wgt_3_82;WeightsStore[3][83]<=Wgt_3_83;WeightsStore[3][84]<=Wgt_3_84;WeightsStore[3][85]<=Wgt_3_85;WeightsStore[3][86]<=Wgt_3_86;WeightsStore[3][87]<=Wgt_3_87;WeightsStore[3][88]<=Wgt_3_88;WeightsStore[3][89]<=Wgt_3_89;WeightsStore[3][90]<=Wgt_3_90;WeightsStore[3][91]<=Wgt_3_91;WeightsStore[3][92]<=Wgt_3_92;WeightsStore[3][93]<=Wgt_3_93;WeightsStore[3][94]<=Wgt_3_94;WeightsStore[3][95]<=Wgt_3_95;WeightsStore[3][96]<=Wgt_3_96;WeightsStore[3][97]<=Wgt_3_97;WeightsStore[3][98]<=Wgt_3_98;WeightsStore[3][99]<=Wgt_3_99;WeightsStore[3][100]<=Wgt_3_100;WeightsStore[3][101]<=Wgt_3_101;WeightsStore[3][102]<=Wgt_3_102;WeightsStore[3][103]<=Wgt_3_103;WeightsStore[3][104]<=Wgt_3_104;WeightsStore[3][105]<=Wgt_3_105;WeightsStore[3][106]<=Wgt_3_106;WeightsStore[3][107]<=Wgt_3_107;WeightsStore[3][108]<=Wgt_3_108;WeightsStore[3][109]<=Wgt_3_109;WeightsStore[3][110]<=Wgt_3_110;WeightsStore[3][111]<=Wgt_3_111;WeightsStore[3][112]<=Wgt_3_112;WeightsStore[3][113]<=Wgt_3_113;WeightsStore[3][114]<=Wgt_3_114;WeightsStore[3][115]<=Wgt_3_115;WeightsStore[3][116]<=Wgt_3_116;WeightsStore[3][117]<=Wgt_3_117;WeightsStore[3][118]<=Wgt_3_118;WeightsStore[3][119]<=Wgt_3_119;WeightsStore[3][120]<=Wgt_3_120;WeightsStore[3][121]<=Wgt_3_121;WeightsStore[3][122]<=Wgt_3_122;WeightsStore[3][123]<=Wgt_3_123;WeightsStore[3][124]<=Wgt_3_124;WeightsStore[3][125]<=Wgt_3_125;WeightsStore[3][126]<=Wgt_3_126;WeightsStore[3][127]<=Wgt_3_127;WeightsStore[3][128]<=Wgt_3_128;WeightsStore[3][129]<=Wgt_3_129;WeightsStore[3][130]<=Wgt_3_130;WeightsStore[3][131]<=Wgt_3_131;WeightsStore[3][132]<=Wgt_3_132;WeightsStore[3][133]<=Wgt_3_133;WeightsStore[3][134]<=Wgt_3_134;WeightsStore[3][135]<=Wgt_3_135;WeightsStore[3][136]<=Wgt_3_136;WeightsStore[3][137]<=Wgt_3_137;WeightsStore[3][138]<=Wgt_3_138;WeightsStore[3][139]<=Wgt_3_139;WeightsStore[3][140]<=Wgt_3_140;WeightsStore[3][141]<=Wgt_3_141;WeightsStore[3][142]<=Wgt_3_142;WeightsStore[3][143]<=Wgt_3_143;WeightsStore[3][144]<=Wgt_3_144;WeightsStore[3][145]<=Wgt_3_145;WeightsStore[3][146]<=Wgt_3_146;WeightsStore[3][147]<=Wgt_3_147;WeightsStore[3][148]<=Wgt_3_148;WeightsStore[3][149]<=Wgt_3_149;WeightsStore[3][150]<=Wgt_3_150;WeightsStore[3][151]<=Wgt_3_151;WeightsStore[3][152]<=Wgt_3_152;WeightsStore[3][153]<=Wgt_3_153;WeightsStore[3][154]<=Wgt_3_154;WeightsStore[3][155]<=Wgt_3_155;WeightsStore[3][156]<=Wgt_3_156;WeightsStore[3][157]<=Wgt_3_157;WeightsStore[3][158]<=Wgt_3_158;WeightsStore[3][159]<=Wgt_3_159;WeightsStore[3][160]<=Wgt_3_160;WeightsStore[3][161]<=Wgt_3_161;WeightsStore[3][162]<=Wgt_3_162;WeightsStore[3][163]<=Wgt_3_163;WeightsStore[3][164]<=Wgt_3_164;WeightsStore[3][165]<=Wgt_3_165;WeightsStore[3][166]<=Wgt_3_166;WeightsStore[3][167]<=Wgt_3_167;WeightsStore[3][168]<=Wgt_3_168;WeightsStore[3][169]<=Wgt_3_169;WeightsStore[3][170]<=Wgt_3_170;WeightsStore[3][171]<=Wgt_3_171;WeightsStore[3][172]<=Wgt_3_172;WeightsStore[3][173]<=Wgt_3_173;WeightsStore[3][174]<=Wgt_3_174;WeightsStore[3][175]<=Wgt_3_175;WeightsStore[3][176]<=Wgt_3_176;WeightsStore[3][177]<=Wgt_3_177;WeightsStore[3][178]<=Wgt_3_178;WeightsStore[3][179]<=Wgt_3_179;WeightsStore[3][180]<=Wgt_3_180;WeightsStore[3][181]<=Wgt_3_181;WeightsStore[3][182]<=Wgt_3_182;WeightsStore[3][183]<=Wgt_3_183;WeightsStore[3][184]<=Wgt_3_184;WeightsStore[3][185]<=Wgt_3_185;WeightsStore[3][186]<=Wgt_3_186;WeightsStore[3][187]<=Wgt_3_187;WeightsStore[3][188]<=Wgt_3_188;WeightsStore[3][189]<=Wgt_3_189;WeightsStore[3][190]<=Wgt_3_190;WeightsStore[3][191]<=Wgt_3_191;WeightsStore[3][192]<=Wgt_3_192;WeightsStore[3][193]<=Wgt_3_193;WeightsStore[3][194]<=Wgt_3_194;WeightsStore[3][195]<=Wgt_3_195;WeightsStore[3][196]<=Wgt_3_196;WeightsStore[3][197]<=Wgt_3_197;WeightsStore[3][198]<=Wgt_3_198;WeightsStore[3][199]<=Wgt_3_199;WeightsStore[3][200]<=Wgt_3_200;WeightsStore[3][201]<=Wgt_3_201;WeightsStore[3][202]<=Wgt_3_202;WeightsStore[3][203]<=Wgt_3_203;WeightsStore[3][204]<=Wgt_3_204;WeightsStore[3][205]<=Wgt_3_205;WeightsStore[3][206]<=Wgt_3_206;WeightsStore[3][207]<=Wgt_3_207;WeightsStore[3][208]<=Wgt_3_208;WeightsStore[3][209]<=Wgt_3_209;WeightsStore[3][210]<=Wgt_3_210;WeightsStore[3][211]<=Wgt_3_211;WeightsStore[3][212]<=Wgt_3_212;WeightsStore[3][213]<=Wgt_3_213;WeightsStore[3][214]<=Wgt_3_214;WeightsStore[3][215]<=Wgt_3_215;WeightsStore[3][216]<=Wgt_3_216;WeightsStore[3][217]<=Wgt_3_217;WeightsStore[3][218]<=Wgt_3_218;WeightsStore[3][219]<=Wgt_3_219;WeightsStore[3][220]<=Wgt_3_220;WeightsStore[3][221]<=Wgt_3_221;WeightsStore[3][222]<=Wgt_3_222;WeightsStore[3][223]<=Wgt_3_223;WeightsStore[3][224]<=Wgt_3_224;WeightsStore[3][225]<=Wgt_3_225;WeightsStore[3][226]<=Wgt_3_226;WeightsStore[3][227]<=Wgt_3_227;WeightsStore[3][228]<=Wgt_3_228;WeightsStore[3][229]<=Wgt_3_229;WeightsStore[3][230]<=Wgt_3_230;WeightsStore[3][231]<=Wgt_3_231;WeightsStore[3][232]<=Wgt_3_232;WeightsStore[3][233]<=Wgt_3_233;WeightsStore[3][234]<=Wgt_3_234;WeightsStore[3][235]<=Wgt_3_235;WeightsStore[3][236]<=Wgt_3_236;WeightsStore[3][237]<=Wgt_3_237;WeightsStore[3][238]<=Wgt_3_238;WeightsStore[3][239]<=Wgt_3_239;WeightsStore[3][240]<=Wgt_3_240;WeightsStore[3][241]<=Wgt_3_241;WeightsStore[3][242]<=Wgt_3_242;WeightsStore[3][243]<=Wgt_3_243;WeightsStore[3][244]<=Wgt_3_244;WeightsStore[3][245]<=Wgt_3_245;WeightsStore[3][246]<=Wgt_3_246;WeightsStore[3][247]<=Wgt_3_247;WeightsStore[3][248]<=Wgt_3_248;WeightsStore[3][249]<=Wgt_3_249;WeightsStore[3][250]<=Wgt_3_250;WeightsStore[3][251]<=Wgt_3_251;WeightsStore[3][252]<=Wgt_3_252;WeightsStore[3][253]<=Wgt_3_253;WeightsStore[3][254]<=Wgt_3_254;WeightsStore[3][255]<=Wgt_3_255;WeightsStore[3][256]<=Wgt_3_256;WeightsStore[3][257]<=Wgt_3_257;WeightsStore[3][258]<=Wgt_3_258;WeightsStore[3][259]<=Wgt_3_259;WeightsStore[3][260]<=Wgt_3_260;WeightsStore[3][261]<=Wgt_3_261;WeightsStore[3][262]<=Wgt_3_262;WeightsStore[3][263]<=Wgt_3_263;WeightsStore[3][264]<=Wgt_3_264;WeightsStore[3][265]<=Wgt_3_265;WeightsStore[3][266]<=Wgt_3_266;WeightsStore[3][267]<=Wgt_3_267;WeightsStore[3][268]<=Wgt_3_268;WeightsStore[3][269]<=Wgt_3_269;WeightsStore[3][270]<=Wgt_3_270;WeightsStore[3][271]<=Wgt_3_271;WeightsStore[3][272]<=Wgt_3_272;WeightsStore[3][273]<=Wgt_3_273;WeightsStore[3][274]<=Wgt_3_274;WeightsStore[3][275]<=Wgt_3_275;WeightsStore[3][276]<=Wgt_3_276;WeightsStore[3][277]<=Wgt_3_277;WeightsStore[3][278]<=Wgt_3_278;WeightsStore[3][279]<=Wgt_3_279;WeightsStore[3][280]<=Wgt_3_280;WeightsStore[3][281]<=Wgt_3_281;WeightsStore[3][282]<=Wgt_3_282;WeightsStore[3][283]<=Wgt_3_283;WeightsStore[3][284]<=Wgt_3_284;WeightsStore[3][285]<=Wgt_3_285;WeightsStore[3][286]<=Wgt_3_286;WeightsStore[3][287]<=Wgt_3_287;WeightsStore[3][288]<=Wgt_3_288;WeightsStore[3][289]<=Wgt_3_289;WeightsStore[3][290]<=Wgt_3_290;WeightsStore[3][291]<=Wgt_3_291;WeightsStore[3][292]<=Wgt_3_292;WeightsStore[3][293]<=Wgt_3_293;WeightsStore[3][294]<=Wgt_3_294;WeightsStore[3][295]<=Wgt_3_295;WeightsStore[3][296]<=Wgt_3_296;WeightsStore[3][297]<=Wgt_3_297;WeightsStore[3][298]<=Wgt_3_298;WeightsStore[3][299]<=Wgt_3_299;WeightsStore[3][300]<=Wgt_3_300;WeightsStore[3][301]<=Wgt_3_301;WeightsStore[3][302]<=Wgt_3_302;WeightsStore[3][303]<=Wgt_3_303;WeightsStore[3][304]<=Wgt_3_304;WeightsStore[3][305]<=Wgt_3_305;WeightsStore[3][306]<=Wgt_3_306;WeightsStore[3][307]<=Wgt_3_307;WeightsStore[3][308]<=Wgt_3_308;WeightsStore[3][309]<=Wgt_3_309;WeightsStore[3][310]<=Wgt_3_310;WeightsStore[3][311]<=Wgt_3_311;WeightsStore[3][312]<=Wgt_3_312;WeightsStore[3][313]<=Wgt_3_313;WeightsStore[3][314]<=Wgt_3_314;WeightsStore[3][315]<=Wgt_3_315;WeightsStore[3][316]<=Wgt_3_316;WeightsStore[3][317]<=Wgt_3_317;WeightsStore[3][318]<=Wgt_3_318;WeightsStore[3][319]<=Wgt_3_319;WeightsStore[3][320]<=Wgt_3_320;WeightsStore[3][321]<=Wgt_3_321;WeightsStore[3][322]<=Wgt_3_322;WeightsStore[3][323]<=Wgt_3_323;WeightsStore[3][324]<=Wgt_3_324;WeightsStore[3][325]<=Wgt_3_325;WeightsStore[3][326]<=Wgt_3_326;WeightsStore[3][327]<=Wgt_3_327;WeightsStore[3][328]<=Wgt_3_328;WeightsStore[3][329]<=Wgt_3_329;WeightsStore[3][330]<=Wgt_3_330;WeightsStore[3][331]<=Wgt_3_331;WeightsStore[3][332]<=Wgt_3_332;WeightsStore[3][333]<=Wgt_3_333;WeightsStore[3][334]<=Wgt_3_334;WeightsStore[3][335]<=Wgt_3_335;WeightsStore[3][336]<=Wgt_3_336;WeightsStore[3][337]<=Wgt_3_337;WeightsStore[3][338]<=Wgt_3_338;WeightsStore[3][339]<=Wgt_3_339;WeightsStore[3][340]<=Wgt_3_340;WeightsStore[3][341]<=Wgt_3_341;WeightsStore[3][342]<=Wgt_3_342;WeightsStore[3][343]<=Wgt_3_343;WeightsStore[3][344]<=Wgt_3_344;WeightsStore[3][345]<=Wgt_3_345;WeightsStore[3][346]<=Wgt_3_346;WeightsStore[3][347]<=Wgt_3_347;WeightsStore[3][348]<=Wgt_3_348;WeightsStore[3][349]<=Wgt_3_349;WeightsStore[3][350]<=Wgt_3_350;WeightsStore[3][351]<=Wgt_3_351;WeightsStore[3][352]<=Wgt_3_352;WeightsStore[3][353]<=Wgt_3_353;WeightsStore[3][354]<=Wgt_3_354;WeightsStore[3][355]<=Wgt_3_355;WeightsStore[3][356]<=Wgt_3_356;WeightsStore[3][357]<=Wgt_3_357;WeightsStore[3][358]<=Wgt_3_358;WeightsStore[3][359]<=Wgt_3_359;WeightsStore[3][360]<=Wgt_3_360;WeightsStore[3][361]<=Wgt_3_361;WeightsStore[3][362]<=Wgt_3_362;WeightsStore[3][363]<=Wgt_3_363;WeightsStore[3][364]<=Wgt_3_364;WeightsStore[3][365]<=Wgt_3_365;WeightsStore[3][366]<=Wgt_3_366;WeightsStore[3][367]<=Wgt_3_367;WeightsStore[3][368]<=Wgt_3_368;WeightsStore[3][369]<=Wgt_3_369;WeightsStore[3][370]<=Wgt_3_370;WeightsStore[3][371]<=Wgt_3_371;WeightsStore[3][372]<=Wgt_3_372;WeightsStore[3][373]<=Wgt_3_373;WeightsStore[3][374]<=Wgt_3_374;WeightsStore[3][375]<=Wgt_3_375;WeightsStore[3][376]<=Wgt_3_376;WeightsStore[3][377]<=Wgt_3_377;WeightsStore[3][378]<=Wgt_3_378;WeightsStore[3][379]<=Wgt_3_379;WeightsStore[3][380]<=Wgt_3_380;WeightsStore[3][381]<=Wgt_3_381;WeightsStore[3][382]<=Wgt_3_382;WeightsStore[3][383]<=Wgt_3_383;WeightsStore[3][384]<=Wgt_3_384;WeightsStore[3][385]<=Wgt_3_385;WeightsStore[3][386]<=Wgt_3_386;WeightsStore[3][387]<=Wgt_3_387;WeightsStore[3][388]<=Wgt_3_388;WeightsStore[3][389]<=Wgt_3_389;WeightsStore[3][390]<=Wgt_3_390;WeightsStore[3][391]<=Wgt_3_391;WeightsStore[3][392]<=Wgt_3_392;WeightsStore[3][393]<=Wgt_3_393;WeightsStore[3][394]<=Wgt_3_394;WeightsStore[3][395]<=Wgt_3_395;WeightsStore[3][396]<=Wgt_3_396;WeightsStore[3][397]<=Wgt_3_397;WeightsStore[3][398]<=Wgt_3_398;WeightsStore[3][399]<=Wgt_3_399;WeightsStore[3][400]<=Wgt_3_400;WeightsStore[3][401]<=Wgt_3_401;WeightsStore[3][402]<=Wgt_3_402;WeightsStore[3][403]<=Wgt_3_403;WeightsStore[3][404]<=Wgt_3_404;WeightsStore[3][405]<=Wgt_3_405;WeightsStore[3][406]<=Wgt_3_406;WeightsStore[3][407]<=Wgt_3_407;WeightsStore[3][408]<=Wgt_3_408;WeightsStore[3][409]<=Wgt_3_409;WeightsStore[3][410]<=Wgt_3_410;WeightsStore[3][411]<=Wgt_3_411;WeightsStore[3][412]<=Wgt_3_412;WeightsStore[3][413]<=Wgt_3_413;WeightsStore[3][414]<=Wgt_3_414;WeightsStore[3][415]<=Wgt_3_415;WeightsStore[3][416]<=Wgt_3_416;WeightsStore[3][417]<=Wgt_3_417;WeightsStore[3][418]<=Wgt_3_418;WeightsStore[3][419]<=Wgt_3_419;WeightsStore[3][420]<=Wgt_3_420;WeightsStore[3][421]<=Wgt_3_421;WeightsStore[3][422]<=Wgt_3_422;WeightsStore[3][423]<=Wgt_3_423;WeightsStore[3][424]<=Wgt_3_424;WeightsStore[3][425]<=Wgt_3_425;WeightsStore[3][426]<=Wgt_3_426;WeightsStore[3][427]<=Wgt_3_427;WeightsStore[3][428]<=Wgt_3_428;WeightsStore[3][429]<=Wgt_3_429;WeightsStore[3][430]<=Wgt_3_430;WeightsStore[3][431]<=Wgt_3_431;WeightsStore[3][432]<=Wgt_3_432;WeightsStore[3][433]<=Wgt_3_433;WeightsStore[3][434]<=Wgt_3_434;WeightsStore[3][435]<=Wgt_3_435;WeightsStore[3][436]<=Wgt_3_436;WeightsStore[3][437]<=Wgt_3_437;WeightsStore[3][438]<=Wgt_3_438;WeightsStore[3][439]<=Wgt_3_439;WeightsStore[3][440]<=Wgt_3_440;WeightsStore[3][441]<=Wgt_3_441;WeightsStore[3][442]<=Wgt_3_442;WeightsStore[3][443]<=Wgt_3_443;WeightsStore[3][444]<=Wgt_3_444;WeightsStore[3][445]<=Wgt_3_445;WeightsStore[3][446]<=Wgt_3_446;WeightsStore[3][447]<=Wgt_3_447;WeightsStore[3][448]<=Wgt_3_448;WeightsStore[3][449]<=Wgt_3_449;WeightsStore[3][450]<=Wgt_3_450;WeightsStore[3][451]<=Wgt_3_451;WeightsStore[3][452]<=Wgt_3_452;WeightsStore[3][453]<=Wgt_3_453;WeightsStore[3][454]<=Wgt_3_454;WeightsStore[3][455]<=Wgt_3_455;WeightsStore[3][456]<=Wgt_3_456;WeightsStore[3][457]<=Wgt_3_457;WeightsStore[3][458]<=Wgt_3_458;WeightsStore[3][459]<=Wgt_3_459;WeightsStore[3][460]<=Wgt_3_460;WeightsStore[3][461]<=Wgt_3_461;WeightsStore[3][462]<=Wgt_3_462;WeightsStore[3][463]<=Wgt_3_463;WeightsStore[3][464]<=Wgt_3_464;WeightsStore[3][465]<=Wgt_3_465;WeightsStore[3][466]<=Wgt_3_466;WeightsStore[3][467]<=Wgt_3_467;WeightsStore[3][468]<=Wgt_3_468;WeightsStore[3][469]<=Wgt_3_469;WeightsStore[3][470]<=Wgt_3_470;WeightsStore[3][471]<=Wgt_3_471;WeightsStore[3][472]<=Wgt_3_472;WeightsStore[3][473]<=Wgt_3_473;WeightsStore[3][474]<=Wgt_3_474;WeightsStore[3][475]<=Wgt_3_475;WeightsStore[3][476]<=Wgt_3_476;WeightsStore[3][477]<=Wgt_3_477;WeightsStore[3][478]<=Wgt_3_478;WeightsStore[3][479]<=Wgt_3_479;WeightsStore[3][480]<=Wgt_3_480;WeightsStore[3][481]<=Wgt_3_481;WeightsStore[3][482]<=Wgt_3_482;WeightsStore[3][483]<=Wgt_3_483;WeightsStore[3][484]<=Wgt_3_484;WeightsStore[3][485]<=Wgt_3_485;WeightsStore[3][486]<=Wgt_3_486;WeightsStore[3][487]<=Wgt_3_487;WeightsStore[3][488]<=Wgt_3_488;WeightsStore[3][489]<=Wgt_3_489;WeightsStore[3][490]<=Wgt_3_490;WeightsStore[3][491]<=Wgt_3_491;WeightsStore[3][492]<=Wgt_3_492;WeightsStore[3][493]<=Wgt_3_493;WeightsStore[3][494]<=Wgt_3_494;WeightsStore[3][495]<=Wgt_3_495;WeightsStore[3][496]<=Wgt_3_496;WeightsStore[3][497]<=Wgt_3_497;WeightsStore[3][498]<=Wgt_3_498;WeightsStore[3][499]<=Wgt_3_499;WeightsStore[3][500]<=Wgt_3_500;WeightsStore[3][501]<=Wgt_3_501;WeightsStore[3][502]<=Wgt_3_502;WeightsStore[3][503]<=Wgt_3_503;WeightsStore[3][504]<=Wgt_3_504;WeightsStore[3][505]<=Wgt_3_505;WeightsStore[3][506]<=Wgt_3_506;WeightsStore[3][507]<=Wgt_3_507;WeightsStore[3][508]<=Wgt_3_508;WeightsStore[3][509]<=Wgt_3_509;WeightsStore[3][510]<=Wgt_3_510;WeightsStore[3][511]<=Wgt_3_511;WeightsStore[3][512]<=Wgt_3_512;WeightsStore[3][513]<=Wgt_3_513;WeightsStore[3][514]<=Wgt_3_514;WeightsStore[3][515]<=Wgt_3_515;WeightsStore[3][516]<=Wgt_3_516;WeightsStore[3][517]<=Wgt_3_517;WeightsStore[3][518]<=Wgt_3_518;WeightsStore[3][519]<=Wgt_3_519;WeightsStore[3][520]<=Wgt_3_520;WeightsStore[3][521]<=Wgt_3_521;WeightsStore[3][522]<=Wgt_3_522;WeightsStore[3][523]<=Wgt_3_523;WeightsStore[3][524]<=Wgt_3_524;WeightsStore[3][525]<=Wgt_3_525;WeightsStore[3][526]<=Wgt_3_526;WeightsStore[3][527]<=Wgt_3_527;WeightsStore[3][528]<=Wgt_3_528;WeightsStore[3][529]<=Wgt_3_529;WeightsStore[3][530]<=Wgt_3_530;WeightsStore[3][531]<=Wgt_3_531;WeightsStore[3][532]<=Wgt_3_532;WeightsStore[3][533]<=Wgt_3_533;WeightsStore[3][534]<=Wgt_3_534;WeightsStore[3][535]<=Wgt_3_535;WeightsStore[3][536]<=Wgt_3_536;WeightsStore[3][537]<=Wgt_3_537;WeightsStore[3][538]<=Wgt_3_538;WeightsStore[3][539]<=Wgt_3_539;WeightsStore[3][540]<=Wgt_3_540;WeightsStore[3][541]<=Wgt_3_541;WeightsStore[3][542]<=Wgt_3_542;WeightsStore[3][543]<=Wgt_3_543;WeightsStore[3][544]<=Wgt_3_544;WeightsStore[3][545]<=Wgt_3_545;WeightsStore[3][546]<=Wgt_3_546;WeightsStore[3][547]<=Wgt_3_547;WeightsStore[3][548]<=Wgt_3_548;WeightsStore[3][549]<=Wgt_3_549;WeightsStore[3][550]<=Wgt_3_550;WeightsStore[3][551]<=Wgt_3_551;WeightsStore[3][552]<=Wgt_3_552;WeightsStore[3][553]<=Wgt_3_553;WeightsStore[3][554]<=Wgt_3_554;WeightsStore[3][555]<=Wgt_3_555;WeightsStore[3][556]<=Wgt_3_556;WeightsStore[3][557]<=Wgt_3_557;WeightsStore[3][558]<=Wgt_3_558;WeightsStore[3][559]<=Wgt_3_559;WeightsStore[3][560]<=Wgt_3_560;WeightsStore[3][561]<=Wgt_3_561;WeightsStore[3][562]<=Wgt_3_562;WeightsStore[3][563]<=Wgt_3_563;WeightsStore[3][564]<=Wgt_3_564;WeightsStore[3][565]<=Wgt_3_565;WeightsStore[3][566]<=Wgt_3_566;WeightsStore[3][567]<=Wgt_3_567;WeightsStore[3][568]<=Wgt_3_568;WeightsStore[3][569]<=Wgt_3_569;WeightsStore[3][570]<=Wgt_3_570;WeightsStore[3][571]<=Wgt_3_571;WeightsStore[3][572]<=Wgt_3_572;WeightsStore[3][573]<=Wgt_3_573;WeightsStore[3][574]<=Wgt_3_574;WeightsStore[3][575]<=Wgt_3_575;WeightsStore[3][576]<=Wgt_3_576;WeightsStore[3][577]<=Wgt_3_577;WeightsStore[3][578]<=Wgt_3_578;WeightsStore[3][579]<=Wgt_3_579;WeightsStore[3][580]<=Wgt_3_580;WeightsStore[3][581]<=Wgt_3_581;WeightsStore[3][582]<=Wgt_3_582;WeightsStore[3][583]<=Wgt_3_583;WeightsStore[3][584]<=Wgt_3_584;WeightsStore[3][585]<=Wgt_3_585;WeightsStore[3][586]<=Wgt_3_586;WeightsStore[3][587]<=Wgt_3_587;WeightsStore[3][588]<=Wgt_3_588;WeightsStore[3][589]<=Wgt_3_589;WeightsStore[3][590]<=Wgt_3_590;WeightsStore[3][591]<=Wgt_3_591;WeightsStore[3][592]<=Wgt_3_592;WeightsStore[3][593]<=Wgt_3_593;WeightsStore[3][594]<=Wgt_3_594;WeightsStore[3][595]<=Wgt_3_595;WeightsStore[3][596]<=Wgt_3_596;WeightsStore[3][597]<=Wgt_3_597;WeightsStore[3][598]<=Wgt_3_598;WeightsStore[3][599]<=Wgt_3_599;WeightsStore[3][600]<=Wgt_3_600;WeightsStore[3][601]<=Wgt_3_601;WeightsStore[3][602]<=Wgt_3_602;WeightsStore[3][603]<=Wgt_3_603;WeightsStore[3][604]<=Wgt_3_604;WeightsStore[3][605]<=Wgt_3_605;WeightsStore[3][606]<=Wgt_3_606;WeightsStore[3][607]<=Wgt_3_607;WeightsStore[3][608]<=Wgt_3_608;WeightsStore[3][609]<=Wgt_3_609;WeightsStore[3][610]<=Wgt_3_610;WeightsStore[3][611]<=Wgt_3_611;WeightsStore[3][612]<=Wgt_3_612;WeightsStore[3][613]<=Wgt_3_613;WeightsStore[3][614]<=Wgt_3_614;WeightsStore[3][615]<=Wgt_3_615;WeightsStore[3][616]<=Wgt_3_616;WeightsStore[3][617]<=Wgt_3_617;WeightsStore[3][618]<=Wgt_3_618;WeightsStore[3][619]<=Wgt_3_619;WeightsStore[3][620]<=Wgt_3_620;WeightsStore[3][621]<=Wgt_3_621;WeightsStore[3][622]<=Wgt_3_622;WeightsStore[3][623]<=Wgt_3_623;WeightsStore[3][624]<=Wgt_3_624;WeightsStore[3][625]<=Wgt_3_625;WeightsStore[3][626]<=Wgt_3_626;WeightsStore[3][627]<=Wgt_3_627;WeightsStore[3][628]<=Wgt_3_628;WeightsStore[3][629]<=Wgt_3_629;WeightsStore[3][630]<=Wgt_3_630;WeightsStore[3][631]<=Wgt_3_631;WeightsStore[3][632]<=Wgt_3_632;WeightsStore[3][633]<=Wgt_3_633;WeightsStore[3][634]<=Wgt_3_634;WeightsStore[3][635]<=Wgt_3_635;WeightsStore[3][636]<=Wgt_3_636;WeightsStore[3][637]<=Wgt_3_637;WeightsStore[3][638]<=Wgt_3_638;WeightsStore[3][639]<=Wgt_3_639;WeightsStore[3][640]<=Wgt_3_640;WeightsStore[3][641]<=Wgt_3_641;WeightsStore[3][642]<=Wgt_3_642;WeightsStore[3][643]<=Wgt_3_643;WeightsStore[3][644]<=Wgt_3_644;WeightsStore[3][645]<=Wgt_3_645;WeightsStore[3][646]<=Wgt_3_646;WeightsStore[3][647]<=Wgt_3_647;WeightsStore[3][648]<=Wgt_3_648;WeightsStore[3][649]<=Wgt_3_649;WeightsStore[3][650]<=Wgt_3_650;WeightsStore[3][651]<=Wgt_3_651;WeightsStore[3][652]<=Wgt_3_652;WeightsStore[3][653]<=Wgt_3_653;WeightsStore[3][654]<=Wgt_3_654;WeightsStore[3][655]<=Wgt_3_655;WeightsStore[3][656]<=Wgt_3_656;WeightsStore[3][657]<=Wgt_3_657;WeightsStore[3][658]<=Wgt_3_658;WeightsStore[3][659]<=Wgt_3_659;WeightsStore[3][660]<=Wgt_3_660;WeightsStore[3][661]<=Wgt_3_661;WeightsStore[3][662]<=Wgt_3_662;WeightsStore[3][663]<=Wgt_3_663;WeightsStore[3][664]<=Wgt_3_664;WeightsStore[3][665]<=Wgt_3_665;WeightsStore[3][666]<=Wgt_3_666;WeightsStore[3][667]<=Wgt_3_667;WeightsStore[3][668]<=Wgt_3_668;WeightsStore[3][669]<=Wgt_3_669;WeightsStore[3][670]<=Wgt_3_670;WeightsStore[3][671]<=Wgt_3_671;WeightsStore[3][672]<=Wgt_3_672;WeightsStore[3][673]<=Wgt_3_673;WeightsStore[3][674]<=Wgt_3_674;WeightsStore[3][675]<=Wgt_3_675;WeightsStore[3][676]<=Wgt_3_676;WeightsStore[3][677]<=Wgt_3_677;WeightsStore[3][678]<=Wgt_3_678;WeightsStore[3][679]<=Wgt_3_679;WeightsStore[3][680]<=Wgt_3_680;WeightsStore[3][681]<=Wgt_3_681;WeightsStore[3][682]<=Wgt_3_682;WeightsStore[3][683]<=Wgt_3_683;WeightsStore[3][684]<=Wgt_3_684;WeightsStore[3][685]<=Wgt_3_685;WeightsStore[3][686]<=Wgt_3_686;WeightsStore[3][687]<=Wgt_3_687;WeightsStore[3][688]<=Wgt_3_688;WeightsStore[3][689]<=Wgt_3_689;WeightsStore[3][690]<=Wgt_3_690;WeightsStore[3][691]<=Wgt_3_691;WeightsStore[3][692]<=Wgt_3_692;WeightsStore[3][693]<=Wgt_3_693;WeightsStore[3][694]<=Wgt_3_694;WeightsStore[3][695]<=Wgt_3_695;WeightsStore[3][696]<=Wgt_3_696;WeightsStore[3][697]<=Wgt_3_697;WeightsStore[3][698]<=Wgt_3_698;WeightsStore[3][699]<=Wgt_3_699;WeightsStore[3][700]<=Wgt_3_700;WeightsStore[3][701]<=Wgt_3_701;WeightsStore[3][702]<=Wgt_3_702;WeightsStore[3][703]<=Wgt_3_703;WeightsStore[3][704]<=Wgt_3_704;WeightsStore[3][705]<=Wgt_3_705;WeightsStore[3][706]<=Wgt_3_706;WeightsStore[3][707]<=Wgt_3_707;WeightsStore[3][708]<=Wgt_3_708;WeightsStore[3][709]<=Wgt_3_709;WeightsStore[3][710]<=Wgt_3_710;WeightsStore[3][711]<=Wgt_3_711;WeightsStore[3][712]<=Wgt_3_712;WeightsStore[3][713]<=Wgt_3_713;WeightsStore[3][714]<=Wgt_3_714;WeightsStore[3][715]<=Wgt_3_715;WeightsStore[3][716]<=Wgt_3_716;WeightsStore[3][717]<=Wgt_3_717;WeightsStore[3][718]<=Wgt_3_718;WeightsStore[3][719]<=Wgt_3_719;WeightsStore[3][720]<=Wgt_3_720;WeightsStore[3][721]<=Wgt_3_721;WeightsStore[3][722]<=Wgt_3_722;WeightsStore[3][723]<=Wgt_3_723;WeightsStore[3][724]<=Wgt_3_724;WeightsStore[3][725]<=Wgt_3_725;WeightsStore[3][726]<=Wgt_3_726;WeightsStore[3][727]<=Wgt_3_727;WeightsStore[3][728]<=Wgt_3_728;WeightsStore[3][729]<=Wgt_3_729;WeightsStore[3][730]<=Wgt_3_730;WeightsStore[3][731]<=Wgt_3_731;WeightsStore[3][732]<=Wgt_3_732;WeightsStore[3][733]<=Wgt_3_733;WeightsStore[3][734]<=Wgt_3_734;WeightsStore[3][735]<=Wgt_3_735;WeightsStore[3][736]<=Wgt_3_736;WeightsStore[3][737]<=Wgt_3_737;WeightsStore[3][738]<=Wgt_3_738;WeightsStore[3][739]<=Wgt_3_739;WeightsStore[3][740]<=Wgt_3_740;WeightsStore[3][741]<=Wgt_3_741;WeightsStore[3][742]<=Wgt_3_742;WeightsStore[3][743]<=Wgt_3_743;WeightsStore[3][744]<=Wgt_3_744;WeightsStore[3][745]<=Wgt_3_745;WeightsStore[3][746]<=Wgt_3_746;WeightsStore[3][747]<=Wgt_3_747;WeightsStore[3][748]<=Wgt_3_748;WeightsStore[3][749]<=Wgt_3_749;WeightsStore[3][750]<=Wgt_3_750;WeightsStore[3][751]<=Wgt_3_751;WeightsStore[3][752]<=Wgt_3_752;WeightsStore[3][753]<=Wgt_3_753;WeightsStore[3][754]<=Wgt_3_754;WeightsStore[3][755]<=Wgt_3_755;WeightsStore[3][756]<=Wgt_3_756;WeightsStore[3][757]<=Wgt_3_757;WeightsStore[3][758]<=Wgt_3_758;WeightsStore[3][759]<=Wgt_3_759;WeightsStore[3][760]<=Wgt_3_760;WeightsStore[3][761]<=Wgt_3_761;WeightsStore[3][762]<=Wgt_3_762;WeightsStore[3][763]<=Wgt_3_763;WeightsStore[3][764]<=Wgt_3_764;WeightsStore[3][765]<=Wgt_3_765;WeightsStore[3][766]<=Wgt_3_766;WeightsStore[3][767]<=Wgt_3_767;WeightsStore[3][768]<=Wgt_3_768;WeightsStore[3][769]<=Wgt_3_769;WeightsStore[3][770]<=Wgt_3_770;WeightsStore[3][771]<=Wgt_3_771;WeightsStore[3][772]<=Wgt_3_772;WeightsStore[3][773]<=Wgt_3_773;WeightsStore[3][774]<=Wgt_3_774;WeightsStore[3][775]<=Wgt_3_775;WeightsStore[3][776]<=Wgt_3_776;WeightsStore[3][777]<=Wgt_3_777;WeightsStore[3][778]<=Wgt_3_778;WeightsStore[3][779]<=Wgt_3_779;WeightsStore[3][780]<=Wgt_3_780;WeightsStore[3][781]<=Wgt_3_781;WeightsStore[3][782]<=Wgt_3_782;WeightsStore[3][783]<=Wgt_3_783;WeightsStore[3][784]<=Wgt_3_784;WeightsStore[4][0]<=Wgt_4_0;WeightsStore[4][1]<=Wgt_4_1;WeightsStore[4][2]<=Wgt_4_2;WeightsStore[4][3]<=Wgt_4_3;WeightsStore[4][4]<=Wgt_4_4;WeightsStore[4][5]<=Wgt_4_5;WeightsStore[4][6]<=Wgt_4_6;WeightsStore[4][7]<=Wgt_4_7;WeightsStore[4][8]<=Wgt_4_8;WeightsStore[4][9]<=Wgt_4_9;WeightsStore[4][10]<=Wgt_4_10;WeightsStore[4][11]<=Wgt_4_11;WeightsStore[4][12]<=Wgt_4_12;WeightsStore[4][13]<=Wgt_4_13;WeightsStore[4][14]<=Wgt_4_14;WeightsStore[4][15]<=Wgt_4_15;WeightsStore[4][16]<=Wgt_4_16;WeightsStore[4][17]<=Wgt_4_17;WeightsStore[4][18]<=Wgt_4_18;WeightsStore[4][19]<=Wgt_4_19;WeightsStore[4][20]<=Wgt_4_20;WeightsStore[4][21]<=Wgt_4_21;WeightsStore[4][22]<=Wgt_4_22;WeightsStore[4][23]<=Wgt_4_23;WeightsStore[4][24]<=Wgt_4_24;WeightsStore[4][25]<=Wgt_4_25;WeightsStore[4][26]<=Wgt_4_26;WeightsStore[4][27]<=Wgt_4_27;WeightsStore[4][28]<=Wgt_4_28;WeightsStore[4][29]<=Wgt_4_29;WeightsStore[4][30]<=Wgt_4_30;WeightsStore[4][31]<=Wgt_4_31;WeightsStore[4][32]<=Wgt_4_32;WeightsStore[4][33]<=Wgt_4_33;WeightsStore[4][34]<=Wgt_4_34;WeightsStore[4][35]<=Wgt_4_35;WeightsStore[4][36]<=Wgt_4_36;WeightsStore[4][37]<=Wgt_4_37;WeightsStore[4][38]<=Wgt_4_38;WeightsStore[4][39]<=Wgt_4_39;WeightsStore[4][40]<=Wgt_4_40;WeightsStore[4][41]<=Wgt_4_41;WeightsStore[4][42]<=Wgt_4_42;WeightsStore[4][43]<=Wgt_4_43;WeightsStore[4][44]<=Wgt_4_44;WeightsStore[4][45]<=Wgt_4_45;WeightsStore[4][46]<=Wgt_4_46;WeightsStore[4][47]<=Wgt_4_47;WeightsStore[4][48]<=Wgt_4_48;WeightsStore[4][49]<=Wgt_4_49;WeightsStore[4][50]<=Wgt_4_50;WeightsStore[4][51]<=Wgt_4_51;WeightsStore[4][52]<=Wgt_4_52;WeightsStore[4][53]<=Wgt_4_53;WeightsStore[4][54]<=Wgt_4_54;WeightsStore[4][55]<=Wgt_4_55;WeightsStore[4][56]<=Wgt_4_56;WeightsStore[4][57]<=Wgt_4_57;WeightsStore[4][58]<=Wgt_4_58;WeightsStore[4][59]<=Wgt_4_59;WeightsStore[4][60]<=Wgt_4_60;WeightsStore[4][61]<=Wgt_4_61;WeightsStore[4][62]<=Wgt_4_62;WeightsStore[4][63]<=Wgt_4_63;WeightsStore[4][64]<=Wgt_4_64;WeightsStore[4][65]<=Wgt_4_65;WeightsStore[4][66]<=Wgt_4_66;WeightsStore[4][67]<=Wgt_4_67;WeightsStore[4][68]<=Wgt_4_68;WeightsStore[4][69]<=Wgt_4_69;WeightsStore[4][70]<=Wgt_4_70;WeightsStore[4][71]<=Wgt_4_71;WeightsStore[4][72]<=Wgt_4_72;WeightsStore[4][73]<=Wgt_4_73;WeightsStore[4][74]<=Wgt_4_74;WeightsStore[4][75]<=Wgt_4_75;WeightsStore[4][76]<=Wgt_4_76;WeightsStore[4][77]<=Wgt_4_77;WeightsStore[4][78]<=Wgt_4_78;WeightsStore[4][79]<=Wgt_4_79;WeightsStore[4][80]<=Wgt_4_80;WeightsStore[4][81]<=Wgt_4_81;WeightsStore[4][82]<=Wgt_4_82;WeightsStore[4][83]<=Wgt_4_83;WeightsStore[4][84]<=Wgt_4_84;WeightsStore[4][85]<=Wgt_4_85;WeightsStore[4][86]<=Wgt_4_86;WeightsStore[4][87]<=Wgt_4_87;WeightsStore[4][88]<=Wgt_4_88;WeightsStore[4][89]<=Wgt_4_89;WeightsStore[4][90]<=Wgt_4_90;WeightsStore[4][91]<=Wgt_4_91;WeightsStore[4][92]<=Wgt_4_92;WeightsStore[4][93]<=Wgt_4_93;WeightsStore[4][94]<=Wgt_4_94;WeightsStore[4][95]<=Wgt_4_95;WeightsStore[4][96]<=Wgt_4_96;WeightsStore[4][97]<=Wgt_4_97;WeightsStore[4][98]<=Wgt_4_98;WeightsStore[4][99]<=Wgt_4_99;WeightsStore[4][100]<=Wgt_4_100;WeightsStore[4][101]<=Wgt_4_101;WeightsStore[4][102]<=Wgt_4_102;WeightsStore[4][103]<=Wgt_4_103;WeightsStore[4][104]<=Wgt_4_104;WeightsStore[4][105]<=Wgt_4_105;WeightsStore[4][106]<=Wgt_4_106;WeightsStore[4][107]<=Wgt_4_107;WeightsStore[4][108]<=Wgt_4_108;WeightsStore[4][109]<=Wgt_4_109;WeightsStore[4][110]<=Wgt_4_110;WeightsStore[4][111]<=Wgt_4_111;WeightsStore[4][112]<=Wgt_4_112;WeightsStore[4][113]<=Wgt_4_113;WeightsStore[4][114]<=Wgt_4_114;WeightsStore[4][115]<=Wgt_4_115;WeightsStore[4][116]<=Wgt_4_116;WeightsStore[4][117]<=Wgt_4_117;WeightsStore[4][118]<=Wgt_4_118;WeightsStore[4][119]<=Wgt_4_119;WeightsStore[4][120]<=Wgt_4_120;WeightsStore[4][121]<=Wgt_4_121;WeightsStore[4][122]<=Wgt_4_122;WeightsStore[4][123]<=Wgt_4_123;WeightsStore[4][124]<=Wgt_4_124;WeightsStore[4][125]<=Wgt_4_125;WeightsStore[4][126]<=Wgt_4_126;WeightsStore[4][127]<=Wgt_4_127;WeightsStore[4][128]<=Wgt_4_128;WeightsStore[4][129]<=Wgt_4_129;WeightsStore[4][130]<=Wgt_4_130;WeightsStore[4][131]<=Wgt_4_131;WeightsStore[4][132]<=Wgt_4_132;WeightsStore[4][133]<=Wgt_4_133;WeightsStore[4][134]<=Wgt_4_134;WeightsStore[4][135]<=Wgt_4_135;WeightsStore[4][136]<=Wgt_4_136;WeightsStore[4][137]<=Wgt_4_137;WeightsStore[4][138]<=Wgt_4_138;WeightsStore[4][139]<=Wgt_4_139;WeightsStore[4][140]<=Wgt_4_140;WeightsStore[4][141]<=Wgt_4_141;WeightsStore[4][142]<=Wgt_4_142;WeightsStore[4][143]<=Wgt_4_143;WeightsStore[4][144]<=Wgt_4_144;WeightsStore[4][145]<=Wgt_4_145;WeightsStore[4][146]<=Wgt_4_146;WeightsStore[4][147]<=Wgt_4_147;WeightsStore[4][148]<=Wgt_4_148;WeightsStore[4][149]<=Wgt_4_149;WeightsStore[4][150]<=Wgt_4_150;WeightsStore[4][151]<=Wgt_4_151;WeightsStore[4][152]<=Wgt_4_152;WeightsStore[4][153]<=Wgt_4_153;WeightsStore[4][154]<=Wgt_4_154;WeightsStore[4][155]<=Wgt_4_155;WeightsStore[4][156]<=Wgt_4_156;WeightsStore[4][157]<=Wgt_4_157;WeightsStore[4][158]<=Wgt_4_158;WeightsStore[4][159]<=Wgt_4_159;WeightsStore[4][160]<=Wgt_4_160;WeightsStore[4][161]<=Wgt_4_161;WeightsStore[4][162]<=Wgt_4_162;WeightsStore[4][163]<=Wgt_4_163;WeightsStore[4][164]<=Wgt_4_164;WeightsStore[4][165]<=Wgt_4_165;WeightsStore[4][166]<=Wgt_4_166;WeightsStore[4][167]<=Wgt_4_167;WeightsStore[4][168]<=Wgt_4_168;WeightsStore[4][169]<=Wgt_4_169;WeightsStore[4][170]<=Wgt_4_170;WeightsStore[4][171]<=Wgt_4_171;WeightsStore[4][172]<=Wgt_4_172;WeightsStore[4][173]<=Wgt_4_173;WeightsStore[4][174]<=Wgt_4_174;WeightsStore[4][175]<=Wgt_4_175;WeightsStore[4][176]<=Wgt_4_176;WeightsStore[4][177]<=Wgt_4_177;WeightsStore[4][178]<=Wgt_4_178;WeightsStore[4][179]<=Wgt_4_179;WeightsStore[4][180]<=Wgt_4_180;WeightsStore[4][181]<=Wgt_4_181;WeightsStore[4][182]<=Wgt_4_182;WeightsStore[4][183]<=Wgt_4_183;WeightsStore[4][184]<=Wgt_4_184;WeightsStore[4][185]<=Wgt_4_185;WeightsStore[4][186]<=Wgt_4_186;WeightsStore[4][187]<=Wgt_4_187;WeightsStore[4][188]<=Wgt_4_188;WeightsStore[4][189]<=Wgt_4_189;WeightsStore[4][190]<=Wgt_4_190;WeightsStore[4][191]<=Wgt_4_191;WeightsStore[4][192]<=Wgt_4_192;WeightsStore[4][193]<=Wgt_4_193;WeightsStore[4][194]<=Wgt_4_194;WeightsStore[4][195]<=Wgt_4_195;WeightsStore[4][196]<=Wgt_4_196;WeightsStore[4][197]<=Wgt_4_197;WeightsStore[4][198]<=Wgt_4_198;WeightsStore[4][199]<=Wgt_4_199;WeightsStore[4][200]<=Wgt_4_200;WeightsStore[4][201]<=Wgt_4_201;WeightsStore[4][202]<=Wgt_4_202;WeightsStore[4][203]<=Wgt_4_203;WeightsStore[4][204]<=Wgt_4_204;WeightsStore[4][205]<=Wgt_4_205;WeightsStore[4][206]<=Wgt_4_206;WeightsStore[4][207]<=Wgt_4_207;WeightsStore[4][208]<=Wgt_4_208;WeightsStore[4][209]<=Wgt_4_209;WeightsStore[4][210]<=Wgt_4_210;WeightsStore[4][211]<=Wgt_4_211;WeightsStore[4][212]<=Wgt_4_212;WeightsStore[4][213]<=Wgt_4_213;WeightsStore[4][214]<=Wgt_4_214;WeightsStore[4][215]<=Wgt_4_215;WeightsStore[4][216]<=Wgt_4_216;WeightsStore[4][217]<=Wgt_4_217;WeightsStore[4][218]<=Wgt_4_218;WeightsStore[4][219]<=Wgt_4_219;WeightsStore[4][220]<=Wgt_4_220;WeightsStore[4][221]<=Wgt_4_221;WeightsStore[4][222]<=Wgt_4_222;WeightsStore[4][223]<=Wgt_4_223;WeightsStore[4][224]<=Wgt_4_224;WeightsStore[4][225]<=Wgt_4_225;WeightsStore[4][226]<=Wgt_4_226;WeightsStore[4][227]<=Wgt_4_227;WeightsStore[4][228]<=Wgt_4_228;WeightsStore[4][229]<=Wgt_4_229;WeightsStore[4][230]<=Wgt_4_230;WeightsStore[4][231]<=Wgt_4_231;WeightsStore[4][232]<=Wgt_4_232;WeightsStore[4][233]<=Wgt_4_233;WeightsStore[4][234]<=Wgt_4_234;WeightsStore[4][235]<=Wgt_4_235;WeightsStore[4][236]<=Wgt_4_236;WeightsStore[4][237]<=Wgt_4_237;WeightsStore[4][238]<=Wgt_4_238;WeightsStore[4][239]<=Wgt_4_239;WeightsStore[4][240]<=Wgt_4_240;WeightsStore[4][241]<=Wgt_4_241;WeightsStore[4][242]<=Wgt_4_242;WeightsStore[4][243]<=Wgt_4_243;WeightsStore[4][244]<=Wgt_4_244;WeightsStore[4][245]<=Wgt_4_245;WeightsStore[4][246]<=Wgt_4_246;WeightsStore[4][247]<=Wgt_4_247;WeightsStore[4][248]<=Wgt_4_248;WeightsStore[4][249]<=Wgt_4_249;WeightsStore[4][250]<=Wgt_4_250;WeightsStore[4][251]<=Wgt_4_251;WeightsStore[4][252]<=Wgt_4_252;WeightsStore[4][253]<=Wgt_4_253;WeightsStore[4][254]<=Wgt_4_254;WeightsStore[4][255]<=Wgt_4_255;WeightsStore[4][256]<=Wgt_4_256;WeightsStore[4][257]<=Wgt_4_257;WeightsStore[4][258]<=Wgt_4_258;WeightsStore[4][259]<=Wgt_4_259;WeightsStore[4][260]<=Wgt_4_260;WeightsStore[4][261]<=Wgt_4_261;WeightsStore[4][262]<=Wgt_4_262;WeightsStore[4][263]<=Wgt_4_263;WeightsStore[4][264]<=Wgt_4_264;WeightsStore[4][265]<=Wgt_4_265;WeightsStore[4][266]<=Wgt_4_266;WeightsStore[4][267]<=Wgt_4_267;WeightsStore[4][268]<=Wgt_4_268;WeightsStore[4][269]<=Wgt_4_269;WeightsStore[4][270]<=Wgt_4_270;WeightsStore[4][271]<=Wgt_4_271;WeightsStore[4][272]<=Wgt_4_272;WeightsStore[4][273]<=Wgt_4_273;WeightsStore[4][274]<=Wgt_4_274;WeightsStore[4][275]<=Wgt_4_275;WeightsStore[4][276]<=Wgt_4_276;WeightsStore[4][277]<=Wgt_4_277;WeightsStore[4][278]<=Wgt_4_278;WeightsStore[4][279]<=Wgt_4_279;WeightsStore[4][280]<=Wgt_4_280;WeightsStore[4][281]<=Wgt_4_281;WeightsStore[4][282]<=Wgt_4_282;WeightsStore[4][283]<=Wgt_4_283;WeightsStore[4][284]<=Wgt_4_284;WeightsStore[4][285]<=Wgt_4_285;WeightsStore[4][286]<=Wgt_4_286;WeightsStore[4][287]<=Wgt_4_287;WeightsStore[4][288]<=Wgt_4_288;WeightsStore[4][289]<=Wgt_4_289;WeightsStore[4][290]<=Wgt_4_290;WeightsStore[4][291]<=Wgt_4_291;WeightsStore[4][292]<=Wgt_4_292;WeightsStore[4][293]<=Wgt_4_293;WeightsStore[4][294]<=Wgt_4_294;WeightsStore[4][295]<=Wgt_4_295;WeightsStore[4][296]<=Wgt_4_296;WeightsStore[4][297]<=Wgt_4_297;WeightsStore[4][298]<=Wgt_4_298;WeightsStore[4][299]<=Wgt_4_299;WeightsStore[4][300]<=Wgt_4_300;WeightsStore[4][301]<=Wgt_4_301;WeightsStore[4][302]<=Wgt_4_302;WeightsStore[4][303]<=Wgt_4_303;WeightsStore[4][304]<=Wgt_4_304;WeightsStore[4][305]<=Wgt_4_305;WeightsStore[4][306]<=Wgt_4_306;WeightsStore[4][307]<=Wgt_4_307;WeightsStore[4][308]<=Wgt_4_308;WeightsStore[4][309]<=Wgt_4_309;WeightsStore[4][310]<=Wgt_4_310;WeightsStore[4][311]<=Wgt_4_311;WeightsStore[4][312]<=Wgt_4_312;WeightsStore[4][313]<=Wgt_4_313;WeightsStore[4][314]<=Wgt_4_314;WeightsStore[4][315]<=Wgt_4_315;WeightsStore[4][316]<=Wgt_4_316;WeightsStore[4][317]<=Wgt_4_317;WeightsStore[4][318]<=Wgt_4_318;WeightsStore[4][319]<=Wgt_4_319;WeightsStore[4][320]<=Wgt_4_320;WeightsStore[4][321]<=Wgt_4_321;WeightsStore[4][322]<=Wgt_4_322;WeightsStore[4][323]<=Wgt_4_323;WeightsStore[4][324]<=Wgt_4_324;WeightsStore[4][325]<=Wgt_4_325;WeightsStore[4][326]<=Wgt_4_326;WeightsStore[4][327]<=Wgt_4_327;WeightsStore[4][328]<=Wgt_4_328;WeightsStore[4][329]<=Wgt_4_329;WeightsStore[4][330]<=Wgt_4_330;WeightsStore[4][331]<=Wgt_4_331;WeightsStore[4][332]<=Wgt_4_332;WeightsStore[4][333]<=Wgt_4_333;WeightsStore[4][334]<=Wgt_4_334;WeightsStore[4][335]<=Wgt_4_335;WeightsStore[4][336]<=Wgt_4_336;WeightsStore[4][337]<=Wgt_4_337;WeightsStore[4][338]<=Wgt_4_338;WeightsStore[4][339]<=Wgt_4_339;WeightsStore[4][340]<=Wgt_4_340;WeightsStore[4][341]<=Wgt_4_341;WeightsStore[4][342]<=Wgt_4_342;WeightsStore[4][343]<=Wgt_4_343;WeightsStore[4][344]<=Wgt_4_344;WeightsStore[4][345]<=Wgt_4_345;WeightsStore[4][346]<=Wgt_4_346;WeightsStore[4][347]<=Wgt_4_347;WeightsStore[4][348]<=Wgt_4_348;WeightsStore[4][349]<=Wgt_4_349;WeightsStore[4][350]<=Wgt_4_350;WeightsStore[4][351]<=Wgt_4_351;WeightsStore[4][352]<=Wgt_4_352;WeightsStore[4][353]<=Wgt_4_353;WeightsStore[4][354]<=Wgt_4_354;WeightsStore[4][355]<=Wgt_4_355;WeightsStore[4][356]<=Wgt_4_356;WeightsStore[4][357]<=Wgt_4_357;WeightsStore[4][358]<=Wgt_4_358;WeightsStore[4][359]<=Wgt_4_359;WeightsStore[4][360]<=Wgt_4_360;WeightsStore[4][361]<=Wgt_4_361;WeightsStore[4][362]<=Wgt_4_362;WeightsStore[4][363]<=Wgt_4_363;WeightsStore[4][364]<=Wgt_4_364;WeightsStore[4][365]<=Wgt_4_365;WeightsStore[4][366]<=Wgt_4_366;WeightsStore[4][367]<=Wgt_4_367;WeightsStore[4][368]<=Wgt_4_368;WeightsStore[4][369]<=Wgt_4_369;WeightsStore[4][370]<=Wgt_4_370;WeightsStore[4][371]<=Wgt_4_371;WeightsStore[4][372]<=Wgt_4_372;WeightsStore[4][373]<=Wgt_4_373;WeightsStore[4][374]<=Wgt_4_374;WeightsStore[4][375]<=Wgt_4_375;WeightsStore[4][376]<=Wgt_4_376;WeightsStore[4][377]<=Wgt_4_377;WeightsStore[4][378]<=Wgt_4_378;WeightsStore[4][379]<=Wgt_4_379;WeightsStore[4][380]<=Wgt_4_380;WeightsStore[4][381]<=Wgt_4_381;WeightsStore[4][382]<=Wgt_4_382;WeightsStore[4][383]<=Wgt_4_383;WeightsStore[4][384]<=Wgt_4_384;WeightsStore[4][385]<=Wgt_4_385;WeightsStore[4][386]<=Wgt_4_386;WeightsStore[4][387]<=Wgt_4_387;WeightsStore[4][388]<=Wgt_4_388;WeightsStore[4][389]<=Wgt_4_389;WeightsStore[4][390]<=Wgt_4_390;WeightsStore[4][391]<=Wgt_4_391;WeightsStore[4][392]<=Wgt_4_392;WeightsStore[4][393]<=Wgt_4_393;WeightsStore[4][394]<=Wgt_4_394;WeightsStore[4][395]<=Wgt_4_395;WeightsStore[4][396]<=Wgt_4_396;WeightsStore[4][397]<=Wgt_4_397;WeightsStore[4][398]<=Wgt_4_398;WeightsStore[4][399]<=Wgt_4_399;WeightsStore[4][400]<=Wgt_4_400;WeightsStore[4][401]<=Wgt_4_401;WeightsStore[4][402]<=Wgt_4_402;WeightsStore[4][403]<=Wgt_4_403;WeightsStore[4][404]<=Wgt_4_404;WeightsStore[4][405]<=Wgt_4_405;WeightsStore[4][406]<=Wgt_4_406;WeightsStore[4][407]<=Wgt_4_407;WeightsStore[4][408]<=Wgt_4_408;WeightsStore[4][409]<=Wgt_4_409;WeightsStore[4][410]<=Wgt_4_410;WeightsStore[4][411]<=Wgt_4_411;WeightsStore[4][412]<=Wgt_4_412;WeightsStore[4][413]<=Wgt_4_413;WeightsStore[4][414]<=Wgt_4_414;WeightsStore[4][415]<=Wgt_4_415;WeightsStore[4][416]<=Wgt_4_416;WeightsStore[4][417]<=Wgt_4_417;WeightsStore[4][418]<=Wgt_4_418;WeightsStore[4][419]<=Wgt_4_419;WeightsStore[4][420]<=Wgt_4_420;WeightsStore[4][421]<=Wgt_4_421;WeightsStore[4][422]<=Wgt_4_422;WeightsStore[4][423]<=Wgt_4_423;WeightsStore[4][424]<=Wgt_4_424;WeightsStore[4][425]<=Wgt_4_425;WeightsStore[4][426]<=Wgt_4_426;WeightsStore[4][427]<=Wgt_4_427;WeightsStore[4][428]<=Wgt_4_428;WeightsStore[4][429]<=Wgt_4_429;WeightsStore[4][430]<=Wgt_4_430;WeightsStore[4][431]<=Wgt_4_431;WeightsStore[4][432]<=Wgt_4_432;WeightsStore[4][433]<=Wgt_4_433;WeightsStore[4][434]<=Wgt_4_434;WeightsStore[4][435]<=Wgt_4_435;WeightsStore[4][436]<=Wgt_4_436;WeightsStore[4][437]<=Wgt_4_437;WeightsStore[4][438]<=Wgt_4_438;WeightsStore[4][439]<=Wgt_4_439;WeightsStore[4][440]<=Wgt_4_440;WeightsStore[4][441]<=Wgt_4_441;WeightsStore[4][442]<=Wgt_4_442;WeightsStore[4][443]<=Wgt_4_443;WeightsStore[4][444]<=Wgt_4_444;WeightsStore[4][445]<=Wgt_4_445;WeightsStore[4][446]<=Wgt_4_446;WeightsStore[4][447]<=Wgt_4_447;WeightsStore[4][448]<=Wgt_4_448;WeightsStore[4][449]<=Wgt_4_449;WeightsStore[4][450]<=Wgt_4_450;WeightsStore[4][451]<=Wgt_4_451;WeightsStore[4][452]<=Wgt_4_452;WeightsStore[4][453]<=Wgt_4_453;WeightsStore[4][454]<=Wgt_4_454;WeightsStore[4][455]<=Wgt_4_455;WeightsStore[4][456]<=Wgt_4_456;WeightsStore[4][457]<=Wgt_4_457;WeightsStore[4][458]<=Wgt_4_458;WeightsStore[4][459]<=Wgt_4_459;WeightsStore[4][460]<=Wgt_4_460;WeightsStore[4][461]<=Wgt_4_461;WeightsStore[4][462]<=Wgt_4_462;WeightsStore[4][463]<=Wgt_4_463;WeightsStore[4][464]<=Wgt_4_464;WeightsStore[4][465]<=Wgt_4_465;WeightsStore[4][466]<=Wgt_4_466;WeightsStore[4][467]<=Wgt_4_467;WeightsStore[4][468]<=Wgt_4_468;WeightsStore[4][469]<=Wgt_4_469;WeightsStore[4][470]<=Wgt_4_470;WeightsStore[4][471]<=Wgt_4_471;WeightsStore[4][472]<=Wgt_4_472;WeightsStore[4][473]<=Wgt_4_473;WeightsStore[4][474]<=Wgt_4_474;WeightsStore[4][475]<=Wgt_4_475;WeightsStore[4][476]<=Wgt_4_476;WeightsStore[4][477]<=Wgt_4_477;WeightsStore[4][478]<=Wgt_4_478;WeightsStore[4][479]<=Wgt_4_479;WeightsStore[4][480]<=Wgt_4_480;WeightsStore[4][481]<=Wgt_4_481;WeightsStore[4][482]<=Wgt_4_482;WeightsStore[4][483]<=Wgt_4_483;WeightsStore[4][484]<=Wgt_4_484;WeightsStore[4][485]<=Wgt_4_485;WeightsStore[4][486]<=Wgt_4_486;WeightsStore[4][487]<=Wgt_4_487;WeightsStore[4][488]<=Wgt_4_488;WeightsStore[4][489]<=Wgt_4_489;WeightsStore[4][490]<=Wgt_4_490;WeightsStore[4][491]<=Wgt_4_491;WeightsStore[4][492]<=Wgt_4_492;WeightsStore[4][493]<=Wgt_4_493;WeightsStore[4][494]<=Wgt_4_494;WeightsStore[4][495]<=Wgt_4_495;WeightsStore[4][496]<=Wgt_4_496;WeightsStore[4][497]<=Wgt_4_497;WeightsStore[4][498]<=Wgt_4_498;WeightsStore[4][499]<=Wgt_4_499;WeightsStore[4][500]<=Wgt_4_500;WeightsStore[4][501]<=Wgt_4_501;WeightsStore[4][502]<=Wgt_4_502;WeightsStore[4][503]<=Wgt_4_503;WeightsStore[4][504]<=Wgt_4_504;WeightsStore[4][505]<=Wgt_4_505;WeightsStore[4][506]<=Wgt_4_506;WeightsStore[4][507]<=Wgt_4_507;WeightsStore[4][508]<=Wgt_4_508;WeightsStore[4][509]<=Wgt_4_509;WeightsStore[4][510]<=Wgt_4_510;WeightsStore[4][511]<=Wgt_4_511;WeightsStore[4][512]<=Wgt_4_512;WeightsStore[4][513]<=Wgt_4_513;WeightsStore[4][514]<=Wgt_4_514;WeightsStore[4][515]<=Wgt_4_515;WeightsStore[4][516]<=Wgt_4_516;WeightsStore[4][517]<=Wgt_4_517;WeightsStore[4][518]<=Wgt_4_518;WeightsStore[4][519]<=Wgt_4_519;WeightsStore[4][520]<=Wgt_4_520;WeightsStore[4][521]<=Wgt_4_521;WeightsStore[4][522]<=Wgt_4_522;WeightsStore[4][523]<=Wgt_4_523;WeightsStore[4][524]<=Wgt_4_524;WeightsStore[4][525]<=Wgt_4_525;WeightsStore[4][526]<=Wgt_4_526;WeightsStore[4][527]<=Wgt_4_527;WeightsStore[4][528]<=Wgt_4_528;WeightsStore[4][529]<=Wgt_4_529;WeightsStore[4][530]<=Wgt_4_530;WeightsStore[4][531]<=Wgt_4_531;WeightsStore[4][532]<=Wgt_4_532;WeightsStore[4][533]<=Wgt_4_533;WeightsStore[4][534]<=Wgt_4_534;WeightsStore[4][535]<=Wgt_4_535;WeightsStore[4][536]<=Wgt_4_536;WeightsStore[4][537]<=Wgt_4_537;WeightsStore[4][538]<=Wgt_4_538;WeightsStore[4][539]<=Wgt_4_539;WeightsStore[4][540]<=Wgt_4_540;WeightsStore[4][541]<=Wgt_4_541;WeightsStore[4][542]<=Wgt_4_542;WeightsStore[4][543]<=Wgt_4_543;WeightsStore[4][544]<=Wgt_4_544;WeightsStore[4][545]<=Wgt_4_545;WeightsStore[4][546]<=Wgt_4_546;WeightsStore[4][547]<=Wgt_4_547;WeightsStore[4][548]<=Wgt_4_548;WeightsStore[4][549]<=Wgt_4_549;WeightsStore[4][550]<=Wgt_4_550;WeightsStore[4][551]<=Wgt_4_551;WeightsStore[4][552]<=Wgt_4_552;WeightsStore[4][553]<=Wgt_4_553;WeightsStore[4][554]<=Wgt_4_554;WeightsStore[4][555]<=Wgt_4_555;WeightsStore[4][556]<=Wgt_4_556;WeightsStore[4][557]<=Wgt_4_557;WeightsStore[4][558]<=Wgt_4_558;WeightsStore[4][559]<=Wgt_4_559;WeightsStore[4][560]<=Wgt_4_560;WeightsStore[4][561]<=Wgt_4_561;WeightsStore[4][562]<=Wgt_4_562;WeightsStore[4][563]<=Wgt_4_563;WeightsStore[4][564]<=Wgt_4_564;WeightsStore[4][565]<=Wgt_4_565;WeightsStore[4][566]<=Wgt_4_566;WeightsStore[4][567]<=Wgt_4_567;WeightsStore[4][568]<=Wgt_4_568;WeightsStore[4][569]<=Wgt_4_569;WeightsStore[4][570]<=Wgt_4_570;WeightsStore[4][571]<=Wgt_4_571;WeightsStore[4][572]<=Wgt_4_572;WeightsStore[4][573]<=Wgt_4_573;WeightsStore[4][574]<=Wgt_4_574;WeightsStore[4][575]<=Wgt_4_575;WeightsStore[4][576]<=Wgt_4_576;WeightsStore[4][577]<=Wgt_4_577;WeightsStore[4][578]<=Wgt_4_578;WeightsStore[4][579]<=Wgt_4_579;WeightsStore[4][580]<=Wgt_4_580;WeightsStore[4][581]<=Wgt_4_581;WeightsStore[4][582]<=Wgt_4_582;WeightsStore[4][583]<=Wgt_4_583;WeightsStore[4][584]<=Wgt_4_584;WeightsStore[4][585]<=Wgt_4_585;WeightsStore[4][586]<=Wgt_4_586;WeightsStore[4][587]<=Wgt_4_587;WeightsStore[4][588]<=Wgt_4_588;WeightsStore[4][589]<=Wgt_4_589;WeightsStore[4][590]<=Wgt_4_590;WeightsStore[4][591]<=Wgt_4_591;WeightsStore[4][592]<=Wgt_4_592;WeightsStore[4][593]<=Wgt_4_593;WeightsStore[4][594]<=Wgt_4_594;WeightsStore[4][595]<=Wgt_4_595;WeightsStore[4][596]<=Wgt_4_596;WeightsStore[4][597]<=Wgt_4_597;WeightsStore[4][598]<=Wgt_4_598;WeightsStore[4][599]<=Wgt_4_599;WeightsStore[4][600]<=Wgt_4_600;WeightsStore[4][601]<=Wgt_4_601;WeightsStore[4][602]<=Wgt_4_602;WeightsStore[4][603]<=Wgt_4_603;WeightsStore[4][604]<=Wgt_4_604;WeightsStore[4][605]<=Wgt_4_605;WeightsStore[4][606]<=Wgt_4_606;WeightsStore[4][607]<=Wgt_4_607;WeightsStore[4][608]<=Wgt_4_608;WeightsStore[4][609]<=Wgt_4_609;WeightsStore[4][610]<=Wgt_4_610;WeightsStore[4][611]<=Wgt_4_611;WeightsStore[4][612]<=Wgt_4_612;WeightsStore[4][613]<=Wgt_4_613;WeightsStore[4][614]<=Wgt_4_614;WeightsStore[4][615]<=Wgt_4_615;WeightsStore[4][616]<=Wgt_4_616;WeightsStore[4][617]<=Wgt_4_617;WeightsStore[4][618]<=Wgt_4_618;WeightsStore[4][619]<=Wgt_4_619;WeightsStore[4][620]<=Wgt_4_620;WeightsStore[4][621]<=Wgt_4_621;WeightsStore[4][622]<=Wgt_4_622;WeightsStore[4][623]<=Wgt_4_623;WeightsStore[4][624]<=Wgt_4_624;WeightsStore[4][625]<=Wgt_4_625;WeightsStore[4][626]<=Wgt_4_626;WeightsStore[4][627]<=Wgt_4_627;WeightsStore[4][628]<=Wgt_4_628;WeightsStore[4][629]<=Wgt_4_629;WeightsStore[4][630]<=Wgt_4_630;WeightsStore[4][631]<=Wgt_4_631;WeightsStore[4][632]<=Wgt_4_632;WeightsStore[4][633]<=Wgt_4_633;WeightsStore[4][634]<=Wgt_4_634;WeightsStore[4][635]<=Wgt_4_635;WeightsStore[4][636]<=Wgt_4_636;WeightsStore[4][637]<=Wgt_4_637;WeightsStore[4][638]<=Wgt_4_638;WeightsStore[4][639]<=Wgt_4_639;WeightsStore[4][640]<=Wgt_4_640;WeightsStore[4][641]<=Wgt_4_641;WeightsStore[4][642]<=Wgt_4_642;WeightsStore[4][643]<=Wgt_4_643;WeightsStore[4][644]<=Wgt_4_644;WeightsStore[4][645]<=Wgt_4_645;WeightsStore[4][646]<=Wgt_4_646;WeightsStore[4][647]<=Wgt_4_647;WeightsStore[4][648]<=Wgt_4_648;WeightsStore[4][649]<=Wgt_4_649;WeightsStore[4][650]<=Wgt_4_650;WeightsStore[4][651]<=Wgt_4_651;WeightsStore[4][652]<=Wgt_4_652;WeightsStore[4][653]<=Wgt_4_653;WeightsStore[4][654]<=Wgt_4_654;WeightsStore[4][655]<=Wgt_4_655;WeightsStore[4][656]<=Wgt_4_656;WeightsStore[4][657]<=Wgt_4_657;WeightsStore[4][658]<=Wgt_4_658;WeightsStore[4][659]<=Wgt_4_659;WeightsStore[4][660]<=Wgt_4_660;WeightsStore[4][661]<=Wgt_4_661;WeightsStore[4][662]<=Wgt_4_662;WeightsStore[4][663]<=Wgt_4_663;WeightsStore[4][664]<=Wgt_4_664;WeightsStore[4][665]<=Wgt_4_665;WeightsStore[4][666]<=Wgt_4_666;WeightsStore[4][667]<=Wgt_4_667;WeightsStore[4][668]<=Wgt_4_668;WeightsStore[4][669]<=Wgt_4_669;WeightsStore[4][670]<=Wgt_4_670;WeightsStore[4][671]<=Wgt_4_671;WeightsStore[4][672]<=Wgt_4_672;WeightsStore[4][673]<=Wgt_4_673;WeightsStore[4][674]<=Wgt_4_674;WeightsStore[4][675]<=Wgt_4_675;WeightsStore[4][676]<=Wgt_4_676;WeightsStore[4][677]<=Wgt_4_677;WeightsStore[4][678]<=Wgt_4_678;WeightsStore[4][679]<=Wgt_4_679;WeightsStore[4][680]<=Wgt_4_680;WeightsStore[4][681]<=Wgt_4_681;WeightsStore[4][682]<=Wgt_4_682;WeightsStore[4][683]<=Wgt_4_683;WeightsStore[4][684]<=Wgt_4_684;WeightsStore[4][685]<=Wgt_4_685;WeightsStore[4][686]<=Wgt_4_686;WeightsStore[4][687]<=Wgt_4_687;WeightsStore[4][688]<=Wgt_4_688;WeightsStore[4][689]<=Wgt_4_689;WeightsStore[4][690]<=Wgt_4_690;WeightsStore[4][691]<=Wgt_4_691;WeightsStore[4][692]<=Wgt_4_692;WeightsStore[4][693]<=Wgt_4_693;WeightsStore[4][694]<=Wgt_4_694;WeightsStore[4][695]<=Wgt_4_695;WeightsStore[4][696]<=Wgt_4_696;WeightsStore[4][697]<=Wgt_4_697;WeightsStore[4][698]<=Wgt_4_698;WeightsStore[4][699]<=Wgt_4_699;WeightsStore[4][700]<=Wgt_4_700;WeightsStore[4][701]<=Wgt_4_701;WeightsStore[4][702]<=Wgt_4_702;WeightsStore[4][703]<=Wgt_4_703;WeightsStore[4][704]<=Wgt_4_704;WeightsStore[4][705]<=Wgt_4_705;WeightsStore[4][706]<=Wgt_4_706;WeightsStore[4][707]<=Wgt_4_707;WeightsStore[4][708]<=Wgt_4_708;WeightsStore[4][709]<=Wgt_4_709;WeightsStore[4][710]<=Wgt_4_710;WeightsStore[4][711]<=Wgt_4_711;WeightsStore[4][712]<=Wgt_4_712;WeightsStore[4][713]<=Wgt_4_713;WeightsStore[4][714]<=Wgt_4_714;WeightsStore[4][715]<=Wgt_4_715;WeightsStore[4][716]<=Wgt_4_716;WeightsStore[4][717]<=Wgt_4_717;WeightsStore[4][718]<=Wgt_4_718;WeightsStore[4][719]<=Wgt_4_719;WeightsStore[4][720]<=Wgt_4_720;WeightsStore[4][721]<=Wgt_4_721;WeightsStore[4][722]<=Wgt_4_722;WeightsStore[4][723]<=Wgt_4_723;WeightsStore[4][724]<=Wgt_4_724;WeightsStore[4][725]<=Wgt_4_725;WeightsStore[4][726]<=Wgt_4_726;WeightsStore[4][727]<=Wgt_4_727;WeightsStore[4][728]<=Wgt_4_728;WeightsStore[4][729]<=Wgt_4_729;WeightsStore[4][730]<=Wgt_4_730;WeightsStore[4][731]<=Wgt_4_731;WeightsStore[4][732]<=Wgt_4_732;WeightsStore[4][733]<=Wgt_4_733;WeightsStore[4][734]<=Wgt_4_734;WeightsStore[4][735]<=Wgt_4_735;WeightsStore[4][736]<=Wgt_4_736;WeightsStore[4][737]<=Wgt_4_737;WeightsStore[4][738]<=Wgt_4_738;WeightsStore[4][739]<=Wgt_4_739;WeightsStore[4][740]<=Wgt_4_740;WeightsStore[4][741]<=Wgt_4_741;WeightsStore[4][742]<=Wgt_4_742;WeightsStore[4][743]<=Wgt_4_743;WeightsStore[4][744]<=Wgt_4_744;WeightsStore[4][745]<=Wgt_4_745;WeightsStore[4][746]<=Wgt_4_746;WeightsStore[4][747]<=Wgt_4_747;WeightsStore[4][748]<=Wgt_4_748;WeightsStore[4][749]<=Wgt_4_749;WeightsStore[4][750]<=Wgt_4_750;WeightsStore[4][751]<=Wgt_4_751;WeightsStore[4][752]<=Wgt_4_752;WeightsStore[4][753]<=Wgt_4_753;WeightsStore[4][754]<=Wgt_4_754;WeightsStore[4][755]<=Wgt_4_755;WeightsStore[4][756]<=Wgt_4_756;WeightsStore[4][757]<=Wgt_4_757;WeightsStore[4][758]<=Wgt_4_758;WeightsStore[4][759]<=Wgt_4_759;WeightsStore[4][760]<=Wgt_4_760;WeightsStore[4][761]<=Wgt_4_761;WeightsStore[4][762]<=Wgt_4_762;WeightsStore[4][763]<=Wgt_4_763;WeightsStore[4][764]<=Wgt_4_764;WeightsStore[4][765]<=Wgt_4_765;WeightsStore[4][766]<=Wgt_4_766;WeightsStore[4][767]<=Wgt_4_767;WeightsStore[4][768]<=Wgt_4_768;WeightsStore[4][769]<=Wgt_4_769;WeightsStore[4][770]<=Wgt_4_770;WeightsStore[4][771]<=Wgt_4_771;WeightsStore[4][772]<=Wgt_4_772;WeightsStore[4][773]<=Wgt_4_773;WeightsStore[4][774]<=Wgt_4_774;WeightsStore[4][775]<=Wgt_4_775;WeightsStore[4][776]<=Wgt_4_776;WeightsStore[4][777]<=Wgt_4_777;WeightsStore[4][778]<=Wgt_4_778;WeightsStore[4][779]<=Wgt_4_779;WeightsStore[4][780]<=Wgt_4_780;WeightsStore[4][781]<=Wgt_4_781;WeightsStore[4][782]<=Wgt_4_782;WeightsStore[4][783]<=Wgt_4_783;WeightsStore[4][784]<=Wgt_4_784;WeightsStore[5][0]<=Wgt_5_0;WeightsStore[5][1]<=Wgt_5_1;WeightsStore[5][2]<=Wgt_5_2;WeightsStore[5][3]<=Wgt_5_3;WeightsStore[5][4]<=Wgt_5_4;WeightsStore[5][5]<=Wgt_5_5;WeightsStore[5][6]<=Wgt_5_6;WeightsStore[5][7]<=Wgt_5_7;WeightsStore[5][8]<=Wgt_5_8;WeightsStore[5][9]<=Wgt_5_9;WeightsStore[5][10]<=Wgt_5_10;WeightsStore[5][11]<=Wgt_5_11;WeightsStore[5][12]<=Wgt_5_12;WeightsStore[5][13]<=Wgt_5_13;WeightsStore[5][14]<=Wgt_5_14;WeightsStore[5][15]<=Wgt_5_15;WeightsStore[5][16]<=Wgt_5_16;WeightsStore[5][17]<=Wgt_5_17;WeightsStore[5][18]<=Wgt_5_18;WeightsStore[5][19]<=Wgt_5_19;WeightsStore[5][20]<=Wgt_5_20;WeightsStore[5][21]<=Wgt_5_21;WeightsStore[5][22]<=Wgt_5_22;WeightsStore[5][23]<=Wgt_5_23;WeightsStore[5][24]<=Wgt_5_24;WeightsStore[5][25]<=Wgt_5_25;WeightsStore[5][26]<=Wgt_5_26;WeightsStore[5][27]<=Wgt_5_27;WeightsStore[5][28]<=Wgt_5_28;WeightsStore[5][29]<=Wgt_5_29;WeightsStore[5][30]<=Wgt_5_30;WeightsStore[5][31]<=Wgt_5_31;WeightsStore[5][32]<=Wgt_5_32;WeightsStore[5][33]<=Wgt_5_33;WeightsStore[5][34]<=Wgt_5_34;WeightsStore[5][35]<=Wgt_5_35;WeightsStore[5][36]<=Wgt_5_36;WeightsStore[5][37]<=Wgt_5_37;WeightsStore[5][38]<=Wgt_5_38;WeightsStore[5][39]<=Wgt_5_39;WeightsStore[5][40]<=Wgt_5_40;WeightsStore[5][41]<=Wgt_5_41;WeightsStore[5][42]<=Wgt_5_42;WeightsStore[5][43]<=Wgt_5_43;WeightsStore[5][44]<=Wgt_5_44;WeightsStore[5][45]<=Wgt_5_45;WeightsStore[5][46]<=Wgt_5_46;WeightsStore[5][47]<=Wgt_5_47;WeightsStore[5][48]<=Wgt_5_48;WeightsStore[5][49]<=Wgt_5_49;WeightsStore[5][50]<=Wgt_5_50;WeightsStore[5][51]<=Wgt_5_51;WeightsStore[5][52]<=Wgt_5_52;WeightsStore[5][53]<=Wgt_5_53;WeightsStore[5][54]<=Wgt_5_54;WeightsStore[5][55]<=Wgt_5_55;WeightsStore[5][56]<=Wgt_5_56;WeightsStore[5][57]<=Wgt_5_57;WeightsStore[5][58]<=Wgt_5_58;WeightsStore[5][59]<=Wgt_5_59;WeightsStore[5][60]<=Wgt_5_60;WeightsStore[5][61]<=Wgt_5_61;WeightsStore[5][62]<=Wgt_5_62;WeightsStore[5][63]<=Wgt_5_63;WeightsStore[5][64]<=Wgt_5_64;WeightsStore[5][65]<=Wgt_5_65;WeightsStore[5][66]<=Wgt_5_66;WeightsStore[5][67]<=Wgt_5_67;WeightsStore[5][68]<=Wgt_5_68;WeightsStore[5][69]<=Wgt_5_69;WeightsStore[5][70]<=Wgt_5_70;WeightsStore[5][71]<=Wgt_5_71;WeightsStore[5][72]<=Wgt_5_72;WeightsStore[5][73]<=Wgt_5_73;WeightsStore[5][74]<=Wgt_5_74;WeightsStore[5][75]<=Wgt_5_75;WeightsStore[5][76]<=Wgt_5_76;WeightsStore[5][77]<=Wgt_5_77;WeightsStore[5][78]<=Wgt_5_78;WeightsStore[5][79]<=Wgt_5_79;WeightsStore[5][80]<=Wgt_5_80;WeightsStore[5][81]<=Wgt_5_81;WeightsStore[5][82]<=Wgt_5_82;WeightsStore[5][83]<=Wgt_5_83;WeightsStore[5][84]<=Wgt_5_84;WeightsStore[5][85]<=Wgt_5_85;WeightsStore[5][86]<=Wgt_5_86;WeightsStore[5][87]<=Wgt_5_87;WeightsStore[5][88]<=Wgt_5_88;WeightsStore[5][89]<=Wgt_5_89;WeightsStore[5][90]<=Wgt_5_90;WeightsStore[5][91]<=Wgt_5_91;WeightsStore[5][92]<=Wgt_5_92;WeightsStore[5][93]<=Wgt_5_93;WeightsStore[5][94]<=Wgt_5_94;WeightsStore[5][95]<=Wgt_5_95;WeightsStore[5][96]<=Wgt_5_96;WeightsStore[5][97]<=Wgt_5_97;WeightsStore[5][98]<=Wgt_5_98;WeightsStore[5][99]<=Wgt_5_99;WeightsStore[5][100]<=Wgt_5_100;WeightsStore[5][101]<=Wgt_5_101;WeightsStore[5][102]<=Wgt_5_102;WeightsStore[5][103]<=Wgt_5_103;WeightsStore[5][104]<=Wgt_5_104;WeightsStore[5][105]<=Wgt_5_105;WeightsStore[5][106]<=Wgt_5_106;WeightsStore[5][107]<=Wgt_5_107;WeightsStore[5][108]<=Wgt_5_108;WeightsStore[5][109]<=Wgt_5_109;WeightsStore[5][110]<=Wgt_5_110;WeightsStore[5][111]<=Wgt_5_111;WeightsStore[5][112]<=Wgt_5_112;WeightsStore[5][113]<=Wgt_5_113;WeightsStore[5][114]<=Wgt_5_114;WeightsStore[5][115]<=Wgt_5_115;WeightsStore[5][116]<=Wgt_5_116;WeightsStore[5][117]<=Wgt_5_117;WeightsStore[5][118]<=Wgt_5_118;WeightsStore[5][119]<=Wgt_5_119;WeightsStore[5][120]<=Wgt_5_120;WeightsStore[5][121]<=Wgt_5_121;WeightsStore[5][122]<=Wgt_5_122;WeightsStore[5][123]<=Wgt_5_123;WeightsStore[5][124]<=Wgt_5_124;WeightsStore[5][125]<=Wgt_5_125;WeightsStore[5][126]<=Wgt_5_126;WeightsStore[5][127]<=Wgt_5_127;WeightsStore[5][128]<=Wgt_5_128;WeightsStore[5][129]<=Wgt_5_129;WeightsStore[5][130]<=Wgt_5_130;WeightsStore[5][131]<=Wgt_5_131;WeightsStore[5][132]<=Wgt_5_132;WeightsStore[5][133]<=Wgt_5_133;WeightsStore[5][134]<=Wgt_5_134;WeightsStore[5][135]<=Wgt_5_135;WeightsStore[5][136]<=Wgt_5_136;WeightsStore[5][137]<=Wgt_5_137;WeightsStore[5][138]<=Wgt_5_138;WeightsStore[5][139]<=Wgt_5_139;WeightsStore[5][140]<=Wgt_5_140;WeightsStore[5][141]<=Wgt_5_141;WeightsStore[5][142]<=Wgt_5_142;WeightsStore[5][143]<=Wgt_5_143;WeightsStore[5][144]<=Wgt_5_144;WeightsStore[5][145]<=Wgt_5_145;WeightsStore[5][146]<=Wgt_5_146;WeightsStore[5][147]<=Wgt_5_147;WeightsStore[5][148]<=Wgt_5_148;WeightsStore[5][149]<=Wgt_5_149;WeightsStore[5][150]<=Wgt_5_150;WeightsStore[5][151]<=Wgt_5_151;WeightsStore[5][152]<=Wgt_5_152;WeightsStore[5][153]<=Wgt_5_153;WeightsStore[5][154]<=Wgt_5_154;WeightsStore[5][155]<=Wgt_5_155;WeightsStore[5][156]<=Wgt_5_156;WeightsStore[5][157]<=Wgt_5_157;WeightsStore[5][158]<=Wgt_5_158;WeightsStore[5][159]<=Wgt_5_159;WeightsStore[5][160]<=Wgt_5_160;WeightsStore[5][161]<=Wgt_5_161;WeightsStore[5][162]<=Wgt_5_162;WeightsStore[5][163]<=Wgt_5_163;WeightsStore[5][164]<=Wgt_5_164;WeightsStore[5][165]<=Wgt_5_165;WeightsStore[5][166]<=Wgt_5_166;WeightsStore[5][167]<=Wgt_5_167;WeightsStore[5][168]<=Wgt_5_168;WeightsStore[5][169]<=Wgt_5_169;WeightsStore[5][170]<=Wgt_5_170;WeightsStore[5][171]<=Wgt_5_171;WeightsStore[5][172]<=Wgt_5_172;WeightsStore[5][173]<=Wgt_5_173;WeightsStore[5][174]<=Wgt_5_174;WeightsStore[5][175]<=Wgt_5_175;WeightsStore[5][176]<=Wgt_5_176;WeightsStore[5][177]<=Wgt_5_177;WeightsStore[5][178]<=Wgt_5_178;WeightsStore[5][179]<=Wgt_5_179;WeightsStore[5][180]<=Wgt_5_180;WeightsStore[5][181]<=Wgt_5_181;WeightsStore[5][182]<=Wgt_5_182;WeightsStore[5][183]<=Wgt_5_183;WeightsStore[5][184]<=Wgt_5_184;WeightsStore[5][185]<=Wgt_5_185;WeightsStore[5][186]<=Wgt_5_186;WeightsStore[5][187]<=Wgt_5_187;WeightsStore[5][188]<=Wgt_5_188;WeightsStore[5][189]<=Wgt_5_189;WeightsStore[5][190]<=Wgt_5_190;WeightsStore[5][191]<=Wgt_5_191;WeightsStore[5][192]<=Wgt_5_192;WeightsStore[5][193]<=Wgt_5_193;WeightsStore[5][194]<=Wgt_5_194;WeightsStore[5][195]<=Wgt_5_195;WeightsStore[5][196]<=Wgt_5_196;WeightsStore[5][197]<=Wgt_5_197;WeightsStore[5][198]<=Wgt_5_198;WeightsStore[5][199]<=Wgt_5_199;WeightsStore[5][200]<=Wgt_5_200;WeightsStore[5][201]<=Wgt_5_201;WeightsStore[5][202]<=Wgt_5_202;WeightsStore[5][203]<=Wgt_5_203;WeightsStore[5][204]<=Wgt_5_204;WeightsStore[5][205]<=Wgt_5_205;WeightsStore[5][206]<=Wgt_5_206;WeightsStore[5][207]<=Wgt_5_207;WeightsStore[5][208]<=Wgt_5_208;WeightsStore[5][209]<=Wgt_5_209;WeightsStore[5][210]<=Wgt_5_210;WeightsStore[5][211]<=Wgt_5_211;WeightsStore[5][212]<=Wgt_5_212;WeightsStore[5][213]<=Wgt_5_213;WeightsStore[5][214]<=Wgt_5_214;WeightsStore[5][215]<=Wgt_5_215;WeightsStore[5][216]<=Wgt_5_216;WeightsStore[5][217]<=Wgt_5_217;WeightsStore[5][218]<=Wgt_5_218;WeightsStore[5][219]<=Wgt_5_219;WeightsStore[5][220]<=Wgt_5_220;WeightsStore[5][221]<=Wgt_5_221;WeightsStore[5][222]<=Wgt_5_222;WeightsStore[5][223]<=Wgt_5_223;WeightsStore[5][224]<=Wgt_5_224;WeightsStore[5][225]<=Wgt_5_225;WeightsStore[5][226]<=Wgt_5_226;WeightsStore[5][227]<=Wgt_5_227;WeightsStore[5][228]<=Wgt_5_228;WeightsStore[5][229]<=Wgt_5_229;WeightsStore[5][230]<=Wgt_5_230;WeightsStore[5][231]<=Wgt_5_231;WeightsStore[5][232]<=Wgt_5_232;WeightsStore[5][233]<=Wgt_5_233;WeightsStore[5][234]<=Wgt_5_234;WeightsStore[5][235]<=Wgt_5_235;WeightsStore[5][236]<=Wgt_5_236;WeightsStore[5][237]<=Wgt_5_237;WeightsStore[5][238]<=Wgt_5_238;WeightsStore[5][239]<=Wgt_5_239;WeightsStore[5][240]<=Wgt_5_240;WeightsStore[5][241]<=Wgt_5_241;WeightsStore[5][242]<=Wgt_5_242;WeightsStore[5][243]<=Wgt_5_243;WeightsStore[5][244]<=Wgt_5_244;WeightsStore[5][245]<=Wgt_5_245;WeightsStore[5][246]<=Wgt_5_246;WeightsStore[5][247]<=Wgt_5_247;WeightsStore[5][248]<=Wgt_5_248;WeightsStore[5][249]<=Wgt_5_249;WeightsStore[5][250]<=Wgt_5_250;WeightsStore[5][251]<=Wgt_5_251;WeightsStore[5][252]<=Wgt_5_252;WeightsStore[5][253]<=Wgt_5_253;WeightsStore[5][254]<=Wgt_5_254;WeightsStore[5][255]<=Wgt_5_255;WeightsStore[5][256]<=Wgt_5_256;WeightsStore[5][257]<=Wgt_5_257;WeightsStore[5][258]<=Wgt_5_258;WeightsStore[5][259]<=Wgt_5_259;WeightsStore[5][260]<=Wgt_5_260;WeightsStore[5][261]<=Wgt_5_261;WeightsStore[5][262]<=Wgt_5_262;WeightsStore[5][263]<=Wgt_5_263;WeightsStore[5][264]<=Wgt_5_264;WeightsStore[5][265]<=Wgt_5_265;WeightsStore[5][266]<=Wgt_5_266;WeightsStore[5][267]<=Wgt_5_267;WeightsStore[5][268]<=Wgt_5_268;WeightsStore[5][269]<=Wgt_5_269;WeightsStore[5][270]<=Wgt_5_270;WeightsStore[5][271]<=Wgt_5_271;WeightsStore[5][272]<=Wgt_5_272;WeightsStore[5][273]<=Wgt_5_273;WeightsStore[5][274]<=Wgt_5_274;WeightsStore[5][275]<=Wgt_5_275;WeightsStore[5][276]<=Wgt_5_276;WeightsStore[5][277]<=Wgt_5_277;WeightsStore[5][278]<=Wgt_5_278;WeightsStore[5][279]<=Wgt_5_279;WeightsStore[5][280]<=Wgt_5_280;WeightsStore[5][281]<=Wgt_5_281;WeightsStore[5][282]<=Wgt_5_282;WeightsStore[5][283]<=Wgt_5_283;WeightsStore[5][284]<=Wgt_5_284;WeightsStore[5][285]<=Wgt_5_285;WeightsStore[5][286]<=Wgt_5_286;WeightsStore[5][287]<=Wgt_5_287;WeightsStore[5][288]<=Wgt_5_288;WeightsStore[5][289]<=Wgt_5_289;WeightsStore[5][290]<=Wgt_5_290;WeightsStore[5][291]<=Wgt_5_291;WeightsStore[5][292]<=Wgt_5_292;WeightsStore[5][293]<=Wgt_5_293;WeightsStore[5][294]<=Wgt_5_294;WeightsStore[5][295]<=Wgt_5_295;WeightsStore[5][296]<=Wgt_5_296;WeightsStore[5][297]<=Wgt_5_297;WeightsStore[5][298]<=Wgt_5_298;WeightsStore[5][299]<=Wgt_5_299;WeightsStore[5][300]<=Wgt_5_300;WeightsStore[5][301]<=Wgt_5_301;WeightsStore[5][302]<=Wgt_5_302;WeightsStore[5][303]<=Wgt_5_303;WeightsStore[5][304]<=Wgt_5_304;WeightsStore[5][305]<=Wgt_5_305;WeightsStore[5][306]<=Wgt_5_306;WeightsStore[5][307]<=Wgt_5_307;WeightsStore[5][308]<=Wgt_5_308;WeightsStore[5][309]<=Wgt_5_309;WeightsStore[5][310]<=Wgt_5_310;WeightsStore[5][311]<=Wgt_5_311;WeightsStore[5][312]<=Wgt_5_312;WeightsStore[5][313]<=Wgt_5_313;WeightsStore[5][314]<=Wgt_5_314;WeightsStore[5][315]<=Wgt_5_315;WeightsStore[5][316]<=Wgt_5_316;WeightsStore[5][317]<=Wgt_5_317;WeightsStore[5][318]<=Wgt_5_318;WeightsStore[5][319]<=Wgt_5_319;WeightsStore[5][320]<=Wgt_5_320;WeightsStore[5][321]<=Wgt_5_321;WeightsStore[5][322]<=Wgt_5_322;WeightsStore[5][323]<=Wgt_5_323;WeightsStore[5][324]<=Wgt_5_324;WeightsStore[5][325]<=Wgt_5_325;WeightsStore[5][326]<=Wgt_5_326;WeightsStore[5][327]<=Wgt_5_327;WeightsStore[5][328]<=Wgt_5_328;WeightsStore[5][329]<=Wgt_5_329;WeightsStore[5][330]<=Wgt_5_330;WeightsStore[5][331]<=Wgt_5_331;WeightsStore[5][332]<=Wgt_5_332;WeightsStore[5][333]<=Wgt_5_333;WeightsStore[5][334]<=Wgt_5_334;WeightsStore[5][335]<=Wgt_5_335;WeightsStore[5][336]<=Wgt_5_336;WeightsStore[5][337]<=Wgt_5_337;WeightsStore[5][338]<=Wgt_5_338;WeightsStore[5][339]<=Wgt_5_339;WeightsStore[5][340]<=Wgt_5_340;WeightsStore[5][341]<=Wgt_5_341;WeightsStore[5][342]<=Wgt_5_342;WeightsStore[5][343]<=Wgt_5_343;WeightsStore[5][344]<=Wgt_5_344;WeightsStore[5][345]<=Wgt_5_345;WeightsStore[5][346]<=Wgt_5_346;WeightsStore[5][347]<=Wgt_5_347;WeightsStore[5][348]<=Wgt_5_348;WeightsStore[5][349]<=Wgt_5_349;WeightsStore[5][350]<=Wgt_5_350;WeightsStore[5][351]<=Wgt_5_351;WeightsStore[5][352]<=Wgt_5_352;WeightsStore[5][353]<=Wgt_5_353;WeightsStore[5][354]<=Wgt_5_354;WeightsStore[5][355]<=Wgt_5_355;WeightsStore[5][356]<=Wgt_5_356;WeightsStore[5][357]<=Wgt_5_357;WeightsStore[5][358]<=Wgt_5_358;WeightsStore[5][359]<=Wgt_5_359;WeightsStore[5][360]<=Wgt_5_360;WeightsStore[5][361]<=Wgt_5_361;WeightsStore[5][362]<=Wgt_5_362;WeightsStore[5][363]<=Wgt_5_363;WeightsStore[5][364]<=Wgt_5_364;WeightsStore[5][365]<=Wgt_5_365;WeightsStore[5][366]<=Wgt_5_366;WeightsStore[5][367]<=Wgt_5_367;WeightsStore[5][368]<=Wgt_5_368;WeightsStore[5][369]<=Wgt_5_369;WeightsStore[5][370]<=Wgt_5_370;WeightsStore[5][371]<=Wgt_5_371;WeightsStore[5][372]<=Wgt_5_372;WeightsStore[5][373]<=Wgt_5_373;WeightsStore[5][374]<=Wgt_5_374;WeightsStore[5][375]<=Wgt_5_375;WeightsStore[5][376]<=Wgt_5_376;WeightsStore[5][377]<=Wgt_5_377;WeightsStore[5][378]<=Wgt_5_378;WeightsStore[5][379]<=Wgt_5_379;WeightsStore[5][380]<=Wgt_5_380;WeightsStore[5][381]<=Wgt_5_381;WeightsStore[5][382]<=Wgt_5_382;WeightsStore[5][383]<=Wgt_5_383;WeightsStore[5][384]<=Wgt_5_384;WeightsStore[5][385]<=Wgt_5_385;WeightsStore[5][386]<=Wgt_5_386;WeightsStore[5][387]<=Wgt_5_387;WeightsStore[5][388]<=Wgt_5_388;WeightsStore[5][389]<=Wgt_5_389;WeightsStore[5][390]<=Wgt_5_390;WeightsStore[5][391]<=Wgt_5_391;WeightsStore[5][392]<=Wgt_5_392;WeightsStore[5][393]<=Wgt_5_393;WeightsStore[5][394]<=Wgt_5_394;WeightsStore[5][395]<=Wgt_5_395;WeightsStore[5][396]<=Wgt_5_396;WeightsStore[5][397]<=Wgt_5_397;WeightsStore[5][398]<=Wgt_5_398;WeightsStore[5][399]<=Wgt_5_399;WeightsStore[5][400]<=Wgt_5_400;WeightsStore[5][401]<=Wgt_5_401;WeightsStore[5][402]<=Wgt_5_402;WeightsStore[5][403]<=Wgt_5_403;WeightsStore[5][404]<=Wgt_5_404;WeightsStore[5][405]<=Wgt_5_405;WeightsStore[5][406]<=Wgt_5_406;WeightsStore[5][407]<=Wgt_5_407;WeightsStore[5][408]<=Wgt_5_408;WeightsStore[5][409]<=Wgt_5_409;WeightsStore[5][410]<=Wgt_5_410;WeightsStore[5][411]<=Wgt_5_411;WeightsStore[5][412]<=Wgt_5_412;WeightsStore[5][413]<=Wgt_5_413;WeightsStore[5][414]<=Wgt_5_414;WeightsStore[5][415]<=Wgt_5_415;WeightsStore[5][416]<=Wgt_5_416;WeightsStore[5][417]<=Wgt_5_417;WeightsStore[5][418]<=Wgt_5_418;WeightsStore[5][419]<=Wgt_5_419;WeightsStore[5][420]<=Wgt_5_420;WeightsStore[5][421]<=Wgt_5_421;WeightsStore[5][422]<=Wgt_5_422;WeightsStore[5][423]<=Wgt_5_423;WeightsStore[5][424]<=Wgt_5_424;WeightsStore[5][425]<=Wgt_5_425;WeightsStore[5][426]<=Wgt_5_426;WeightsStore[5][427]<=Wgt_5_427;WeightsStore[5][428]<=Wgt_5_428;WeightsStore[5][429]<=Wgt_5_429;WeightsStore[5][430]<=Wgt_5_430;WeightsStore[5][431]<=Wgt_5_431;WeightsStore[5][432]<=Wgt_5_432;WeightsStore[5][433]<=Wgt_5_433;WeightsStore[5][434]<=Wgt_5_434;WeightsStore[5][435]<=Wgt_5_435;WeightsStore[5][436]<=Wgt_5_436;WeightsStore[5][437]<=Wgt_5_437;WeightsStore[5][438]<=Wgt_5_438;WeightsStore[5][439]<=Wgt_5_439;WeightsStore[5][440]<=Wgt_5_440;WeightsStore[5][441]<=Wgt_5_441;WeightsStore[5][442]<=Wgt_5_442;WeightsStore[5][443]<=Wgt_5_443;WeightsStore[5][444]<=Wgt_5_444;WeightsStore[5][445]<=Wgt_5_445;WeightsStore[5][446]<=Wgt_5_446;WeightsStore[5][447]<=Wgt_5_447;WeightsStore[5][448]<=Wgt_5_448;WeightsStore[5][449]<=Wgt_5_449;WeightsStore[5][450]<=Wgt_5_450;WeightsStore[5][451]<=Wgt_5_451;WeightsStore[5][452]<=Wgt_5_452;WeightsStore[5][453]<=Wgt_5_453;WeightsStore[5][454]<=Wgt_5_454;WeightsStore[5][455]<=Wgt_5_455;WeightsStore[5][456]<=Wgt_5_456;WeightsStore[5][457]<=Wgt_5_457;WeightsStore[5][458]<=Wgt_5_458;WeightsStore[5][459]<=Wgt_5_459;WeightsStore[5][460]<=Wgt_5_460;WeightsStore[5][461]<=Wgt_5_461;WeightsStore[5][462]<=Wgt_5_462;WeightsStore[5][463]<=Wgt_5_463;WeightsStore[5][464]<=Wgt_5_464;WeightsStore[5][465]<=Wgt_5_465;WeightsStore[5][466]<=Wgt_5_466;WeightsStore[5][467]<=Wgt_5_467;WeightsStore[5][468]<=Wgt_5_468;WeightsStore[5][469]<=Wgt_5_469;WeightsStore[5][470]<=Wgt_5_470;WeightsStore[5][471]<=Wgt_5_471;WeightsStore[5][472]<=Wgt_5_472;WeightsStore[5][473]<=Wgt_5_473;WeightsStore[5][474]<=Wgt_5_474;WeightsStore[5][475]<=Wgt_5_475;WeightsStore[5][476]<=Wgt_5_476;WeightsStore[5][477]<=Wgt_5_477;WeightsStore[5][478]<=Wgt_5_478;WeightsStore[5][479]<=Wgt_5_479;WeightsStore[5][480]<=Wgt_5_480;WeightsStore[5][481]<=Wgt_5_481;WeightsStore[5][482]<=Wgt_5_482;WeightsStore[5][483]<=Wgt_5_483;WeightsStore[5][484]<=Wgt_5_484;WeightsStore[5][485]<=Wgt_5_485;WeightsStore[5][486]<=Wgt_5_486;WeightsStore[5][487]<=Wgt_5_487;WeightsStore[5][488]<=Wgt_5_488;WeightsStore[5][489]<=Wgt_5_489;WeightsStore[5][490]<=Wgt_5_490;WeightsStore[5][491]<=Wgt_5_491;WeightsStore[5][492]<=Wgt_5_492;WeightsStore[5][493]<=Wgt_5_493;WeightsStore[5][494]<=Wgt_5_494;WeightsStore[5][495]<=Wgt_5_495;WeightsStore[5][496]<=Wgt_5_496;WeightsStore[5][497]<=Wgt_5_497;WeightsStore[5][498]<=Wgt_5_498;WeightsStore[5][499]<=Wgt_5_499;WeightsStore[5][500]<=Wgt_5_500;WeightsStore[5][501]<=Wgt_5_501;WeightsStore[5][502]<=Wgt_5_502;WeightsStore[5][503]<=Wgt_5_503;WeightsStore[5][504]<=Wgt_5_504;WeightsStore[5][505]<=Wgt_5_505;WeightsStore[5][506]<=Wgt_5_506;WeightsStore[5][507]<=Wgt_5_507;WeightsStore[5][508]<=Wgt_5_508;WeightsStore[5][509]<=Wgt_5_509;WeightsStore[5][510]<=Wgt_5_510;WeightsStore[5][511]<=Wgt_5_511;WeightsStore[5][512]<=Wgt_5_512;WeightsStore[5][513]<=Wgt_5_513;WeightsStore[5][514]<=Wgt_5_514;WeightsStore[5][515]<=Wgt_5_515;WeightsStore[5][516]<=Wgt_5_516;WeightsStore[5][517]<=Wgt_5_517;WeightsStore[5][518]<=Wgt_5_518;WeightsStore[5][519]<=Wgt_5_519;WeightsStore[5][520]<=Wgt_5_520;WeightsStore[5][521]<=Wgt_5_521;WeightsStore[5][522]<=Wgt_5_522;WeightsStore[5][523]<=Wgt_5_523;WeightsStore[5][524]<=Wgt_5_524;WeightsStore[5][525]<=Wgt_5_525;WeightsStore[5][526]<=Wgt_5_526;WeightsStore[5][527]<=Wgt_5_527;WeightsStore[5][528]<=Wgt_5_528;WeightsStore[5][529]<=Wgt_5_529;WeightsStore[5][530]<=Wgt_5_530;WeightsStore[5][531]<=Wgt_5_531;WeightsStore[5][532]<=Wgt_5_532;WeightsStore[5][533]<=Wgt_5_533;WeightsStore[5][534]<=Wgt_5_534;WeightsStore[5][535]<=Wgt_5_535;WeightsStore[5][536]<=Wgt_5_536;WeightsStore[5][537]<=Wgt_5_537;WeightsStore[5][538]<=Wgt_5_538;WeightsStore[5][539]<=Wgt_5_539;WeightsStore[5][540]<=Wgt_5_540;WeightsStore[5][541]<=Wgt_5_541;WeightsStore[5][542]<=Wgt_5_542;WeightsStore[5][543]<=Wgt_5_543;WeightsStore[5][544]<=Wgt_5_544;WeightsStore[5][545]<=Wgt_5_545;WeightsStore[5][546]<=Wgt_5_546;WeightsStore[5][547]<=Wgt_5_547;WeightsStore[5][548]<=Wgt_5_548;WeightsStore[5][549]<=Wgt_5_549;WeightsStore[5][550]<=Wgt_5_550;WeightsStore[5][551]<=Wgt_5_551;WeightsStore[5][552]<=Wgt_5_552;WeightsStore[5][553]<=Wgt_5_553;WeightsStore[5][554]<=Wgt_5_554;WeightsStore[5][555]<=Wgt_5_555;WeightsStore[5][556]<=Wgt_5_556;WeightsStore[5][557]<=Wgt_5_557;WeightsStore[5][558]<=Wgt_5_558;WeightsStore[5][559]<=Wgt_5_559;WeightsStore[5][560]<=Wgt_5_560;WeightsStore[5][561]<=Wgt_5_561;WeightsStore[5][562]<=Wgt_5_562;WeightsStore[5][563]<=Wgt_5_563;WeightsStore[5][564]<=Wgt_5_564;WeightsStore[5][565]<=Wgt_5_565;WeightsStore[5][566]<=Wgt_5_566;WeightsStore[5][567]<=Wgt_5_567;WeightsStore[5][568]<=Wgt_5_568;WeightsStore[5][569]<=Wgt_5_569;WeightsStore[5][570]<=Wgt_5_570;WeightsStore[5][571]<=Wgt_5_571;WeightsStore[5][572]<=Wgt_5_572;WeightsStore[5][573]<=Wgt_5_573;WeightsStore[5][574]<=Wgt_5_574;WeightsStore[5][575]<=Wgt_5_575;WeightsStore[5][576]<=Wgt_5_576;WeightsStore[5][577]<=Wgt_5_577;WeightsStore[5][578]<=Wgt_5_578;WeightsStore[5][579]<=Wgt_5_579;WeightsStore[5][580]<=Wgt_5_580;WeightsStore[5][581]<=Wgt_5_581;WeightsStore[5][582]<=Wgt_5_582;WeightsStore[5][583]<=Wgt_5_583;WeightsStore[5][584]<=Wgt_5_584;WeightsStore[5][585]<=Wgt_5_585;WeightsStore[5][586]<=Wgt_5_586;WeightsStore[5][587]<=Wgt_5_587;WeightsStore[5][588]<=Wgt_5_588;WeightsStore[5][589]<=Wgt_5_589;WeightsStore[5][590]<=Wgt_5_590;WeightsStore[5][591]<=Wgt_5_591;WeightsStore[5][592]<=Wgt_5_592;WeightsStore[5][593]<=Wgt_5_593;WeightsStore[5][594]<=Wgt_5_594;WeightsStore[5][595]<=Wgt_5_595;WeightsStore[5][596]<=Wgt_5_596;WeightsStore[5][597]<=Wgt_5_597;WeightsStore[5][598]<=Wgt_5_598;WeightsStore[5][599]<=Wgt_5_599;WeightsStore[5][600]<=Wgt_5_600;WeightsStore[5][601]<=Wgt_5_601;WeightsStore[5][602]<=Wgt_5_602;WeightsStore[5][603]<=Wgt_5_603;WeightsStore[5][604]<=Wgt_5_604;WeightsStore[5][605]<=Wgt_5_605;WeightsStore[5][606]<=Wgt_5_606;WeightsStore[5][607]<=Wgt_5_607;WeightsStore[5][608]<=Wgt_5_608;WeightsStore[5][609]<=Wgt_5_609;WeightsStore[5][610]<=Wgt_5_610;WeightsStore[5][611]<=Wgt_5_611;WeightsStore[5][612]<=Wgt_5_612;WeightsStore[5][613]<=Wgt_5_613;WeightsStore[5][614]<=Wgt_5_614;WeightsStore[5][615]<=Wgt_5_615;WeightsStore[5][616]<=Wgt_5_616;WeightsStore[5][617]<=Wgt_5_617;WeightsStore[5][618]<=Wgt_5_618;WeightsStore[5][619]<=Wgt_5_619;WeightsStore[5][620]<=Wgt_5_620;WeightsStore[5][621]<=Wgt_5_621;WeightsStore[5][622]<=Wgt_5_622;WeightsStore[5][623]<=Wgt_5_623;WeightsStore[5][624]<=Wgt_5_624;WeightsStore[5][625]<=Wgt_5_625;WeightsStore[5][626]<=Wgt_5_626;WeightsStore[5][627]<=Wgt_5_627;WeightsStore[5][628]<=Wgt_5_628;WeightsStore[5][629]<=Wgt_5_629;WeightsStore[5][630]<=Wgt_5_630;WeightsStore[5][631]<=Wgt_5_631;WeightsStore[5][632]<=Wgt_5_632;WeightsStore[5][633]<=Wgt_5_633;WeightsStore[5][634]<=Wgt_5_634;WeightsStore[5][635]<=Wgt_5_635;WeightsStore[5][636]<=Wgt_5_636;WeightsStore[5][637]<=Wgt_5_637;WeightsStore[5][638]<=Wgt_5_638;WeightsStore[5][639]<=Wgt_5_639;WeightsStore[5][640]<=Wgt_5_640;WeightsStore[5][641]<=Wgt_5_641;WeightsStore[5][642]<=Wgt_5_642;WeightsStore[5][643]<=Wgt_5_643;WeightsStore[5][644]<=Wgt_5_644;WeightsStore[5][645]<=Wgt_5_645;WeightsStore[5][646]<=Wgt_5_646;WeightsStore[5][647]<=Wgt_5_647;WeightsStore[5][648]<=Wgt_5_648;WeightsStore[5][649]<=Wgt_5_649;WeightsStore[5][650]<=Wgt_5_650;WeightsStore[5][651]<=Wgt_5_651;WeightsStore[5][652]<=Wgt_5_652;WeightsStore[5][653]<=Wgt_5_653;WeightsStore[5][654]<=Wgt_5_654;WeightsStore[5][655]<=Wgt_5_655;WeightsStore[5][656]<=Wgt_5_656;WeightsStore[5][657]<=Wgt_5_657;WeightsStore[5][658]<=Wgt_5_658;WeightsStore[5][659]<=Wgt_5_659;WeightsStore[5][660]<=Wgt_5_660;WeightsStore[5][661]<=Wgt_5_661;WeightsStore[5][662]<=Wgt_5_662;WeightsStore[5][663]<=Wgt_5_663;WeightsStore[5][664]<=Wgt_5_664;WeightsStore[5][665]<=Wgt_5_665;WeightsStore[5][666]<=Wgt_5_666;WeightsStore[5][667]<=Wgt_5_667;WeightsStore[5][668]<=Wgt_5_668;WeightsStore[5][669]<=Wgt_5_669;WeightsStore[5][670]<=Wgt_5_670;WeightsStore[5][671]<=Wgt_5_671;WeightsStore[5][672]<=Wgt_5_672;WeightsStore[5][673]<=Wgt_5_673;WeightsStore[5][674]<=Wgt_5_674;WeightsStore[5][675]<=Wgt_5_675;WeightsStore[5][676]<=Wgt_5_676;WeightsStore[5][677]<=Wgt_5_677;WeightsStore[5][678]<=Wgt_5_678;WeightsStore[5][679]<=Wgt_5_679;WeightsStore[5][680]<=Wgt_5_680;WeightsStore[5][681]<=Wgt_5_681;WeightsStore[5][682]<=Wgt_5_682;WeightsStore[5][683]<=Wgt_5_683;WeightsStore[5][684]<=Wgt_5_684;WeightsStore[5][685]<=Wgt_5_685;WeightsStore[5][686]<=Wgt_5_686;WeightsStore[5][687]<=Wgt_5_687;WeightsStore[5][688]<=Wgt_5_688;WeightsStore[5][689]<=Wgt_5_689;WeightsStore[5][690]<=Wgt_5_690;WeightsStore[5][691]<=Wgt_5_691;WeightsStore[5][692]<=Wgt_5_692;WeightsStore[5][693]<=Wgt_5_693;WeightsStore[5][694]<=Wgt_5_694;WeightsStore[5][695]<=Wgt_5_695;WeightsStore[5][696]<=Wgt_5_696;WeightsStore[5][697]<=Wgt_5_697;WeightsStore[5][698]<=Wgt_5_698;WeightsStore[5][699]<=Wgt_5_699;WeightsStore[5][700]<=Wgt_5_700;WeightsStore[5][701]<=Wgt_5_701;WeightsStore[5][702]<=Wgt_5_702;WeightsStore[5][703]<=Wgt_5_703;WeightsStore[5][704]<=Wgt_5_704;WeightsStore[5][705]<=Wgt_5_705;WeightsStore[5][706]<=Wgt_5_706;WeightsStore[5][707]<=Wgt_5_707;WeightsStore[5][708]<=Wgt_5_708;WeightsStore[5][709]<=Wgt_5_709;WeightsStore[5][710]<=Wgt_5_710;WeightsStore[5][711]<=Wgt_5_711;WeightsStore[5][712]<=Wgt_5_712;WeightsStore[5][713]<=Wgt_5_713;WeightsStore[5][714]<=Wgt_5_714;WeightsStore[5][715]<=Wgt_5_715;WeightsStore[5][716]<=Wgt_5_716;WeightsStore[5][717]<=Wgt_5_717;WeightsStore[5][718]<=Wgt_5_718;WeightsStore[5][719]<=Wgt_5_719;WeightsStore[5][720]<=Wgt_5_720;WeightsStore[5][721]<=Wgt_5_721;WeightsStore[5][722]<=Wgt_5_722;WeightsStore[5][723]<=Wgt_5_723;WeightsStore[5][724]<=Wgt_5_724;WeightsStore[5][725]<=Wgt_5_725;WeightsStore[5][726]<=Wgt_5_726;WeightsStore[5][727]<=Wgt_5_727;WeightsStore[5][728]<=Wgt_5_728;WeightsStore[5][729]<=Wgt_5_729;WeightsStore[5][730]<=Wgt_5_730;WeightsStore[5][731]<=Wgt_5_731;WeightsStore[5][732]<=Wgt_5_732;WeightsStore[5][733]<=Wgt_5_733;WeightsStore[5][734]<=Wgt_5_734;WeightsStore[5][735]<=Wgt_5_735;WeightsStore[5][736]<=Wgt_5_736;WeightsStore[5][737]<=Wgt_5_737;WeightsStore[5][738]<=Wgt_5_738;WeightsStore[5][739]<=Wgt_5_739;WeightsStore[5][740]<=Wgt_5_740;WeightsStore[5][741]<=Wgt_5_741;WeightsStore[5][742]<=Wgt_5_742;WeightsStore[5][743]<=Wgt_5_743;WeightsStore[5][744]<=Wgt_5_744;WeightsStore[5][745]<=Wgt_5_745;WeightsStore[5][746]<=Wgt_5_746;WeightsStore[5][747]<=Wgt_5_747;WeightsStore[5][748]<=Wgt_5_748;WeightsStore[5][749]<=Wgt_5_749;WeightsStore[5][750]<=Wgt_5_750;WeightsStore[5][751]<=Wgt_5_751;WeightsStore[5][752]<=Wgt_5_752;WeightsStore[5][753]<=Wgt_5_753;WeightsStore[5][754]<=Wgt_5_754;WeightsStore[5][755]<=Wgt_5_755;WeightsStore[5][756]<=Wgt_5_756;WeightsStore[5][757]<=Wgt_5_757;WeightsStore[5][758]<=Wgt_5_758;WeightsStore[5][759]<=Wgt_5_759;WeightsStore[5][760]<=Wgt_5_760;WeightsStore[5][761]<=Wgt_5_761;WeightsStore[5][762]<=Wgt_5_762;WeightsStore[5][763]<=Wgt_5_763;WeightsStore[5][764]<=Wgt_5_764;WeightsStore[5][765]<=Wgt_5_765;WeightsStore[5][766]<=Wgt_5_766;WeightsStore[5][767]<=Wgt_5_767;WeightsStore[5][768]<=Wgt_5_768;WeightsStore[5][769]<=Wgt_5_769;WeightsStore[5][770]<=Wgt_5_770;WeightsStore[5][771]<=Wgt_5_771;WeightsStore[5][772]<=Wgt_5_772;WeightsStore[5][773]<=Wgt_5_773;WeightsStore[5][774]<=Wgt_5_774;WeightsStore[5][775]<=Wgt_5_775;WeightsStore[5][776]<=Wgt_5_776;WeightsStore[5][777]<=Wgt_5_777;WeightsStore[5][778]<=Wgt_5_778;WeightsStore[5][779]<=Wgt_5_779;WeightsStore[5][780]<=Wgt_5_780;WeightsStore[5][781]<=Wgt_5_781;WeightsStore[5][782]<=Wgt_5_782;WeightsStore[5][783]<=Wgt_5_783;WeightsStore[5][784]<=Wgt_5_784;WeightsStore[6][0]<=Wgt_6_0;WeightsStore[6][1]<=Wgt_6_1;WeightsStore[6][2]<=Wgt_6_2;WeightsStore[6][3]<=Wgt_6_3;WeightsStore[6][4]<=Wgt_6_4;WeightsStore[6][5]<=Wgt_6_5;WeightsStore[6][6]<=Wgt_6_6;WeightsStore[6][7]<=Wgt_6_7;WeightsStore[6][8]<=Wgt_6_8;WeightsStore[6][9]<=Wgt_6_9;WeightsStore[6][10]<=Wgt_6_10;WeightsStore[6][11]<=Wgt_6_11;WeightsStore[6][12]<=Wgt_6_12;WeightsStore[6][13]<=Wgt_6_13;WeightsStore[6][14]<=Wgt_6_14;WeightsStore[6][15]<=Wgt_6_15;WeightsStore[6][16]<=Wgt_6_16;WeightsStore[6][17]<=Wgt_6_17;WeightsStore[6][18]<=Wgt_6_18;WeightsStore[6][19]<=Wgt_6_19;WeightsStore[6][20]<=Wgt_6_20;WeightsStore[6][21]<=Wgt_6_21;WeightsStore[6][22]<=Wgt_6_22;WeightsStore[6][23]<=Wgt_6_23;WeightsStore[6][24]<=Wgt_6_24;WeightsStore[6][25]<=Wgt_6_25;WeightsStore[6][26]<=Wgt_6_26;WeightsStore[6][27]<=Wgt_6_27;WeightsStore[6][28]<=Wgt_6_28;WeightsStore[6][29]<=Wgt_6_29;WeightsStore[6][30]<=Wgt_6_30;WeightsStore[6][31]<=Wgt_6_31;WeightsStore[6][32]<=Wgt_6_32;WeightsStore[6][33]<=Wgt_6_33;WeightsStore[6][34]<=Wgt_6_34;WeightsStore[6][35]<=Wgt_6_35;WeightsStore[6][36]<=Wgt_6_36;WeightsStore[6][37]<=Wgt_6_37;WeightsStore[6][38]<=Wgt_6_38;WeightsStore[6][39]<=Wgt_6_39;WeightsStore[6][40]<=Wgt_6_40;WeightsStore[6][41]<=Wgt_6_41;WeightsStore[6][42]<=Wgt_6_42;WeightsStore[6][43]<=Wgt_6_43;WeightsStore[6][44]<=Wgt_6_44;WeightsStore[6][45]<=Wgt_6_45;WeightsStore[6][46]<=Wgt_6_46;WeightsStore[6][47]<=Wgt_6_47;WeightsStore[6][48]<=Wgt_6_48;WeightsStore[6][49]<=Wgt_6_49;WeightsStore[6][50]<=Wgt_6_50;WeightsStore[6][51]<=Wgt_6_51;WeightsStore[6][52]<=Wgt_6_52;WeightsStore[6][53]<=Wgt_6_53;WeightsStore[6][54]<=Wgt_6_54;WeightsStore[6][55]<=Wgt_6_55;WeightsStore[6][56]<=Wgt_6_56;WeightsStore[6][57]<=Wgt_6_57;WeightsStore[6][58]<=Wgt_6_58;WeightsStore[6][59]<=Wgt_6_59;WeightsStore[6][60]<=Wgt_6_60;WeightsStore[6][61]<=Wgt_6_61;WeightsStore[6][62]<=Wgt_6_62;WeightsStore[6][63]<=Wgt_6_63;WeightsStore[6][64]<=Wgt_6_64;WeightsStore[6][65]<=Wgt_6_65;WeightsStore[6][66]<=Wgt_6_66;WeightsStore[6][67]<=Wgt_6_67;WeightsStore[6][68]<=Wgt_6_68;WeightsStore[6][69]<=Wgt_6_69;WeightsStore[6][70]<=Wgt_6_70;WeightsStore[6][71]<=Wgt_6_71;WeightsStore[6][72]<=Wgt_6_72;WeightsStore[6][73]<=Wgt_6_73;WeightsStore[6][74]<=Wgt_6_74;WeightsStore[6][75]<=Wgt_6_75;WeightsStore[6][76]<=Wgt_6_76;WeightsStore[6][77]<=Wgt_6_77;WeightsStore[6][78]<=Wgt_6_78;WeightsStore[6][79]<=Wgt_6_79;WeightsStore[6][80]<=Wgt_6_80;WeightsStore[6][81]<=Wgt_6_81;WeightsStore[6][82]<=Wgt_6_82;WeightsStore[6][83]<=Wgt_6_83;WeightsStore[6][84]<=Wgt_6_84;WeightsStore[6][85]<=Wgt_6_85;WeightsStore[6][86]<=Wgt_6_86;WeightsStore[6][87]<=Wgt_6_87;WeightsStore[6][88]<=Wgt_6_88;WeightsStore[6][89]<=Wgt_6_89;WeightsStore[6][90]<=Wgt_6_90;WeightsStore[6][91]<=Wgt_6_91;WeightsStore[6][92]<=Wgt_6_92;WeightsStore[6][93]<=Wgt_6_93;WeightsStore[6][94]<=Wgt_6_94;WeightsStore[6][95]<=Wgt_6_95;WeightsStore[6][96]<=Wgt_6_96;WeightsStore[6][97]<=Wgt_6_97;WeightsStore[6][98]<=Wgt_6_98;WeightsStore[6][99]<=Wgt_6_99;WeightsStore[6][100]<=Wgt_6_100;WeightsStore[6][101]<=Wgt_6_101;WeightsStore[6][102]<=Wgt_6_102;WeightsStore[6][103]<=Wgt_6_103;WeightsStore[6][104]<=Wgt_6_104;WeightsStore[6][105]<=Wgt_6_105;WeightsStore[6][106]<=Wgt_6_106;WeightsStore[6][107]<=Wgt_6_107;WeightsStore[6][108]<=Wgt_6_108;WeightsStore[6][109]<=Wgt_6_109;WeightsStore[6][110]<=Wgt_6_110;WeightsStore[6][111]<=Wgt_6_111;WeightsStore[6][112]<=Wgt_6_112;WeightsStore[6][113]<=Wgt_6_113;WeightsStore[6][114]<=Wgt_6_114;WeightsStore[6][115]<=Wgt_6_115;WeightsStore[6][116]<=Wgt_6_116;WeightsStore[6][117]<=Wgt_6_117;WeightsStore[6][118]<=Wgt_6_118;WeightsStore[6][119]<=Wgt_6_119;WeightsStore[6][120]<=Wgt_6_120;WeightsStore[6][121]<=Wgt_6_121;WeightsStore[6][122]<=Wgt_6_122;WeightsStore[6][123]<=Wgt_6_123;WeightsStore[6][124]<=Wgt_6_124;WeightsStore[6][125]<=Wgt_6_125;WeightsStore[6][126]<=Wgt_6_126;WeightsStore[6][127]<=Wgt_6_127;WeightsStore[6][128]<=Wgt_6_128;WeightsStore[6][129]<=Wgt_6_129;WeightsStore[6][130]<=Wgt_6_130;WeightsStore[6][131]<=Wgt_6_131;WeightsStore[6][132]<=Wgt_6_132;WeightsStore[6][133]<=Wgt_6_133;WeightsStore[6][134]<=Wgt_6_134;WeightsStore[6][135]<=Wgt_6_135;WeightsStore[6][136]<=Wgt_6_136;WeightsStore[6][137]<=Wgt_6_137;WeightsStore[6][138]<=Wgt_6_138;WeightsStore[6][139]<=Wgt_6_139;WeightsStore[6][140]<=Wgt_6_140;WeightsStore[6][141]<=Wgt_6_141;WeightsStore[6][142]<=Wgt_6_142;WeightsStore[6][143]<=Wgt_6_143;WeightsStore[6][144]<=Wgt_6_144;WeightsStore[6][145]<=Wgt_6_145;WeightsStore[6][146]<=Wgt_6_146;WeightsStore[6][147]<=Wgt_6_147;WeightsStore[6][148]<=Wgt_6_148;WeightsStore[6][149]<=Wgt_6_149;WeightsStore[6][150]<=Wgt_6_150;WeightsStore[6][151]<=Wgt_6_151;WeightsStore[6][152]<=Wgt_6_152;WeightsStore[6][153]<=Wgt_6_153;WeightsStore[6][154]<=Wgt_6_154;WeightsStore[6][155]<=Wgt_6_155;WeightsStore[6][156]<=Wgt_6_156;WeightsStore[6][157]<=Wgt_6_157;WeightsStore[6][158]<=Wgt_6_158;WeightsStore[6][159]<=Wgt_6_159;WeightsStore[6][160]<=Wgt_6_160;WeightsStore[6][161]<=Wgt_6_161;WeightsStore[6][162]<=Wgt_6_162;WeightsStore[6][163]<=Wgt_6_163;WeightsStore[6][164]<=Wgt_6_164;WeightsStore[6][165]<=Wgt_6_165;WeightsStore[6][166]<=Wgt_6_166;WeightsStore[6][167]<=Wgt_6_167;WeightsStore[6][168]<=Wgt_6_168;WeightsStore[6][169]<=Wgt_6_169;WeightsStore[6][170]<=Wgt_6_170;WeightsStore[6][171]<=Wgt_6_171;WeightsStore[6][172]<=Wgt_6_172;WeightsStore[6][173]<=Wgt_6_173;WeightsStore[6][174]<=Wgt_6_174;WeightsStore[6][175]<=Wgt_6_175;WeightsStore[6][176]<=Wgt_6_176;WeightsStore[6][177]<=Wgt_6_177;WeightsStore[6][178]<=Wgt_6_178;WeightsStore[6][179]<=Wgt_6_179;WeightsStore[6][180]<=Wgt_6_180;WeightsStore[6][181]<=Wgt_6_181;WeightsStore[6][182]<=Wgt_6_182;WeightsStore[6][183]<=Wgt_6_183;WeightsStore[6][184]<=Wgt_6_184;WeightsStore[6][185]<=Wgt_6_185;WeightsStore[6][186]<=Wgt_6_186;WeightsStore[6][187]<=Wgt_6_187;WeightsStore[6][188]<=Wgt_6_188;WeightsStore[6][189]<=Wgt_6_189;WeightsStore[6][190]<=Wgt_6_190;WeightsStore[6][191]<=Wgt_6_191;WeightsStore[6][192]<=Wgt_6_192;WeightsStore[6][193]<=Wgt_6_193;WeightsStore[6][194]<=Wgt_6_194;WeightsStore[6][195]<=Wgt_6_195;WeightsStore[6][196]<=Wgt_6_196;WeightsStore[6][197]<=Wgt_6_197;WeightsStore[6][198]<=Wgt_6_198;WeightsStore[6][199]<=Wgt_6_199;WeightsStore[6][200]<=Wgt_6_200;WeightsStore[6][201]<=Wgt_6_201;WeightsStore[6][202]<=Wgt_6_202;WeightsStore[6][203]<=Wgt_6_203;WeightsStore[6][204]<=Wgt_6_204;WeightsStore[6][205]<=Wgt_6_205;WeightsStore[6][206]<=Wgt_6_206;WeightsStore[6][207]<=Wgt_6_207;WeightsStore[6][208]<=Wgt_6_208;WeightsStore[6][209]<=Wgt_6_209;WeightsStore[6][210]<=Wgt_6_210;WeightsStore[6][211]<=Wgt_6_211;WeightsStore[6][212]<=Wgt_6_212;WeightsStore[6][213]<=Wgt_6_213;WeightsStore[6][214]<=Wgt_6_214;WeightsStore[6][215]<=Wgt_6_215;WeightsStore[6][216]<=Wgt_6_216;WeightsStore[6][217]<=Wgt_6_217;WeightsStore[6][218]<=Wgt_6_218;WeightsStore[6][219]<=Wgt_6_219;WeightsStore[6][220]<=Wgt_6_220;WeightsStore[6][221]<=Wgt_6_221;WeightsStore[6][222]<=Wgt_6_222;WeightsStore[6][223]<=Wgt_6_223;WeightsStore[6][224]<=Wgt_6_224;WeightsStore[6][225]<=Wgt_6_225;WeightsStore[6][226]<=Wgt_6_226;WeightsStore[6][227]<=Wgt_6_227;WeightsStore[6][228]<=Wgt_6_228;WeightsStore[6][229]<=Wgt_6_229;WeightsStore[6][230]<=Wgt_6_230;WeightsStore[6][231]<=Wgt_6_231;WeightsStore[6][232]<=Wgt_6_232;WeightsStore[6][233]<=Wgt_6_233;WeightsStore[6][234]<=Wgt_6_234;WeightsStore[6][235]<=Wgt_6_235;WeightsStore[6][236]<=Wgt_6_236;WeightsStore[6][237]<=Wgt_6_237;WeightsStore[6][238]<=Wgt_6_238;WeightsStore[6][239]<=Wgt_6_239;WeightsStore[6][240]<=Wgt_6_240;WeightsStore[6][241]<=Wgt_6_241;WeightsStore[6][242]<=Wgt_6_242;WeightsStore[6][243]<=Wgt_6_243;WeightsStore[6][244]<=Wgt_6_244;WeightsStore[6][245]<=Wgt_6_245;WeightsStore[6][246]<=Wgt_6_246;WeightsStore[6][247]<=Wgt_6_247;WeightsStore[6][248]<=Wgt_6_248;WeightsStore[6][249]<=Wgt_6_249;WeightsStore[6][250]<=Wgt_6_250;WeightsStore[6][251]<=Wgt_6_251;WeightsStore[6][252]<=Wgt_6_252;WeightsStore[6][253]<=Wgt_6_253;WeightsStore[6][254]<=Wgt_6_254;WeightsStore[6][255]<=Wgt_6_255;WeightsStore[6][256]<=Wgt_6_256;WeightsStore[6][257]<=Wgt_6_257;WeightsStore[6][258]<=Wgt_6_258;WeightsStore[6][259]<=Wgt_6_259;WeightsStore[6][260]<=Wgt_6_260;WeightsStore[6][261]<=Wgt_6_261;WeightsStore[6][262]<=Wgt_6_262;WeightsStore[6][263]<=Wgt_6_263;WeightsStore[6][264]<=Wgt_6_264;WeightsStore[6][265]<=Wgt_6_265;WeightsStore[6][266]<=Wgt_6_266;WeightsStore[6][267]<=Wgt_6_267;WeightsStore[6][268]<=Wgt_6_268;WeightsStore[6][269]<=Wgt_6_269;WeightsStore[6][270]<=Wgt_6_270;WeightsStore[6][271]<=Wgt_6_271;WeightsStore[6][272]<=Wgt_6_272;WeightsStore[6][273]<=Wgt_6_273;WeightsStore[6][274]<=Wgt_6_274;WeightsStore[6][275]<=Wgt_6_275;WeightsStore[6][276]<=Wgt_6_276;WeightsStore[6][277]<=Wgt_6_277;WeightsStore[6][278]<=Wgt_6_278;WeightsStore[6][279]<=Wgt_6_279;WeightsStore[6][280]<=Wgt_6_280;WeightsStore[6][281]<=Wgt_6_281;WeightsStore[6][282]<=Wgt_6_282;WeightsStore[6][283]<=Wgt_6_283;WeightsStore[6][284]<=Wgt_6_284;WeightsStore[6][285]<=Wgt_6_285;WeightsStore[6][286]<=Wgt_6_286;WeightsStore[6][287]<=Wgt_6_287;WeightsStore[6][288]<=Wgt_6_288;WeightsStore[6][289]<=Wgt_6_289;WeightsStore[6][290]<=Wgt_6_290;WeightsStore[6][291]<=Wgt_6_291;WeightsStore[6][292]<=Wgt_6_292;WeightsStore[6][293]<=Wgt_6_293;WeightsStore[6][294]<=Wgt_6_294;WeightsStore[6][295]<=Wgt_6_295;WeightsStore[6][296]<=Wgt_6_296;WeightsStore[6][297]<=Wgt_6_297;WeightsStore[6][298]<=Wgt_6_298;WeightsStore[6][299]<=Wgt_6_299;WeightsStore[6][300]<=Wgt_6_300;WeightsStore[6][301]<=Wgt_6_301;WeightsStore[6][302]<=Wgt_6_302;WeightsStore[6][303]<=Wgt_6_303;WeightsStore[6][304]<=Wgt_6_304;WeightsStore[6][305]<=Wgt_6_305;WeightsStore[6][306]<=Wgt_6_306;WeightsStore[6][307]<=Wgt_6_307;WeightsStore[6][308]<=Wgt_6_308;WeightsStore[6][309]<=Wgt_6_309;WeightsStore[6][310]<=Wgt_6_310;WeightsStore[6][311]<=Wgt_6_311;WeightsStore[6][312]<=Wgt_6_312;WeightsStore[6][313]<=Wgt_6_313;WeightsStore[6][314]<=Wgt_6_314;WeightsStore[6][315]<=Wgt_6_315;WeightsStore[6][316]<=Wgt_6_316;WeightsStore[6][317]<=Wgt_6_317;WeightsStore[6][318]<=Wgt_6_318;WeightsStore[6][319]<=Wgt_6_319;WeightsStore[6][320]<=Wgt_6_320;WeightsStore[6][321]<=Wgt_6_321;WeightsStore[6][322]<=Wgt_6_322;WeightsStore[6][323]<=Wgt_6_323;WeightsStore[6][324]<=Wgt_6_324;WeightsStore[6][325]<=Wgt_6_325;WeightsStore[6][326]<=Wgt_6_326;WeightsStore[6][327]<=Wgt_6_327;WeightsStore[6][328]<=Wgt_6_328;WeightsStore[6][329]<=Wgt_6_329;WeightsStore[6][330]<=Wgt_6_330;WeightsStore[6][331]<=Wgt_6_331;WeightsStore[6][332]<=Wgt_6_332;WeightsStore[6][333]<=Wgt_6_333;WeightsStore[6][334]<=Wgt_6_334;WeightsStore[6][335]<=Wgt_6_335;WeightsStore[6][336]<=Wgt_6_336;WeightsStore[6][337]<=Wgt_6_337;WeightsStore[6][338]<=Wgt_6_338;WeightsStore[6][339]<=Wgt_6_339;WeightsStore[6][340]<=Wgt_6_340;WeightsStore[6][341]<=Wgt_6_341;WeightsStore[6][342]<=Wgt_6_342;WeightsStore[6][343]<=Wgt_6_343;WeightsStore[6][344]<=Wgt_6_344;WeightsStore[6][345]<=Wgt_6_345;WeightsStore[6][346]<=Wgt_6_346;WeightsStore[6][347]<=Wgt_6_347;WeightsStore[6][348]<=Wgt_6_348;WeightsStore[6][349]<=Wgt_6_349;WeightsStore[6][350]<=Wgt_6_350;WeightsStore[6][351]<=Wgt_6_351;WeightsStore[6][352]<=Wgt_6_352;WeightsStore[6][353]<=Wgt_6_353;WeightsStore[6][354]<=Wgt_6_354;WeightsStore[6][355]<=Wgt_6_355;WeightsStore[6][356]<=Wgt_6_356;WeightsStore[6][357]<=Wgt_6_357;WeightsStore[6][358]<=Wgt_6_358;WeightsStore[6][359]<=Wgt_6_359;WeightsStore[6][360]<=Wgt_6_360;WeightsStore[6][361]<=Wgt_6_361;WeightsStore[6][362]<=Wgt_6_362;WeightsStore[6][363]<=Wgt_6_363;WeightsStore[6][364]<=Wgt_6_364;WeightsStore[6][365]<=Wgt_6_365;WeightsStore[6][366]<=Wgt_6_366;WeightsStore[6][367]<=Wgt_6_367;WeightsStore[6][368]<=Wgt_6_368;WeightsStore[6][369]<=Wgt_6_369;WeightsStore[6][370]<=Wgt_6_370;WeightsStore[6][371]<=Wgt_6_371;WeightsStore[6][372]<=Wgt_6_372;WeightsStore[6][373]<=Wgt_6_373;WeightsStore[6][374]<=Wgt_6_374;WeightsStore[6][375]<=Wgt_6_375;WeightsStore[6][376]<=Wgt_6_376;WeightsStore[6][377]<=Wgt_6_377;WeightsStore[6][378]<=Wgt_6_378;WeightsStore[6][379]<=Wgt_6_379;WeightsStore[6][380]<=Wgt_6_380;WeightsStore[6][381]<=Wgt_6_381;WeightsStore[6][382]<=Wgt_6_382;WeightsStore[6][383]<=Wgt_6_383;WeightsStore[6][384]<=Wgt_6_384;WeightsStore[6][385]<=Wgt_6_385;WeightsStore[6][386]<=Wgt_6_386;WeightsStore[6][387]<=Wgt_6_387;WeightsStore[6][388]<=Wgt_6_388;WeightsStore[6][389]<=Wgt_6_389;WeightsStore[6][390]<=Wgt_6_390;WeightsStore[6][391]<=Wgt_6_391;WeightsStore[6][392]<=Wgt_6_392;WeightsStore[6][393]<=Wgt_6_393;WeightsStore[6][394]<=Wgt_6_394;WeightsStore[6][395]<=Wgt_6_395;WeightsStore[6][396]<=Wgt_6_396;WeightsStore[6][397]<=Wgt_6_397;WeightsStore[6][398]<=Wgt_6_398;WeightsStore[6][399]<=Wgt_6_399;WeightsStore[6][400]<=Wgt_6_400;WeightsStore[6][401]<=Wgt_6_401;WeightsStore[6][402]<=Wgt_6_402;WeightsStore[6][403]<=Wgt_6_403;WeightsStore[6][404]<=Wgt_6_404;WeightsStore[6][405]<=Wgt_6_405;WeightsStore[6][406]<=Wgt_6_406;WeightsStore[6][407]<=Wgt_6_407;WeightsStore[6][408]<=Wgt_6_408;WeightsStore[6][409]<=Wgt_6_409;WeightsStore[6][410]<=Wgt_6_410;WeightsStore[6][411]<=Wgt_6_411;WeightsStore[6][412]<=Wgt_6_412;WeightsStore[6][413]<=Wgt_6_413;WeightsStore[6][414]<=Wgt_6_414;WeightsStore[6][415]<=Wgt_6_415;WeightsStore[6][416]<=Wgt_6_416;WeightsStore[6][417]<=Wgt_6_417;WeightsStore[6][418]<=Wgt_6_418;WeightsStore[6][419]<=Wgt_6_419;WeightsStore[6][420]<=Wgt_6_420;WeightsStore[6][421]<=Wgt_6_421;WeightsStore[6][422]<=Wgt_6_422;WeightsStore[6][423]<=Wgt_6_423;WeightsStore[6][424]<=Wgt_6_424;WeightsStore[6][425]<=Wgt_6_425;WeightsStore[6][426]<=Wgt_6_426;WeightsStore[6][427]<=Wgt_6_427;WeightsStore[6][428]<=Wgt_6_428;WeightsStore[6][429]<=Wgt_6_429;WeightsStore[6][430]<=Wgt_6_430;WeightsStore[6][431]<=Wgt_6_431;WeightsStore[6][432]<=Wgt_6_432;WeightsStore[6][433]<=Wgt_6_433;WeightsStore[6][434]<=Wgt_6_434;WeightsStore[6][435]<=Wgt_6_435;WeightsStore[6][436]<=Wgt_6_436;WeightsStore[6][437]<=Wgt_6_437;WeightsStore[6][438]<=Wgt_6_438;WeightsStore[6][439]<=Wgt_6_439;WeightsStore[6][440]<=Wgt_6_440;WeightsStore[6][441]<=Wgt_6_441;WeightsStore[6][442]<=Wgt_6_442;WeightsStore[6][443]<=Wgt_6_443;WeightsStore[6][444]<=Wgt_6_444;WeightsStore[6][445]<=Wgt_6_445;WeightsStore[6][446]<=Wgt_6_446;WeightsStore[6][447]<=Wgt_6_447;WeightsStore[6][448]<=Wgt_6_448;WeightsStore[6][449]<=Wgt_6_449;WeightsStore[6][450]<=Wgt_6_450;WeightsStore[6][451]<=Wgt_6_451;WeightsStore[6][452]<=Wgt_6_452;WeightsStore[6][453]<=Wgt_6_453;WeightsStore[6][454]<=Wgt_6_454;WeightsStore[6][455]<=Wgt_6_455;WeightsStore[6][456]<=Wgt_6_456;WeightsStore[6][457]<=Wgt_6_457;WeightsStore[6][458]<=Wgt_6_458;WeightsStore[6][459]<=Wgt_6_459;WeightsStore[6][460]<=Wgt_6_460;WeightsStore[6][461]<=Wgt_6_461;WeightsStore[6][462]<=Wgt_6_462;WeightsStore[6][463]<=Wgt_6_463;WeightsStore[6][464]<=Wgt_6_464;WeightsStore[6][465]<=Wgt_6_465;WeightsStore[6][466]<=Wgt_6_466;WeightsStore[6][467]<=Wgt_6_467;WeightsStore[6][468]<=Wgt_6_468;WeightsStore[6][469]<=Wgt_6_469;WeightsStore[6][470]<=Wgt_6_470;WeightsStore[6][471]<=Wgt_6_471;WeightsStore[6][472]<=Wgt_6_472;WeightsStore[6][473]<=Wgt_6_473;WeightsStore[6][474]<=Wgt_6_474;WeightsStore[6][475]<=Wgt_6_475;WeightsStore[6][476]<=Wgt_6_476;WeightsStore[6][477]<=Wgt_6_477;WeightsStore[6][478]<=Wgt_6_478;WeightsStore[6][479]<=Wgt_6_479;WeightsStore[6][480]<=Wgt_6_480;WeightsStore[6][481]<=Wgt_6_481;WeightsStore[6][482]<=Wgt_6_482;WeightsStore[6][483]<=Wgt_6_483;WeightsStore[6][484]<=Wgt_6_484;WeightsStore[6][485]<=Wgt_6_485;WeightsStore[6][486]<=Wgt_6_486;WeightsStore[6][487]<=Wgt_6_487;WeightsStore[6][488]<=Wgt_6_488;WeightsStore[6][489]<=Wgt_6_489;WeightsStore[6][490]<=Wgt_6_490;WeightsStore[6][491]<=Wgt_6_491;WeightsStore[6][492]<=Wgt_6_492;WeightsStore[6][493]<=Wgt_6_493;WeightsStore[6][494]<=Wgt_6_494;WeightsStore[6][495]<=Wgt_6_495;WeightsStore[6][496]<=Wgt_6_496;WeightsStore[6][497]<=Wgt_6_497;WeightsStore[6][498]<=Wgt_6_498;WeightsStore[6][499]<=Wgt_6_499;WeightsStore[6][500]<=Wgt_6_500;WeightsStore[6][501]<=Wgt_6_501;WeightsStore[6][502]<=Wgt_6_502;WeightsStore[6][503]<=Wgt_6_503;WeightsStore[6][504]<=Wgt_6_504;WeightsStore[6][505]<=Wgt_6_505;WeightsStore[6][506]<=Wgt_6_506;WeightsStore[6][507]<=Wgt_6_507;WeightsStore[6][508]<=Wgt_6_508;WeightsStore[6][509]<=Wgt_6_509;WeightsStore[6][510]<=Wgt_6_510;WeightsStore[6][511]<=Wgt_6_511;WeightsStore[6][512]<=Wgt_6_512;WeightsStore[6][513]<=Wgt_6_513;WeightsStore[6][514]<=Wgt_6_514;WeightsStore[6][515]<=Wgt_6_515;WeightsStore[6][516]<=Wgt_6_516;WeightsStore[6][517]<=Wgt_6_517;WeightsStore[6][518]<=Wgt_6_518;WeightsStore[6][519]<=Wgt_6_519;WeightsStore[6][520]<=Wgt_6_520;WeightsStore[6][521]<=Wgt_6_521;WeightsStore[6][522]<=Wgt_6_522;WeightsStore[6][523]<=Wgt_6_523;WeightsStore[6][524]<=Wgt_6_524;WeightsStore[6][525]<=Wgt_6_525;WeightsStore[6][526]<=Wgt_6_526;WeightsStore[6][527]<=Wgt_6_527;WeightsStore[6][528]<=Wgt_6_528;WeightsStore[6][529]<=Wgt_6_529;WeightsStore[6][530]<=Wgt_6_530;WeightsStore[6][531]<=Wgt_6_531;WeightsStore[6][532]<=Wgt_6_532;WeightsStore[6][533]<=Wgt_6_533;WeightsStore[6][534]<=Wgt_6_534;WeightsStore[6][535]<=Wgt_6_535;WeightsStore[6][536]<=Wgt_6_536;WeightsStore[6][537]<=Wgt_6_537;WeightsStore[6][538]<=Wgt_6_538;WeightsStore[6][539]<=Wgt_6_539;WeightsStore[6][540]<=Wgt_6_540;WeightsStore[6][541]<=Wgt_6_541;WeightsStore[6][542]<=Wgt_6_542;WeightsStore[6][543]<=Wgt_6_543;WeightsStore[6][544]<=Wgt_6_544;WeightsStore[6][545]<=Wgt_6_545;WeightsStore[6][546]<=Wgt_6_546;WeightsStore[6][547]<=Wgt_6_547;WeightsStore[6][548]<=Wgt_6_548;WeightsStore[6][549]<=Wgt_6_549;WeightsStore[6][550]<=Wgt_6_550;WeightsStore[6][551]<=Wgt_6_551;WeightsStore[6][552]<=Wgt_6_552;WeightsStore[6][553]<=Wgt_6_553;WeightsStore[6][554]<=Wgt_6_554;WeightsStore[6][555]<=Wgt_6_555;WeightsStore[6][556]<=Wgt_6_556;WeightsStore[6][557]<=Wgt_6_557;WeightsStore[6][558]<=Wgt_6_558;WeightsStore[6][559]<=Wgt_6_559;WeightsStore[6][560]<=Wgt_6_560;WeightsStore[6][561]<=Wgt_6_561;WeightsStore[6][562]<=Wgt_6_562;WeightsStore[6][563]<=Wgt_6_563;WeightsStore[6][564]<=Wgt_6_564;WeightsStore[6][565]<=Wgt_6_565;WeightsStore[6][566]<=Wgt_6_566;WeightsStore[6][567]<=Wgt_6_567;WeightsStore[6][568]<=Wgt_6_568;WeightsStore[6][569]<=Wgt_6_569;WeightsStore[6][570]<=Wgt_6_570;WeightsStore[6][571]<=Wgt_6_571;WeightsStore[6][572]<=Wgt_6_572;WeightsStore[6][573]<=Wgt_6_573;WeightsStore[6][574]<=Wgt_6_574;WeightsStore[6][575]<=Wgt_6_575;WeightsStore[6][576]<=Wgt_6_576;WeightsStore[6][577]<=Wgt_6_577;WeightsStore[6][578]<=Wgt_6_578;WeightsStore[6][579]<=Wgt_6_579;WeightsStore[6][580]<=Wgt_6_580;WeightsStore[6][581]<=Wgt_6_581;WeightsStore[6][582]<=Wgt_6_582;WeightsStore[6][583]<=Wgt_6_583;WeightsStore[6][584]<=Wgt_6_584;WeightsStore[6][585]<=Wgt_6_585;WeightsStore[6][586]<=Wgt_6_586;WeightsStore[6][587]<=Wgt_6_587;WeightsStore[6][588]<=Wgt_6_588;WeightsStore[6][589]<=Wgt_6_589;WeightsStore[6][590]<=Wgt_6_590;WeightsStore[6][591]<=Wgt_6_591;WeightsStore[6][592]<=Wgt_6_592;WeightsStore[6][593]<=Wgt_6_593;WeightsStore[6][594]<=Wgt_6_594;WeightsStore[6][595]<=Wgt_6_595;WeightsStore[6][596]<=Wgt_6_596;WeightsStore[6][597]<=Wgt_6_597;WeightsStore[6][598]<=Wgt_6_598;WeightsStore[6][599]<=Wgt_6_599;WeightsStore[6][600]<=Wgt_6_600;WeightsStore[6][601]<=Wgt_6_601;WeightsStore[6][602]<=Wgt_6_602;WeightsStore[6][603]<=Wgt_6_603;WeightsStore[6][604]<=Wgt_6_604;WeightsStore[6][605]<=Wgt_6_605;WeightsStore[6][606]<=Wgt_6_606;WeightsStore[6][607]<=Wgt_6_607;WeightsStore[6][608]<=Wgt_6_608;WeightsStore[6][609]<=Wgt_6_609;WeightsStore[6][610]<=Wgt_6_610;WeightsStore[6][611]<=Wgt_6_611;WeightsStore[6][612]<=Wgt_6_612;WeightsStore[6][613]<=Wgt_6_613;WeightsStore[6][614]<=Wgt_6_614;WeightsStore[6][615]<=Wgt_6_615;WeightsStore[6][616]<=Wgt_6_616;WeightsStore[6][617]<=Wgt_6_617;WeightsStore[6][618]<=Wgt_6_618;WeightsStore[6][619]<=Wgt_6_619;WeightsStore[6][620]<=Wgt_6_620;WeightsStore[6][621]<=Wgt_6_621;WeightsStore[6][622]<=Wgt_6_622;WeightsStore[6][623]<=Wgt_6_623;WeightsStore[6][624]<=Wgt_6_624;WeightsStore[6][625]<=Wgt_6_625;WeightsStore[6][626]<=Wgt_6_626;WeightsStore[6][627]<=Wgt_6_627;WeightsStore[6][628]<=Wgt_6_628;WeightsStore[6][629]<=Wgt_6_629;WeightsStore[6][630]<=Wgt_6_630;WeightsStore[6][631]<=Wgt_6_631;WeightsStore[6][632]<=Wgt_6_632;WeightsStore[6][633]<=Wgt_6_633;WeightsStore[6][634]<=Wgt_6_634;WeightsStore[6][635]<=Wgt_6_635;WeightsStore[6][636]<=Wgt_6_636;WeightsStore[6][637]<=Wgt_6_637;WeightsStore[6][638]<=Wgt_6_638;WeightsStore[6][639]<=Wgt_6_639;WeightsStore[6][640]<=Wgt_6_640;WeightsStore[6][641]<=Wgt_6_641;WeightsStore[6][642]<=Wgt_6_642;WeightsStore[6][643]<=Wgt_6_643;WeightsStore[6][644]<=Wgt_6_644;WeightsStore[6][645]<=Wgt_6_645;WeightsStore[6][646]<=Wgt_6_646;WeightsStore[6][647]<=Wgt_6_647;WeightsStore[6][648]<=Wgt_6_648;WeightsStore[6][649]<=Wgt_6_649;WeightsStore[6][650]<=Wgt_6_650;WeightsStore[6][651]<=Wgt_6_651;WeightsStore[6][652]<=Wgt_6_652;WeightsStore[6][653]<=Wgt_6_653;WeightsStore[6][654]<=Wgt_6_654;WeightsStore[6][655]<=Wgt_6_655;WeightsStore[6][656]<=Wgt_6_656;WeightsStore[6][657]<=Wgt_6_657;WeightsStore[6][658]<=Wgt_6_658;WeightsStore[6][659]<=Wgt_6_659;WeightsStore[6][660]<=Wgt_6_660;WeightsStore[6][661]<=Wgt_6_661;WeightsStore[6][662]<=Wgt_6_662;WeightsStore[6][663]<=Wgt_6_663;WeightsStore[6][664]<=Wgt_6_664;WeightsStore[6][665]<=Wgt_6_665;WeightsStore[6][666]<=Wgt_6_666;WeightsStore[6][667]<=Wgt_6_667;WeightsStore[6][668]<=Wgt_6_668;WeightsStore[6][669]<=Wgt_6_669;WeightsStore[6][670]<=Wgt_6_670;WeightsStore[6][671]<=Wgt_6_671;WeightsStore[6][672]<=Wgt_6_672;WeightsStore[6][673]<=Wgt_6_673;WeightsStore[6][674]<=Wgt_6_674;WeightsStore[6][675]<=Wgt_6_675;WeightsStore[6][676]<=Wgt_6_676;WeightsStore[6][677]<=Wgt_6_677;WeightsStore[6][678]<=Wgt_6_678;WeightsStore[6][679]<=Wgt_6_679;WeightsStore[6][680]<=Wgt_6_680;WeightsStore[6][681]<=Wgt_6_681;WeightsStore[6][682]<=Wgt_6_682;WeightsStore[6][683]<=Wgt_6_683;WeightsStore[6][684]<=Wgt_6_684;WeightsStore[6][685]<=Wgt_6_685;WeightsStore[6][686]<=Wgt_6_686;WeightsStore[6][687]<=Wgt_6_687;WeightsStore[6][688]<=Wgt_6_688;WeightsStore[6][689]<=Wgt_6_689;WeightsStore[6][690]<=Wgt_6_690;WeightsStore[6][691]<=Wgt_6_691;WeightsStore[6][692]<=Wgt_6_692;WeightsStore[6][693]<=Wgt_6_693;WeightsStore[6][694]<=Wgt_6_694;WeightsStore[6][695]<=Wgt_6_695;WeightsStore[6][696]<=Wgt_6_696;WeightsStore[6][697]<=Wgt_6_697;WeightsStore[6][698]<=Wgt_6_698;WeightsStore[6][699]<=Wgt_6_699;WeightsStore[6][700]<=Wgt_6_700;WeightsStore[6][701]<=Wgt_6_701;WeightsStore[6][702]<=Wgt_6_702;WeightsStore[6][703]<=Wgt_6_703;WeightsStore[6][704]<=Wgt_6_704;WeightsStore[6][705]<=Wgt_6_705;WeightsStore[6][706]<=Wgt_6_706;WeightsStore[6][707]<=Wgt_6_707;WeightsStore[6][708]<=Wgt_6_708;WeightsStore[6][709]<=Wgt_6_709;WeightsStore[6][710]<=Wgt_6_710;WeightsStore[6][711]<=Wgt_6_711;WeightsStore[6][712]<=Wgt_6_712;WeightsStore[6][713]<=Wgt_6_713;WeightsStore[6][714]<=Wgt_6_714;WeightsStore[6][715]<=Wgt_6_715;WeightsStore[6][716]<=Wgt_6_716;WeightsStore[6][717]<=Wgt_6_717;WeightsStore[6][718]<=Wgt_6_718;WeightsStore[6][719]<=Wgt_6_719;WeightsStore[6][720]<=Wgt_6_720;WeightsStore[6][721]<=Wgt_6_721;WeightsStore[6][722]<=Wgt_6_722;WeightsStore[6][723]<=Wgt_6_723;WeightsStore[6][724]<=Wgt_6_724;WeightsStore[6][725]<=Wgt_6_725;WeightsStore[6][726]<=Wgt_6_726;WeightsStore[6][727]<=Wgt_6_727;WeightsStore[6][728]<=Wgt_6_728;WeightsStore[6][729]<=Wgt_6_729;WeightsStore[6][730]<=Wgt_6_730;WeightsStore[6][731]<=Wgt_6_731;WeightsStore[6][732]<=Wgt_6_732;WeightsStore[6][733]<=Wgt_6_733;WeightsStore[6][734]<=Wgt_6_734;WeightsStore[6][735]<=Wgt_6_735;WeightsStore[6][736]<=Wgt_6_736;WeightsStore[6][737]<=Wgt_6_737;WeightsStore[6][738]<=Wgt_6_738;WeightsStore[6][739]<=Wgt_6_739;WeightsStore[6][740]<=Wgt_6_740;WeightsStore[6][741]<=Wgt_6_741;WeightsStore[6][742]<=Wgt_6_742;WeightsStore[6][743]<=Wgt_6_743;WeightsStore[6][744]<=Wgt_6_744;WeightsStore[6][745]<=Wgt_6_745;WeightsStore[6][746]<=Wgt_6_746;WeightsStore[6][747]<=Wgt_6_747;WeightsStore[6][748]<=Wgt_6_748;WeightsStore[6][749]<=Wgt_6_749;WeightsStore[6][750]<=Wgt_6_750;WeightsStore[6][751]<=Wgt_6_751;WeightsStore[6][752]<=Wgt_6_752;WeightsStore[6][753]<=Wgt_6_753;WeightsStore[6][754]<=Wgt_6_754;WeightsStore[6][755]<=Wgt_6_755;WeightsStore[6][756]<=Wgt_6_756;WeightsStore[6][757]<=Wgt_6_757;WeightsStore[6][758]<=Wgt_6_758;WeightsStore[6][759]<=Wgt_6_759;WeightsStore[6][760]<=Wgt_6_760;WeightsStore[6][761]<=Wgt_6_761;WeightsStore[6][762]<=Wgt_6_762;WeightsStore[6][763]<=Wgt_6_763;WeightsStore[6][764]<=Wgt_6_764;WeightsStore[6][765]<=Wgt_6_765;WeightsStore[6][766]<=Wgt_6_766;WeightsStore[6][767]<=Wgt_6_767;WeightsStore[6][768]<=Wgt_6_768;WeightsStore[6][769]<=Wgt_6_769;WeightsStore[6][770]<=Wgt_6_770;WeightsStore[6][771]<=Wgt_6_771;WeightsStore[6][772]<=Wgt_6_772;WeightsStore[6][773]<=Wgt_6_773;WeightsStore[6][774]<=Wgt_6_774;WeightsStore[6][775]<=Wgt_6_775;WeightsStore[6][776]<=Wgt_6_776;WeightsStore[6][777]<=Wgt_6_777;WeightsStore[6][778]<=Wgt_6_778;WeightsStore[6][779]<=Wgt_6_779;WeightsStore[6][780]<=Wgt_6_780;WeightsStore[6][781]<=Wgt_6_781;WeightsStore[6][782]<=Wgt_6_782;WeightsStore[6][783]<=Wgt_6_783;WeightsStore[6][784]<=Wgt_6_784;WeightsStore[7][0]<=Wgt_7_0;WeightsStore[7][1]<=Wgt_7_1;WeightsStore[7][2]<=Wgt_7_2;WeightsStore[7][3]<=Wgt_7_3;WeightsStore[7][4]<=Wgt_7_4;WeightsStore[7][5]<=Wgt_7_5;WeightsStore[7][6]<=Wgt_7_6;WeightsStore[7][7]<=Wgt_7_7;WeightsStore[7][8]<=Wgt_7_8;WeightsStore[7][9]<=Wgt_7_9;WeightsStore[7][10]<=Wgt_7_10;WeightsStore[7][11]<=Wgt_7_11;WeightsStore[7][12]<=Wgt_7_12;WeightsStore[7][13]<=Wgt_7_13;WeightsStore[7][14]<=Wgt_7_14;WeightsStore[7][15]<=Wgt_7_15;WeightsStore[7][16]<=Wgt_7_16;WeightsStore[7][17]<=Wgt_7_17;WeightsStore[7][18]<=Wgt_7_18;WeightsStore[7][19]<=Wgt_7_19;WeightsStore[7][20]<=Wgt_7_20;WeightsStore[7][21]<=Wgt_7_21;WeightsStore[7][22]<=Wgt_7_22;WeightsStore[7][23]<=Wgt_7_23;WeightsStore[7][24]<=Wgt_7_24;WeightsStore[7][25]<=Wgt_7_25;WeightsStore[7][26]<=Wgt_7_26;WeightsStore[7][27]<=Wgt_7_27;WeightsStore[7][28]<=Wgt_7_28;WeightsStore[7][29]<=Wgt_7_29;WeightsStore[7][30]<=Wgt_7_30;WeightsStore[7][31]<=Wgt_7_31;WeightsStore[7][32]<=Wgt_7_32;WeightsStore[7][33]<=Wgt_7_33;WeightsStore[7][34]<=Wgt_7_34;WeightsStore[7][35]<=Wgt_7_35;WeightsStore[7][36]<=Wgt_7_36;WeightsStore[7][37]<=Wgt_7_37;WeightsStore[7][38]<=Wgt_7_38;WeightsStore[7][39]<=Wgt_7_39;WeightsStore[7][40]<=Wgt_7_40;WeightsStore[7][41]<=Wgt_7_41;WeightsStore[7][42]<=Wgt_7_42;WeightsStore[7][43]<=Wgt_7_43;WeightsStore[7][44]<=Wgt_7_44;WeightsStore[7][45]<=Wgt_7_45;WeightsStore[7][46]<=Wgt_7_46;WeightsStore[7][47]<=Wgt_7_47;WeightsStore[7][48]<=Wgt_7_48;WeightsStore[7][49]<=Wgt_7_49;WeightsStore[7][50]<=Wgt_7_50;WeightsStore[7][51]<=Wgt_7_51;WeightsStore[7][52]<=Wgt_7_52;WeightsStore[7][53]<=Wgt_7_53;WeightsStore[7][54]<=Wgt_7_54;WeightsStore[7][55]<=Wgt_7_55;WeightsStore[7][56]<=Wgt_7_56;WeightsStore[7][57]<=Wgt_7_57;WeightsStore[7][58]<=Wgt_7_58;WeightsStore[7][59]<=Wgt_7_59;WeightsStore[7][60]<=Wgt_7_60;WeightsStore[7][61]<=Wgt_7_61;WeightsStore[7][62]<=Wgt_7_62;WeightsStore[7][63]<=Wgt_7_63;WeightsStore[7][64]<=Wgt_7_64;WeightsStore[7][65]<=Wgt_7_65;WeightsStore[7][66]<=Wgt_7_66;WeightsStore[7][67]<=Wgt_7_67;WeightsStore[7][68]<=Wgt_7_68;WeightsStore[7][69]<=Wgt_7_69;WeightsStore[7][70]<=Wgt_7_70;WeightsStore[7][71]<=Wgt_7_71;WeightsStore[7][72]<=Wgt_7_72;WeightsStore[7][73]<=Wgt_7_73;WeightsStore[7][74]<=Wgt_7_74;WeightsStore[7][75]<=Wgt_7_75;WeightsStore[7][76]<=Wgt_7_76;WeightsStore[7][77]<=Wgt_7_77;WeightsStore[7][78]<=Wgt_7_78;WeightsStore[7][79]<=Wgt_7_79;WeightsStore[7][80]<=Wgt_7_80;WeightsStore[7][81]<=Wgt_7_81;WeightsStore[7][82]<=Wgt_7_82;WeightsStore[7][83]<=Wgt_7_83;WeightsStore[7][84]<=Wgt_7_84;WeightsStore[7][85]<=Wgt_7_85;WeightsStore[7][86]<=Wgt_7_86;WeightsStore[7][87]<=Wgt_7_87;WeightsStore[7][88]<=Wgt_7_88;WeightsStore[7][89]<=Wgt_7_89;WeightsStore[7][90]<=Wgt_7_90;WeightsStore[7][91]<=Wgt_7_91;WeightsStore[7][92]<=Wgt_7_92;WeightsStore[7][93]<=Wgt_7_93;WeightsStore[7][94]<=Wgt_7_94;WeightsStore[7][95]<=Wgt_7_95;WeightsStore[7][96]<=Wgt_7_96;WeightsStore[7][97]<=Wgt_7_97;WeightsStore[7][98]<=Wgt_7_98;WeightsStore[7][99]<=Wgt_7_99;WeightsStore[7][100]<=Wgt_7_100;WeightsStore[7][101]<=Wgt_7_101;WeightsStore[7][102]<=Wgt_7_102;WeightsStore[7][103]<=Wgt_7_103;WeightsStore[7][104]<=Wgt_7_104;WeightsStore[7][105]<=Wgt_7_105;WeightsStore[7][106]<=Wgt_7_106;WeightsStore[7][107]<=Wgt_7_107;WeightsStore[7][108]<=Wgt_7_108;WeightsStore[7][109]<=Wgt_7_109;WeightsStore[7][110]<=Wgt_7_110;WeightsStore[7][111]<=Wgt_7_111;WeightsStore[7][112]<=Wgt_7_112;WeightsStore[7][113]<=Wgt_7_113;WeightsStore[7][114]<=Wgt_7_114;WeightsStore[7][115]<=Wgt_7_115;WeightsStore[7][116]<=Wgt_7_116;WeightsStore[7][117]<=Wgt_7_117;WeightsStore[7][118]<=Wgt_7_118;WeightsStore[7][119]<=Wgt_7_119;WeightsStore[7][120]<=Wgt_7_120;WeightsStore[7][121]<=Wgt_7_121;WeightsStore[7][122]<=Wgt_7_122;WeightsStore[7][123]<=Wgt_7_123;WeightsStore[7][124]<=Wgt_7_124;WeightsStore[7][125]<=Wgt_7_125;WeightsStore[7][126]<=Wgt_7_126;WeightsStore[7][127]<=Wgt_7_127;WeightsStore[7][128]<=Wgt_7_128;WeightsStore[7][129]<=Wgt_7_129;WeightsStore[7][130]<=Wgt_7_130;WeightsStore[7][131]<=Wgt_7_131;WeightsStore[7][132]<=Wgt_7_132;WeightsStore[7][133]<=Wgt_7_133;WeightsStore[7][134]<=Wgt_7_134;WeightsStore[7][135]<=Wgt_7_135;WeightsStore[7][136]<=Wgt_7_136;WeightsStore[7][137]<=Wgt_7_137;WeightsStore[7][138]<=Wgt_7_138;WeightsStore[7][139]<=Wgt_7_139;WeightsStore[7][140]<=Wgt_7_140;WeightsStore[7][141]<=Wgt_7_141;WeightsStore[7][142]<=Wgt_7_142;WeightsStore[7][143]<=Wgt_7_143;WeightsStore[7][144]<=Wgt_7_144;WeightsStore[7][145]<=Wgt_7_145;WeightsStore[7][146]<=Wgt_7_146;WeightsStore[7][147]<=Wgt_7_147;WeightsStore[7][148]<=Wgt_7_148;WeightsStore[7][149]<=Wgt_7_149;WeightsStore[7][150]<=Wgt_7_150;WeightsStore[7][151]<=Wgt_7_151;WeightsStore[7][152]<=Wgt_7_152;WeightsStore[7][153]<=Wgt_7_153;WeightsStore[7][154]<=Wgt_7_154;WeightsStore[7][155]<=Wgt_7_155;WeightsStore[7][156]<=Wgt_7_156;WeightsStore[7][157]<=Wgt_7_157;WeightsStore[7][158]<=Wgt_7_158;WeightsStore[7][159]<=Wgt_7_159;WeightsStore[7][160]<=Wgt_7_160;WeightsStore[7][161]<=Wgt_7_161;WeightsStore[7][162]<=Wgt_7_162;WeightsStore[7][163]<=Wgt_7_163;WeightsStore[7][164]<=Wgt_7_164;WeightsStore[7][165]<=Wgt_7_165;WeightsStore[7][166]<=Wgt_7_166;WeightsStore[7][167]<=Wgt_7_167;WeightsStore[7][168]<=Wgt_7_168;WeightsStore[7][169]<=Wgt_7_169;WeightsStore[7][170]<=Wgt_7_170;WeightsStore[7][171]<=Wgt_7_171;WeightsStore[7][172]<=Wgt_7_172;WeightsStore[7][173]<=Wgt_7_173;WeightsStore[7][174]<=Wgt_7_174;WeightsStore[7][175]<=Wgt_7_175;WeightsStore[7][176]<=Wgt_7_176;WeightsStore[7][177]<=Wgt_7_177;WeightsStore[7][178]<=Wgt_7_178;WeightsStore[7][179]<=Wgt_7_179;WeightsStore[7][180]<=Wgt_7_180;WeightsStore[7][181]<=Wgt_7_181;WeightsStore[7][182]<=Wgt_7_182;WeightsStore[7][183]<=Wgt_7_183;WeightsStore[7][184]<=Wgt_7_184;WeightsStore[7][185]<=Wgt_7_185;WeightsStore[7][186]<=Wgt_7_186;WeightsStore[7][187]<=Wgt_7_187;WeightsStore[7][188]<=Wgt_7_188;WeightsStore[7][189]<=Wgt_7_189;WeightsStore[7][190]<=Wgt_7_190;WeightsStore[7][191]<=Wgt_7_191;WeightsStore[7][192]<=Wgt_7_192;WeightsStore[7][193]<=Wgt_7_193;WeightsStore[7][194]<=Wgt_7_194;WeightsStore[7][195]<=Wgt_7_195;WeightsStore[7][196]<=Wgt_7_196;WeightsStore[7][197]<=Wgt_7_197;WeightsStore[7][198]<=Wgt_7_198;WeightsStore[7][199]<=Wgt_7_199;WeightsStore[7][200]<=Wgt_7_200;WeightsStore[7][201]<=Wgt_7_201;WeightsStore[7][202]<=Wgt_7_202;WeightsStore[7][203]<=Wgt_7_203;WeightsStore[7][204]<=Wgt_7_204;WeightsStore[7][205]<=Wgt_7_205;WeightsStore[7][206]<=Wgt_7_206;WeightsStore[7][207]<=Wgt_7_207;WeightsStore[7][208]<=Wgt_7_208;WeightsStore[7][209]<=Wgt_7_209;WeightsStore[7][210]<=Wgt_7_210;WeightsStore[7][211]<=Wgt_7_211;WeightsStore[7][212]<=Wgt_7_212;WeightsStore[7][213]<=Wgt_7_213;WeightsStore[7][214]<=Wgt_7_214;WeightsStore[7][215]<=Wgt_7_215;WeightsStore[7][216]<=Wgt_7_216;WeightsStore[7][217]<=Wgt_7_217;WeightsStore[7][218]<=Wgt_7_218;WeightsStore[7][219]<=Wgt_7_219;WeightsStore[7][220]<=Wgt_7_220;WeightsStore[7][221]<=Wgt_7_221;WeightsStore[7][222]<=Wgt_7_222;WeightsStore[7][223]<=Wgt_7_223;WeightsStore[7][224]<=Wgt_7_224;WeightsStore[7][225]<=Wgt_7_225;WeightsStore[7][226]<=Wgt_7_226;WeightsStore[7][227]<=Wgt_7_227;WeightsStore[7][228]<=Wgt_7_228;WeightsStore[7][229]<=Wgt_7_229;WeightsStore[7][230]<=Wgt_7_230;WeightsStore[7][231]<=Wgt_7_231;WeightsStore[7][232]<=Wgt_7_232;WeightsStore[7][233]<=Wgt_7_233;WeightsStore[7][234]<=Wgt_7_234;WeightsStore[7][235]<=Wgt_7_235;WeightsStore[7][236]<=Wgt_7_236;WeightsStore[7][237]<=Wgt_7_237;WeightsStore[7][238]<=Wgt_7_238;WeightsStore[7][239]<=Wgt_7_239;WeightsStore[7][240]<=Wgt_7_240;WeightsStore[7][241]<=Wgt_7_241;WeightsStore[7][242]<=Wgt_7_242;WeightsStore[7][243]<=Wgt_7_243;WeightsStore[7][244]<=Wgt_7_244;WeightsStore[7][245]<=Wgt_7_245;WeightsStore[7][246]<=Wgt_7_246;WeightsStore[7][247]<=Wgt_7_247;WeightsStore[7][248]<=Wgt_7_248;WeightsStore[7][249]<=Wgt_7_249;WeightsStore[7][250]<=Wgt_7_250;WeightsStore[7][251]<=Wgt_7_251;WeightsStore[7][252]<=Wgt_7_252;WeightsStore[7][253]<=Wgt_7_253;WeightsStore[7][254]<=Wgt_7_254;WeightsStore[7][255]<=Wgt_7_255;WeightsStore[7][256]<=Wgt_7_256;WeightsStore[7][257]<=Wgt_7_257;WeightsStore[7][258]<=Wgt_7_258;WeightsStore[7][259]<=Wgt_7_259;WeightsStore[7][260]<=Wgt_7_260;WeightsStore[7][261]<=Wgt_7_261;WeightsStore[7][262]<=Wgt_7_262;WeightsStore[7][263]<=Wgt_7_263;WeightsStore[7][264]<=Wgt_7_264;WeightsStore[7][265]<=Wgt_7_265;WeightsStore[7][266]<=Wgt_7_266;WeightsStore[7][267]<=Wgt_7_267;WeightsStore[7][268]<=Wgt_7_268;WeightsStore[7][269]<=Wgt_7_269;WeightsStore[7][270]<=Wgt_7_270;WeightsStore[7][271]<=Wgt_7_271;WeightsStore[7][272]<=Wgt_7_272;WeightsStore[7][273]<=Wgt_7_273;WeightsStore[7][274]<=Wgt_7_274;WeightsStore[7][275]<=Wgt_7_275;WeightsStore[7][276]<=Wgt_7_276;WeightsStore[7][277]<=Wgt_7_277;WeightsStore[7][278]<=Wgt_7_278;WeightsStore[7][279]<=Wgt_7_279;WeightsStore[7][280]<=Wgt_7_280;WeightsStore[7][281]<=Wgt_7_281;WeightsStore[7][282]<=Wgt_7_282;WeightsStore[7][283]<=Wgt_7_283;WeightsStore[7][284]<=Wgt_7_284;WeightsStore[7][285]<=Wgt_7_285;WeightsStore[7][286]<=Wgt_7_286;WeightsStore[7][287]<=Wgt_7_287;WeightsStore[7][288]<=Wgt_7_288;WeightsStore[7][289]<=Wgt_7_289;WeightsStore[7][290]<=Wgt_7_290;WeightsStore[7][291]<=Wgt_7_291;WeightsStore[7][292]<=Wgt_7_292;WeightsStore[7][293]<=Wgt_7_293;WeightsStore[7][294]<=Wgt_7_294;WeightsStore[7][295]<=Wgt_7_295;WeightsStore[7][296]<=Wgt_7_296;WeightsStore[7][297]<=Wgt_7_297;WeightsStore[7][298]<=Wgt_7_298;WeightsStore[7][299]<=Wgt_7_299;WeightsStore[7][300]<=Wgt_7_300;WeightsStore[7][301]<=Wgt_7_301;WeightsStore[7][302]<=Wgt_7_302;WeightsStore[7][303]<=Wgt_7_303;WeightsStore[7][304]<=Wgt_7_304;WeightsStore[7][305]<=Wgt_7_305;WeightsStore[7][306]<=Wgt_7_306;WeightsStore[7][307]<=Wgt_7_307;WeightsStore[7][308]<=Wgt_7_308;WeightsStore[7][309]<=Wgt_7_309;WeightsStore[7][310]<=Wgt_7_310;WeightsStore[7][311]<=Wgt_7_311;WeightsStore[7][312]<=Wgt_7_312;WeightsStore[7][313]<=Wgt_7_313;WeightsStore[7][314]<=Wgt_7_314;WeightsStore[7][315]<=Wgt_7_315;WeightsStore[7][316]<=Wgt_7_316;WeightsStore[7][317]<=Wgt_7_317;WeightsStore[7][318]<=Wgt_7_318;WeightsStore[7][319]<=Wgt_7_319;WeightsStore[7][320]<=Wgt_7_320;WeightsStore[7][321]<=Wgt_7_321;WeightsStore[7][322]<=Wgt_7_322;WeightsStore[7][323]<=Wgt_7_323;WeightsStore[7][324]<=Wgt_7_324;WeightsStore[7][325]<=Wgt_7_325;WeightsStore[7][326]<=Wgt_7_326;WeightsStore[7][327]<=Wgt_7_327;WeightsStore[7][328]<=Wgt_7_328;WeightsStore[7][329]<=Wgt_7_329;WeightsStore[7][330]<=Wgt_7_330;WeightsStore[7][331]<=Wgt_7_331;WeightsStore[7][332]<=Wgt_7_332;WeightsStore[7][333]<=Wgt_7_333;WeightsStore[7][334]<=Wgt_7_334;WeightsStore[7][335]<=Wgt_7_335;WeightsStore[7][336]<=Wgt_7_336;WeightsStore[7][337]<=Wgt_7_337;WeightsStore[7][338]<=Wgt_7_338;WeightsStore[7][339]<=Wgt_7_339;WeightsStore[7][340]<=Wgt_7_340;WeightsStore[7][341]<=Wgt_7_341;WeightsStore[7][342]<=Wgt_7_342;WeightsStore[7][343]<=Wgt_7_343;WeightsStore[7][344]<=Wgt_7_344;WeightsStore[7][345]<=Wgt_7_345;WeightsStore[7][346]<=Wgt_7_346;WeightsStore[7][347]<=Wgt_7_347;WeightsStore[7][348]<=Wgt_7_348;WeightsStore[7][349]<=Wgt_7_349;WeightsStore[7][350]<=Wgt_7_350;WeightsStore[7][351]<=Wgt_7_351;WeightsStore[7][352]<=Wgt_7_352;WeightsStore[7][353]<=Wgt_7_353;WeightsStore[7][354]<=Wgt_7_354;WeightsStore[7][355]<=Wgt_7_355;WeightsStore[7][356]<=Wgt_7_356;WeightsStore[7][357]<=Wgt_7_357;WeightsStore[7][358]<=Wgt_7_358;WeightsStore[7][359]<=Wgt_7_359;WeightsStore[7][360]<=Wgt_7_360;WeightsStore[7][361]<=Wgt_7_361;WeightsStore[7][362]<=Wgt_7_362;WeightsStore[7][363]<=Wgt_7_363;WeightsStore[7][364]<=Wgt_7_364;WeightsStore[7][365]<=Wgt_7_365;WeightsStore[7][366]<=Wgt_7_366;WeightsStore[7][367]<=Wgt_7_367;WeightsStore[7][368]<=Wgt_7_368;WeightsStore[7][369]<=Wgt_7_369;WeightsStore[7][370]<=Wgt_7_370;WeightsStore[7][371]<=Wgt_7_371;WeightsStore[7][372]<=Wgt_7_372;WeightsStore[7][373]<=Wgt_7_373;WeightsStore[7][374]<=Wgt_7_374;WeightsStore[7][375]<=Wgt_7_375;WeightsStore[7][376]<=Wgt_7_376;WeightsStore[7][377]<=Wgt_7_377;WeightsStore[7][378]<=Wgt_7_378;WeightsStore[7][379]<=Wgt_7_379;WeightsStore[7][380]<=Wgt_7_380;WeightsStore[7][381]<=Wgt_7_381;WeightsStore[7][382]<=Wgt_7_382;WeightsStore[7][383]<=Wgt_7_383;WeightsStore[7][384]<=Wgt_7_384;WeightsStore[7][385]<=Wgt_7_385;WeightsStore[7][386]<=Wgt_7_386;WeightsStore[7][387]<=Wgt_7_387;WeightsStore[7][388]<=Wgt_7_388;WeightsStore[7][389]<=Wgt_7_389;WeightsStore[7][390]<=Wgt_7_390;WeightsStore[7][391]<=Wgt_7_391;WeightsStore[7][392]<=Wgt_7_392;WeightsStore[7][393]<=Wgt_7_393;WeightsStore[7][394]<=Wgt_7_394;WeightsStore[7][395]<=Wgt_7_395;WeightsStore[7][396]<=Wgt_7_396;WeightsStore[7][397]<=Wgt_7_397;WeightsStore[7][398]<=Wgt_7_398;WeightsStore[7][399]<=Wgt_7_399;WeightsStore[7][400]<=Wgt_7_400;WeightsStore[7][401]<=Wgt_7_401;WeightsStore[7][402]<=Wgt_7_402;WeightsStore[7][403]<=Wgt_7_403;WeightsStore[7][404]<=Wgt_7_404;WeightsStore[7][405]<=Wgt_7_405;WeightsStore[7][406]<=Wgt_7_406;WeightsStore[7][407]<=Wgt_7_407;WeightsStore[7][408]<=Wgt_7_408;WeightsStore[7][409]<=Wgt_7_409;WeightsStore[7][410]<=Wgt_7_410;WeightsStore[7][411]<=Wgt_7_411;WeightsStore[7][412]<=Wgt_7_412;WeightsStore[7][413]<=Wgt_7_413;WeightsStore[7][414]<=Wgt_7_414;WeightsStore[7][415]<=Wgt_7_415;WeightsStore[7][416]<=Wgt_7_416;WeightsStore[7][417]<=Wgt_7_417;WeightsStore[7][418]<=Wgt_7_418;WeightsStore[7][419]<=Wgt_7_419;WeightsStore[7][420]<=Wgt_7_420;WeightsStore[7][421]<=Wgt_7_421;WeightsStore[7][422]<=Wgt_7_422;WeightsStore[7][423]<=Wgt_7_423;WeightsStore[7][424]<=Wgt_7_424;WeightsStore[7][425]<=Wgt_7_425;WeightsStore[7][426]<=Wgt_7_426;WeightsStore[7][427]<=Wgt_7_427;WeightsStore[7][428]<=Wgt_7_428;WeightsStore[7][429]<=Wgt_7_429;WeightsStore[7][430]<=Wgt_7_430;WeightsStore[7][431]<=Wgt_7_431;WeightsStore[7][432]<=Wgt_7_432;WeightsStore[7][433]<=Wgt_7_433;WeightsStore[7][434]<=Wgt_7_434;WeightsStore[7][435]<=Wgt_7_435;WeightsStore[7][436]<=Wgt_7_436;WeightsStore[7][437]<=Wgt_7_437;WeightsStore[7][438]<=Wgt_7_438;WeightsStore[7][439]<=Wgt_7_439;WeightsStore[7][440]<=Wgt_7_440;WeightsStore[7][441]<=Wgt_7_441;WeightsStore[7][442]<=Wgt_7_442;WeightsStore[7][443]<=Wgt_7_443;WeightsStore[7][444]<=Wgt_7_444;WeightsStore[7][445]<=Wgt_7_445;WeightsStore[7][446]<=Wgt_7_446;WeightsStore[7][447]<=Wgt_7_447;WeightsStore[7][448]<=Wgt_7_448;WeightsStore[7][449]<=Wgt_7_449;WeightsStore[7][450]<=Wgt_7_450;WeightsStore[7][451]<=Wgt_7_451;WeightsStore[7][452]<=Wgt_7_452;WeightsStore[7][453]<=Wgt_7_453;WeightsStore[7][454]<=Wgt_7_454;WeightsStore[7][455]<=Wgt_7_455;WeightsStore[7][456]<=Wgt_7_456;WeightsStore[7][457]<=Wgt_7_457;WeightsStore[7][458]<=Wgt_7_458;WeightsStore[7][459]<=Wgt_7_459;WeightsStore[7][460]<=Wgt_7_460;WeightsStore[7][461]<=Wgt_7_461;WeightsStore[7][462]<=Wgt_7_462;WeightsStore[7][463]<=Wgt_7_463;WeightsStore[7][464]<=Wgt_7_464;WeightsStore[7][465]<=Wgt_7_465;WeightsStore[7][466]<=Wgt_7_466;WeightsStore[7][467]<=Wgt_7_467;WeightsStore[7][468]<=Wgt_7_468;WeightsStore[7][469]<=Wgt_7_469;WeightsStore[7][470]<=Wgt_7_470;WeightsStore[7][471]<=Wgt_7_471;WeightsStore[7][472]<=Wgt_7_472;WeightsStore[7][473]<=Wgt_7_473;WeightsStore[7][474]<=Wgt_7_474;WeightsStore[7][475]<=Wgt_7_475;WeightsStore[7][476]<=Wgt_7_476;WeightsStore[7][477]<=Wgt_7_477;WeightsStore[7][478]<=Wgt_7_478;WeightsStore[7][479]<=Wgt_7_479;WeightsStore[7][480]<=Wgt_7_480;WeightsStore[7][481]<=Wgt_7_481;WeightsStore[7][482]<=Wgt_7_482;WeightsStore[7][483]<=Wgt_7_483;WeightsStore[7][484]<=Wgt_7_484;WeightsStore[7][485]<=Wgt_7_485;WeightsStore[7][486]<=Wgt_7_486;WeightsStore[7][487]<=Wgt_7_487;WeightsStore[7][488]<=Wgt_7_488;WeightsStore[7][489]<=Wgt_7_489;WeightsStore[7][490]<=Wgt_7_490;WeightsStore[7][491]<=Wgt_7_491;WeightsStore[7][492]<=Wgt_7_492;WeightsStore[7][493]<=Wgt_7_493;WeightsStore[7][494]<=Wgt_7_494;WeightsStore[7][495]<=Wgt_7_495;WeightsStore[7][496]<=Wgt_7_496;WeightsStore[7][497]<=Wgt_7_497;WeightsStore[7][498]<=Wgt_7_498;WeightsStore[7][499]<=Wgt_7_499;WeightsStore[7][500]<=Wgt_7_500;WeightsStore[7][501]<=Wgt_7_501;WeightsStore[7][502]<=Wgt_7_502;WeightsStore[7][503]<=Wgt_7_503;WeightsStore[7][504]<=Wgt_7_504;WeightsStore[7][505]<=Wgt_7_505;WeightsStore[7][506]<=Wgt_7_506;WeightsStore[7][507]<=Wgt_7_507;WeightsStore[7][508]<=Wgt_7_508;WeightsStore[7][509]<=Wgt_7_509;WeightsStore[7][510]<=Wgt_7_510;WeightsStore[7][511]<=Wgt_7_511;WeightsStore[7][512]<=Wgt_7_512;WeightsStore[7][513]<=Wgt_7_513;WeightsStore[7][514]<=Wgt_7_514;WeightsStore[7][515]<=Wgt_7_515;WeightsStore[7][516]<=Wgt_7_516;WeightsStore[7][517]<=Wgt_7_517;WeightsStore[7][518]<=Wgt_7_518;WeightsStore[7][519]<=Wgt_7_519;WeightsStore[7][520]<=Wgt_7_520;WeightsStore[7][521]<=Wgt_7_521;WeightsStore[7][522]<=Wgt_7_522;WeightsStore[7][523]<=Wgt_7_523;WeightsStore[7][524]<=Wgt_7_524;WeightsStore[7][525]<=Wgt_7_525;WeightsStore[7][526]<=Wgt_7_526;WeightsStore[7][527]<=Wgt_7_527;WeightsStore[7][528]<=Wgt_7_528;WeightsStore[7][529]<=Wgt_7_529;WeightsStore[7][530]<=Wgt_7_530;WeightsStore[7][531]<=Wgt_7_531;WeightsStore[7][532]<=Wgt_7_532;WeightsStore[7][533]<=Wgt_7_533;WeightsStore[7][534]<=Wgt_7_534;WeightsStore[7][535]<=Wgt_7_535;WeightsStore[7][536]<=Wgt_7_536;WeightsStore[7][537]<=Wgt_7_537;WeightsStore[7][538]<=Wgt_7_538;WeightsStore[7][539]<=Wgt_7_539;WeightsStore[7][540]<=Wgt_7_540;WeightsStore[7][541]<=Wgt_7_541;WeightsStore[7][542]<=Wgt_7_542;WeightsStore[7][543]<=Wgt_7_543;WeightsStore[7][544]<=Wgt_7_544;WeightsStore[7][545]<=Wgt_7_545;WeightsStore[7][546]<=Wgt_7_546;WeightsStore[7][547]<=Wgt_7_547;WeightsStore[7][548]<=Wgt_7_548;WeightsStore[7][549]<=Wgt_7_549;WeightsStore[7][550]<=Wgt_7_550;WeightsStore[7][551]<=Wgt_7_551;WeightsStore[7][552]<=Wgt_7_552;WeightsStore[7][553]<=Wgt_7_553;WeightsStore[7][554]<=Wgt_7_554;WeightsStore[7][555]<=Wgt_7_555;WeightsStore[7][556]<=Wgt_7_556;WeightsStore[7][557]<=Wgt_7_557;WeightsStore[7][558]<=Wgt_7_558;WeightsStore[7][559]<=Wgt_7_559;WeightsStore[7][560]<=Wgt_7_560;WeightsStore[7][561]<=Wgt_7_561;WeightsStore[7][562]<=Wgt_7_562;WeightsStore[7][563]<=Wgt_7_563;WeightsStore[7][564]<=Wgt_7_564;WeightsStore[7][565]<=Wgt_7_565;WeightsStore[7][566]<=Wgt_7_566;WeightsStore[7][567]<=Wgt_7_567;WeightsStore[7][568]<=Wgt_7_568;WeightsStore[7][569]<=Wgt_7_569;WeightsStore[7][570]<=Wgt_7_570;WeightsStore[7][571]<=Wgt_7_571;WeightsStore[7][572]<=Wgt_7_572;WeightsStore[7][573]<=Wgt_7_573;WeightsStore[7][574]<=Wgt_7_574;WeightsStore[7][575]<=Wgt_7_575;WeightsStore[7][576]<=Wgt_7_576;WeightsStore[7][577]<=Wgt_7_577;WeightsStore[7][578]<=Wgt_7_578;WeightsStore[7][579]<=Wgt_7_579;WeightsStore[7][580]<=Wgt_7_580;WeightsStore[7][581]<=Wgt_7_581;WeightsStore[7][582]<=Wgt_7_582;WeightsStore[7][583]<=Wgt_7_583;WeightsStore[7][584]<=Wgt_7_584;WeightsStore[7][585]<=Wgt_7_585;WeightsStore[7][586]<=Wgt_7_586;WeightsStore[7][587]<=Wgt_7_587;WeightsStore[7][588]<=Wgt_7_588;WeightsStore[7][589]<=Wgt_7_589;WeightsStore[7][590]<=Wgt_7_590;WeightsStore[7][591]<=Wgt_7_591;WeightsStore[7][592]<=Wgt_7_592;WeightsStore[7][593]<=Wgt_7_593;WeightsStore[7][594]<=Wgt_7_594;WeightsStore[7][595]<=Wgt_7_595;WeightsStore[7][596]<=Wgt_7_596;WeightsStore[7][597]<=Wgt_7_597;WeightsStore[7][598]<=Wgt_7_598;WeightsStore[7][599]<=Wgt_7_599;WeightsStore[7][600]<=Wgt_7_600;WeightsStore[7][601]<=Wgt_7_601;WeightsStore[7][602]<=Wgt_7_602;WeightsStore[7][603]<=Wgt_7_603;WeightsStore[7][604]<=Wgt_7_604;WeightsStore[7][605]<=Wgt_7_605;WeightsStore[7][606]<=Wgt_7_606;WeightsStore[7][607]<=Wgt_7_607;WeightsStore[7][608]<=Wgt_7_608;WeightsStore[7][609]<=Wgt_7_609;WeightsStore[7][610]<=Wgt_7_610;WeightsStore[7][611]<=Wgt_7_611;WeightsStore[7][612]<=Wgt_7_612;WeightsStore[7][613]<=Wgt_7_613;WeightsStore[7][614]<=Wgt_7_614;WeightsStore[7][615]<=Wgt_7_615;WeightsStore[7][616]<=Wgt_7_616;WeightsStore[7][617]<=Wgt_7_617;WeightsStore[7][618]<=Wgt_7_618;WeightsStore[7][619]<=Wgt_7_619;WeightsStore[7][620]<=Wgt_7_620;WeightsStore[7][621]<=Wgt_7_621;WeightsStore[7][622]<=Wgt_7_622;WeightsStore[7][623]<=Wgt_7_623;WeightsStore[7][624]<=Wgt_7_624;WeightsStore[7][625]<=Wgt_7_625;WeightsStore[7][626]<=Wgt_7_626;WeightsStore[7][627]<=Wgt_7_627;WeightsStore[7][628]<=Wgt_7_628;WeightsStore[7][629]<=Wgt_7_629;WeightsStore[7][630]<=Wgt_7_630;WeightsStore[7][631]<=Wgt_7_631;WeightsStore[7][632]<=Wgt_7_632;WeightsStore[7][633]<=Wgt_7_633;WeightsStore[7][634]<=Wgt_7_634;WeightsStore[7][635]<=Wgt_7_635;WeightsStore[7][636]<=Wgt_7_636;WeightsStore[7][637]<=Wgt_7_637;WeightsStore[7][638]<=Wgt_7_638;WeightsStore[7][639]<=Wgt_7_639;WeightsStore[7][640]<=Wgt_7_640;WeightsStore[7][641]<=Wgt_7_641;WeightsStore[7][642]<=Wgt_7_642;WeightsStore[7][643]<=Wgt_7_643;WeightsStore[7][644]<=Wgt_7_644;WeightsStore[7][645]<=Wgt_7_645;WeightsStore[7][646]<=Wgt_7_646;WeightsStore[7][647]<=Wgt_7_647;WeightsStore[7][648]<=Wgt_7_648;WeightsStore[7][649]<=Wgt_7_649;WeightsStore[7][650]<=Wgt_7_650;WeightsStore[7][651]<=Wgt_7_651;WeightsStore[7][652]<=Wgt_7_652;WeightsStore[7][653]<=Wgt_7_653;WeightsStore[7][654]<=Wgt_7_654;WeightsStore[7][655]<=Wgt_7_655;WeightsStore[7][656]<=Wgt_7_656;WeightsStore[7][657]<=Wgt_7_657;WeightsStore[7][658]<=Wgt_7_658;WeightsStore[7][659]<=Wgt_7_659;WeightsStore[7][660]<=Wgt_7_660;WeightsStore[7][661]<=Wgt_7_661;WeightsStore[7][662]<=Wgt_7_662;WeightsStore[7][663]<=Wgt_7_663;WeightsStore[7][664]<=Wgt_7_664;WeightsStore[7][665]<=Wgt_7_665;WeightsStore[7][666]<=Wgt_7_666;WeightsStore[7][667]<=Wgt_7_667;WeightsStore[7][668]<=Wgt_7_668;WeightsStore[7][669]<=Wgt_7_669;WeightsStore[7][670]<=Wgt_7_670;WeightsStore[7][671]<=Wgt_7_671;WeightsStore[7][672]<=Wgt_7_672;WeightsStore[7][673]<=Wgt_7_673;WeightsStore[7][674]<=Wgt_7_674;WeightsStore[7][675]<=Wgt_7_675;WeightsStore[7][676]<=Wgt_7_676;WeightsStore[7][677]<=Wgt_7_677;WeightsStore[7][678]<=Wgt_7_678;WeightsStore[7][679]<=Wgt_7_679;WeightsStore[7][680]<=Wgt_7_680;WeightsStore[7][681]<=Wgt_7_681;WeightsStore[7][682]<=Wgt_7_682;WeightsStore[7][683]<=Wgt_7_683;WeightsStore[7][684]<=Wgt_7_684;WeightsStore[7][685]<=Wgt_7_685;WeightsStore[7][686]<=Wgt_7_686;WeightsStore[7][687]<=Wgt_7_687;WeightsStore[7][688]<=Wgt_7_688;WeightsStore[7][689]<=Wgt_7_689;WeightsStore[7][690]<=Wgt_7_690;WeightsStore[7][691]<=Wgt_7_691;WeightsStore[7][692]<=Wgt_7_692;WeightsStore[7][693]<=Wgt_7_693;WeightsStore[7][694]<=Wgt_7_694;WeightsStore[7][695]<=Wgt_7_695;WeightsStore[7][696]<=Wgt_7_696;WeightsStore[7][697]<=Wgt_7_697;WeightsStore[7][698]<=Wgt_7_698;WeightsStore[7][699]<=Wgt_7_699;WeightsStore[7][700]<=Wgt_7_700;WeightsStore[7][701]<=Wgt_7_701;WeightsStore[7][702]<=Wgt_7_702;WeightsStore[7][703]<=Wgt_7_703;WeightsStore[7][704]<=Wgt_7_704;WeightsStore[7][705]<=Wgt_7_705;WeightsStore[7][706]<=Wgt_7_706;WeightsStore[7][707]<=Wgt_7_707;WeightsStore[7][708]<=Wgt_7_708;WeightsStore[7][709]<=Wgt_7_709;WeightsStore[7][710]<=Wgt_7_710;WeightsStore[7][711]<=Wgt_7_711;WeightsStore[7][712]<=Wgt_7_712;WeightsStore[7][713]<=Wgt_7_713;WeightsStore[7][714]<=Wgt_7_714;WeightsStore[7][715]<=Wgt_7_715;WeightsStore[7][716]<=Wgt_7_716;WeightsStore[7][717]<=Wgt_7_717;WeightsStore[7][718]<=Wgt_7_718;WeightsStore[7][719]<=Wgt_7_719;WeightsStore[7][720]<=Wgt_7_720;WeightsStore[7][721]<=Wgt_7_721;WeightsStore[7][722]<=Wgt_7_722;WeightsStore[7][723]<=Wgt_7_723;WeightsStore[7][724]<=Wgt_7_724;WeightsStore[7][725]<=Wgt_7_725;WeightsStore[7][726]<=Wgt_7_726;WeightsStore[7][727]<=Wgt_7_727;WeightsStore[7][728]<=Wgt_7_728;WeightsStore[7][729]<=Wgt_7_729;WeightsStore[7][730]<=Wgt_7_730;WeightsStore[7][731]<=Wgt_7_731;WeightsStore[7][732]<=Wgt_7_732;WeightsStore[7][733]<=Wgt_7_733;WeightsStore[7][734]<=Wgt_7_734;WeightsStore[7][735]<=Wgt_7_735;WeightsStore[7][736]<=Wgt_7_736;WeightsStore[7][737]<=Wgt_7_737;WeightsStore[7][738]<=Wgt_7_738;WeightsStore[7][739]<=Wgt_7_739;WeightsStore[7][740]<=Wgt_7_740;WeightsStore[7][741]<=Wgt_7_741;WeightsStore[7][742]<=Wgt_7_742;WeightsStore[7][743]<=Wgt_7_743;WeightsStore[7][744]<=Wgt_7_744;WeightsStore[7][745]<=Wgt_7_745;WeightsStore[7][746]<=Wgt_7_746;WeightsStore[7][747]<=Wgt_7_747;WeightsStore[7][748]<=Wgt_7_748;WeightsStore[7][749]<=Wgt_7_749;WeightsStore[7][750]<=Wgt_7_750;WeightsStore[7][751]<=Wgt_7_751;WeightsStore[7][752]<=Wgt_7_752;WeightsStore[7][753]<=Wgt_7_753;WeightsStore[7][754]<=Wgt_7_754;WeightsStore[7][755]<=Wgt_7_755;WeightsStore[7][756]<=Wgt_7_756;WeightsStore[7][757]<=Wgt_7_757;WeightsStore[7][758]<=Wgt_7_758;WeightsStore[7][759]<=Wgt_7_759;WeightsStore[7][760]<=Wgt_7_760;WeightsStore[7][761]<=Wgt_7_761;WeightsStore[7][762]<=Wgt_7_762;WeightsStore[7][763]<=Wgt_7_763;WeightsStore[7][764]<=Wgt_7_764;WeightsStore[7][765]<=Wgt_7_765;WeightsStore[7][766]<=Wgt_7_766;WeightsStore[7][767]<=Wgt_7_767;WeightsStore[7][768]<=Wgt_7_768;WeightsStore[7][769]<=Wgt_7_769;WeightsStore[7][770]<=Wgt_7_770;WeightsStore[7][771]<=Wgt_7_771;WeightsStore[7][772]<=Wgt_7_772;WeightsStore[7][773]<=Wgt_7_773;WeightsStore[7][774]<=Wgt_7_774;WeightsStore[7][775]<=Wgt_7_775;WeightsStore[7][776]<=Wgt_7_776;WeightsStore[7][777]<=Wgt_7_777;WeightsStore[7][778]<=Wgt_7_778;WeightsStore[7][779]<=Wgt_7_779;WeightsStore[7][780]<=Wgt_7_780;WeightsStore[7][781]<=Wgt_7_781;WeightsStore[7][782]<=Wgt_7_782;WeightsStore[7][783]<=Wgt_7_783;WeightsStore[7][784]<=Wgt_7_784;WeightsStore[8][0]<=Wgt_8_0;WeightsStore[8][1]<=Wgt_8_1;WeightsStore[8][2]<=Wgt_8_2;WeightsStore[8][3]<=Wgt_8_3;WeightsStore[8][4]<=Wgt_8_4;WeightsStore[8][5]<=Wgt_8_5;WeightsStore[8][6]<=Wgt_8_6;WeightsStore[8][7]<=Wgt_8_7;WeightsStore[8][8]<=Wgt_8_8;WeightsStore[8][9]<=Wgt_8_9;WeightsStore[8][10]<=Wgt_8_10;WeightsStore[8][11]<=Wgt_8_11;WeightsStore[8][12]<=Wgt_8_12;WeightsStore[8][13]<=Wgt_8_13;WeightsStore[8][14]<=Wgt_8_14;WeightsStore[8][15]<=Wgt_8_15;WeightsStore[8][16]<=Wgt_8_16;WeightsStore[8][17]<=Wgt_8_17;WeightsStore[8][18]<=Wgt_8_18;WeightsStore[8][19]<=Wgt_8_19;WeightsStore[8][20]<=Wgt_8_20;WeightsStore[8][21]<=Wgt_8_21;WeightsStore[8][22]<=Wgt_8_22;WeightsStore[8][23]<=Wgt_8_23;WeightsStore[8][24]<=Wgt_8_24;WeightsStore[8][25]<=Wgt_8_25;WeightsStore[8][26]<=Wgt_8_26;WeightsStore[8][27]<=Wgt_8_27;WeightsStore[8][28]<=Wgt_8_28;WeightsStore[8][29]<=Wgt_8_29;WeightsStore[8][30]<=Wgt_8_30;WeightsStore[8][31]<=Wgt_8_31;WeightsStore[8][32]<=Wgt_8_32;WeightsStore[8][33]<=Wgt_8_33;WeightsStore[8][34]<=Wgt_8_34;WeightsStore[8][35]<=Wgt_8_35;WeightsStore[8][36]<=Wgt_8_36;WeightsStore[8][37]<=Wgt_8_37;WeightsStore[8][38]<=Wgt_8_38;WeightsStore[8][39]<=Wgt_8_39;WeightsStore[8][40]<=Wgt_8_40;WeightsStore[8][41]<=Wgt_8_41;WeightsStore[8][42]<=Wgt_8_42;WeightsStore[8][43]<=Wgt_8_43;WeightsStore[8][44]<=Wgt_8_44;WeightsStore[8][45]<=Wgt_8_45;WeightsStore[8][46]<=Wgt_8_46;WeightsStore[8][47]<=Wgt_8_47;WeightsStore[8][48]<=Wgt_8_48;WeightsStore[8][49]<=Wgt_8_49;WeightsStore[8][50]<=Wgt_8_50;WeightsStore[8][51]<=Wgt_8_51;WeightsStore[8][52]<=Wgt_8_52;WeightsStore[8][53]<=Wgt_8_53;WeightsStore[8][54]<=Wgt_8_54;WeightsStore[8][55]<=Wgt_8_55;WeightsStore[8][56]<=Wgt_8_56;WeightsStore[8][57]<=Wgt_8_57;WeightsStore[8][58]<=Wgt_8_58;WeightsStore[8][59]<=Wgt_8_59;WeightsStore[8][60]<=Wgt_8_60;WeightsStore[8][61]<=Wgt_8_61;WeightsStore[8][62]<=Wgt_8_62;WeightsStore[8][63]<=Wgt_8_63;WeightsStore[8][64]<=Wgt_8_64;WeightsStore[8][65]<=Wgt_8_65;WeightsStore[8][66]<=Wgt_8_66;WeightsStore[8][67]<=Wgt_8_67;WeightsStore[8][68]<=Wgt_8_68;WeightsStore[8][69]<=Wgt_8_69;WeightsStore[8][70]<=Wgt_8_70;WeightsStore[8][71]<=Wgt_8_71;WeightsStore[8][72]<=Wgt_8_72;WeightsStore[8][73]<=Wgt_8_73;WeightsStore[8][74]<=Wgt_8_74;WeightsStore[8][75]<=Wgt_8_75;WeightsStore[8][76]<=Wgt_8_76;WeightsStore[8][77]<=Wgt_8_77;WeightsStore[8][78]<=Wgt_8_78;WeightsStore[8][79]<=Wgt_8_79;WeightsStore[8][80]<=Wgt_8_80;WeightsStore[8][81]<=Wgt_8_81;WeightsStore[8][82]<=Wgt_8_82;WeightsStore[8][83]<=Wgt_8_83;WeightsStore[8][84]<=Wgt_8_84;WeightsStore[8][85]<=Wgt_8_85;WeightsStore[8][86]<=Wgt_8_86;WeightsStore[8][87]<=Wgt_8_87;WeightsStore[8][88]<=Wgt_8_88;WeightsStore[8][89]<=Wgt_8_89;WeightsStore[8][90]<=Wgt_8_90;WeightsStore[8][91]<=Wgt_8_91;WeightsStore[8][92]<=Wgt_8_92;WeightsStore[8][93]<=Wgt_8_93;WeightsStore[8][94]<=Wgt_8_94;WeightsStore[8][95]<=Wgt_8_95;WeightsStore[8][96]<=Wgt_8_96;WeightsStore[8][97]<=Wgt_8_97;WeightsStore[8][98]<=Wgt_8_98;WeightsStore[8][99]<=Wgt_8_99;WeightsStore[8][100]<=Wgt_8_100;WeightsStore[8][101]<=Wgt_8_101;WeightsStore[8][102]<=Wgt_8_102;WeightsStore[8][103]<=Wgt_8_103;WeightsStore[8][104]<=Wgt_8_104;WeightsStore[8][105]<=Wgt_8_105;WeightsStore[8][106]<=Wgt_8_106;WeightsStore[8][107]<=Wgt_8_107;WeightsStore[8][108]<=Wgt_8_108;WeightsStore[8][109]<=Wgt_8_109;WeightsStore[8][110]<=Wgt_8_110;WeightsStore[8][111]<=Wgt_8_111;WeightsStore[8][112]<=Wgt_8_112;WeightsStore[8][113]<=Wgt_8_113;WeightsStore[8][114]<=Wgt_8_114;WeightsStore[8][115]<=Wgt_8_115;WeightsStore[8][116]<=Wgt_8_116;WeightsStore[8][117]<=Wgt_8_117;WeightsStore[8][118]<=Wgt_8_118;WeightsStore[8][119]<=Wgt_8_119;WeightsStore[8][120]<=Wgt_8_120;WeightsStore[8][121]<=Wgt_8_121;WeightsStore[8][122]<=Wgt_8_122;WeightsStore[8][123]<=Wgt_8_123;WeightsStore[8][124]<=Wgt_8_124;WeightsStore[8][125]<=Wgt_8_125;WeightsStore[8][126]<=Wgt_8_126;WeightsStore[8][127]<=Wgt_8_127;WeightsStore[8][128]<=Wgt_8_128;WeightsStore[8][129]<=Wgt_8_129;WeightsStore[8][130]<=Wgt_8_130;WeightsStore[8][131]<=Wgt_8_131;WeightsStore[8][132]<=Wgt_8_132;WeightsStore[8][133]<=Wgt_8_133;WeightsStore[8][134]<=Wgt_8_134;WeightsStore[8][135]<=Wgt_8_135;WeightsStore[8][136]<=Wgt_8_136;WeightsStore[8][137]<=Wgt_8_137;WeightsStore[8][138]<=Wgt_8_138;WeightsStore[8][139]<=Wgt_8_139;WeightsStore[8][140]<=Wgt_8_140;WeightsStore[8][141]<=Wgt_8_141;WeightsStore[8][142]<=Wgt_8_142;WeightsStore[8][143]<=Wgt_8_143;WeightsStore[8][144]<=Wgt_8_144;WeightsStore[8][145]<=Wgt_8_145;WeightsStore[8][146]<=Wgt_8_146;WeightsStore[8][147]<=Wgt_8_147;WeightsStore[8][148]<=Wgt_8_148;WeightsStore[8][149]<=Wgt_8_149;WeightsStore[8][150]<=Wgt_8_150;WeightsStore[8][151]<=Wgt_8_151;WeightsStore[8][152]<=Wgt_8_152;WeightsStore[8][153]<=Wgt_8_153;WeightsStore[8][154]<=Wgt_8_154;WeightsStore[8][155]<=Wgt_8_155;WeightsStore[8][156]<=Wgt_8_156;WeightsStore[8][157]<=Wgt_8_157;WeightsStore[8][158]<=Wgt_8_158;WeightsStore[8][159]<=Wgt_8_159;WeightsStore[8][160]<=Wgt_8_160;WeightsStore[8][161]<=Wgt_8_161;WeightsStore[8][162]<=Wgt_8_162;WeightsStore[8][163]<=Wgt_8_163;WeightsStore[8][164]<=Wgt_8_164;WeightsStore[8][165]<=Wgt_8_165;WeightsStore[8][166]<=Wgt_8_166;WeightsStore[8][167]<=Wgt_8_167;WeightsStore[8][168]<=Wgt_8_168;WeightsStore[8][169]<=Wgt_8_169;WeightsStore[8][170]<=Wgt_8_170;WeightsStore[8][171]<=Wgt_8_171;WeightsStore[8][172]<=Wgt_8_172;WeightsStore[8][173]<=Wgt_8_173;WeightsStore[8][174]<=Wgt_8_174;WeightsStore[8][175]<=Wgt_8_175;WeightsStore[8][176]<=Wgt_8_176;WeightsStore[8][177]<=Wgt_8_177;WeightsStore[8][178]<=Wgt_8_178;WeightsStore[8][179]<=Wgt_8_179;WeightsStore[8][180]<=Wgt_8_180;WeightsStore[8][181]<=Wgt_8_181;WeightsStore[8][182]<=Wgt_8_182;WeightsStore[8][183]<=Wgt_8_183;WeightsStore[8][184]<=Wgt_8_184;WeightsStore[8][185]<=Wgt_8_185;WeightsStore[8][186]<=Wgt_8_186;WeightsStore[8][187]<=Wgt_8_187;WeightsStore[8][188]<=Wgt_8_188;WeightsStore[8][189]<=Wgt_8_189;WeightsStore[8][190]<=Wgt_8_190;WeightsStore[8][191]<=Wgt_8_191;WeightsStore[8][192]<=Wgt_8_192;WeightsStore[8][193]<=Wgt_8_193;WeightsStore[8][194]<=Wgt_8_194;WeightsStore[8][195]<=Wgt_8_195;WeightsStore[8][196]<=Wgt_8_196;WeightsStore[8][197]<=Wgt_8_197;WeightsStore[8][198]<=Wgt_8_198;WeightsStore[8][199]<=Wgt_8_199;WeightsStore[8][200]<=Wgt_8_200;WeightsStore[8][201]<=Wgt_8_201;WeightsStore[8][202]<=Wgt_8_202;WeightsStore[8][203]<=Wgt_8_203;WeightsStore[8][204]<=Wgt_8_204;WeightsStore[8][205]<=Wgt_8_205;WeightsStore[8][206]<=Wgt_8_206;WeightsStore[8][207]<=Wgt_8_207;WeightsStore[8][208]<=Wgt_8_208;WeightsStore[8][209]<=Wgt_8_209;WeightsStore[8][210]<=Wgt_8_210;WeightsStore[8][211]<=Wgt_8_211;WeightsStore[8][212]<=Wgt_8_212;WeightsStore[8][213]<=Wgt_8_213;WeightsStore[8][214]<=Wgt_8_214;WeightsStore[8][215]<=Wgt_8_215;WeightsStore[8][216]<=Wgt_8_216;WeightsStore[8][217]<=Wgt_8_217;WeightsStore[8][218]<=Wgt_8_218;WeightsStore[8][219]<=Wgt_8_219;WeightsStore[8][220]<=Wgt_8_220;WeightsStore[8][221]<=Wgt_8_221;WeightsStore[8][222]<=Wgt_8_222;WeightsStore[8][223]<=Wgt_8_223;WeightsStore[8][224]<=Wgt_8_224;WeightsStore[8][225]<=Wgt_8_225;WeightsStore[8][226]<=Wgt_8_226;WeightsStore[8][227]<=Wgt_8_227;WeightsStore[8][228]<=Wgt_8_228;WeightsStore[8][229]<=Wgt_8_229;WeightsStore[8][230]<=Wgt_8_230;WeightsStore[8][231]<=Wgt_8_231;WeightsStore[8][232]<=Wgt_8_232;WeightsStore[8][233]<=Wgt_8_233;WeightsStore[8][234]<=Wgt_8_234;WeightsStore[8][235]<=Wgt_8_235;WeightsStore[8][236]<=Wgt_8_236;WeightsStore[8][237]<=Wgt_8_237;WeightsStore[8][238]<=Wgt_8_238;WeightsStore[8][239]<=Wgt_8_239;WeightsStore[8][240]<=Wgt_8_240;WeightsStore[8][241]<=Wgt_8_241;WeightsStore[8][242]<=Wgt_8_242;WeightsStore[8][243]<=Wgt_8_243;WeightsStore[8][244]<=Wgt_8_244;WeightsStore[8][245]<=Wgt_8_245;WeightsStore[8][246]<=Wgt_8_246;WeightsStore[8][247]<=Wgt_8_247;WeightsStore[8][248]<=Wgt_8_248;WeightsStore[8][249]<=Wgt_8_249;WeightsStore[8][250]<=Wgt_8_250;WeightsStore[8][251]<=Wgt_8_251;WeightsStore[8][252]<=Wgt_8_252;WeightsStore[8][253]<=Wgt_8_253;WeightsStore[8][254]<=Wgt_8_254;WeightsStore[8][255]<=Wgt_8_255;WeightsStore[8][256]<=Wgt_8_256;WeightsStore[8][257]<=Wgt_8_257;WeightsStore[8][258]<=Wgt_8_258;WeightsStore[8][259]<=Wgt_8_259;WeightsStore[8][260]<=Wgt_8_260;WeightsStore[8][261]<=Wgt_8_261;WeightsStore[8][262]<=Wgt_8_262;WeightsStore[8][263]<=Wgt_8_263;WeightsStore[8][264]<=Wgt_8_264;WeightsStore[8][265]<=Wgt_8_265;WeightsStore[8][266]<=Wgt_8_266;WeightsStore[8][267]<=Wgt_8_267;WeightsStore[8][268]<=Wgt_8_268;WeightsStore[8][269]<=Wgt_8_269;WeightsStore[8][270]<=Wgt_8_270;WeightsStore[8][271]<=Wgt_8_271;WeightsStore[8][272]<=Wgt_8_272;WeightsStore[8][273]<=Wgt_8_273;WeightsStore[8][274]<=Wgt_8_274;WeightsStore[8][275]<=Wgt_8_275;WeightsStore[8][276]<=Wgt_8_276;WeightsStore[8][277]<=Wgt_8_277;WeightsStore[8][278]<=Wgt_8_278;WeightsStore[8][279]<=Wgt_8_279;WeightsStore[8][280]<=Wgt_8_280;WeightsStore[8][281]<=Wgt_8_281;WeightsStore[8][282]<=Wgt_8_282;WeightsStore[8][283]<=Wgt_8_283;WeightsStore[8][284]<=Wgt_8_284;WeightsStore[8][285]<=Wgt_8_285;WeightsStore[8][286]<=Wgt_8_286;WeightsStore[8][287]<=Wgt_8_287;WeightsStore[8][288]<=Wgt_8_288;WeightsStore[8][289]<=Wgt_8_289;WeightsStore[8][290]<=Wgt_8_290;WeightsStore[8][291]<=Wgt_8_291;WeightsStore[8][292]<=Wgt_8_292;WeightsStore[8][293]<=Wgt_8_293;WeightsStore[8][294]<=Wgt_8_294;WeightsStore[8][295]<=Wgt_8_295;WeightsStore[8][296]<=Wgt_8_296;WeightsStore[8][297]<=Wgt_8_297;WeightsStore[8][298]<=Wgt_8_298;WeightsStore[8][299]<=Wgt_8_299;WeightsStore[8][300]<=Wgt_8_300;WeightsStore[8][301]<=Wgt_8_301;WeightsStore[8][302]<=Wgt_8_302;WeightsStore[8][303]<=Wgt_8_303;WeightsStore[8][304]<=Wgt_8_304;WeightsStore[8][305]<=Wgt_8_305;WeightsStore[8][306]<=Wgt_8_306;WeightsStore[8][307]<=Wgt_8_307;WeightsStore[8][308]<=Wgt_8_308;WeightsStore[8][309]<=Wgt_8_309;WeightsStore[8][310]<=Wgt_8_310;WeightsStore[8][311]<=Wgt_8_311;WeightsStore[8][312]<=Wgt_8_312;WeightsStore[8][313]<=Wgt_8_313;WeightsStore[8][314]<=Wgt_8_314;WeightsStore[8][315]<=Wgt_8_315;WeightsStore[8][316]<=Wgt_8_316;WeightsStore[8][317]<=Wgt_8_317;WeightsStore[8][318]<=Wgt_8_318;WeightsStore[8][319]<=Wgt_8_319;WeightsStore[8][320]<=Wgt_8_320;WeightsStore[8][321]<=Wgt_8_321;WeightsStore[8][322]<=Wgt_8_322;WeightsStore[8][323]<=Wgt_8_323;WeightsStore[8][324]<=Wgt_8_324;WeightsStore[8][325]<=Wgt_8_325;WeightsStore[8][326]<=Wgt_8_326;WeightsStore[8][327]<=Wgt_8_327;WeightsStore[8][328]<=Wgt_8_328;WeightsStore[8][329]<=Wgt_8_329;WeightsStore[8][330]<=Wgt_8_330;WeightsStore[8][331]<=Wgt_8_331;WeightsStore[8][332]<=Wgt_8_332;WeightsStore[8][333]<=Wgt_8_333;WeightsStore[8][334]<=Wgt_8_334;WeightsStore[8][335]<=Wgt_8_335;WeightsStore[8][336]<=Wgt_8_336;WeightsStore[8][337]<=Wgt_8_337;WeightsStore[8][338]<=Wgt_8_338;WeightsStore[8][339]<=Wgt_8_339;WeightsStore[8][340]<=Wgt_8_340;WeightsStore[8][341]<=Wgt_8_341;WeightsStore[8][342]<=Wgt_8_342;WeightsStore[8][343]<=Wgt_8_343;WeightsStore[8][344]<=Wgt_8_344;WeightsStore[8][345]<=Wgt_8_345;WeightsStore[8][346]<=Wgt_8_346;WeightsStore[8][347]<=Wgt_8_347;WeightsStore[8][348]<=Wgt_8_348;WeightsStore[8][349]<=Wgt_8_349;WeightsStore[8][350]<=Wgt_8_350;WeightsStore[8][351]<=Wgt_8_351;WeightsStore[8][352]<=Wgt_8_352;WeightsStore[8][353]<=Wgt_8_353;WeightsStore[8][354]<=Wgt_8_354;WeightsStore[8][355]<=Wgt_8_355;WeightsStore[8][356]<=Wgt_8_356;WeightsStore[8][357]<=Wgt_8_357;WeightsStore[8][358]<=Wgt_8_358;WeightsStore[8][359]<=Wgt_8_359;WeightsStore[8][360]<=Wgt_8_360;WeightsStore[8][361]<=Wgt_8_361;WeightsStore[8][362]<=Wgt_8_362;WeightsStore[8][363]<=Wgt_8_363;WeightsStore[8][364]<=Wgt_8_364;WeightsStore[8][365]<=Wgt_8_365;WeightsStore[8][366]<=Wgt_8_366;WeightsStore[8][367]<=Wgt_8_367;WeightsStore[8][368]<=Wgt_8_368;WeightsStore[8][369]<=Wgt_8_369;WeightsStore[8][370]<=Wgt_8_370;WeightsStore[8][371]<=Wgt_8_371;WeightsStore[8][372]<=Wgt_8_372;WeightsStore[8][373]<=Wgt_8_373;WeightsStore[8][374]<=Wgt_8_374;WeightsStore[8][375]<=Wgt_8_375;WeightsStore[8][376]<=Wgt_8_376;WeightsStore[8][377]<=Wgt_8_377;WeightsStore[8][378]<=Wgt_8_378;WeightsStore[8][379]<=Wgt_8_379;WeightsStore[8][380]<=Wgt_8_380;WeightsStore[8][381]<=Wgt_8_381;WeightsStore[8][382]<=Wgt_8_382;WeightsStore[8][383]<=Wgt_8_383;WeightsStore[8][384]<=Wgt_8_384;WeightsStore[8][385]<=Wgt_8_385;WeightsStore[8][386]<=Wgt_8_386;WeightsStore[8][387]<=Wgt_8_387;WeightsStore[8][388]<=Wgt_8_388;WeightsStore[8][389]<=Wgt_8_389;WeightsStore[8][390]<=Wgt_8_390;WeightsStore[8][391]<=Wgt_8_391;WeightsStore[8][392]<=Wgt_8_392;WeightsStore[8][393]<=Wgt_8_393;WeightsStore[8][394]<=Wgt_8_394;WeightsStore[8][395]<=Wgt_8_395;WeightsStore[8][396]<=Wgt_8_396;WeightsStore[8][397]<=Wgt_8_397;WeightsStore[8][398]<=Wgt_8_398;WeightsStore[8][399]<=Wgt_8_399;WeightsStore[8][400]<=Wgt_8_400;WeightsStore[8][401]<=Wgt_8_401;WeightsStore[8][402]<=Wgt_8_402;WeightsStore[8][403]<=Wgt_8_403;WeightsStore[8][404]<=Wgt_8_404;WeightsStore[8][405]<=Wgt_8_405;WeightsStore[8][406]<=Wgt_8_406;WeightsStore[8][407]<=Wgt_8_407;WeightsStore[8][408]<=Wgt_8_408;WeightsStore[8][409]<=Wgt_8_409;WeightsStore[8][410]<=Wgt_8_410;WeightsStore[8][411]<=Wgt_8_411;WeightsStore[8][412]<=Wgt_8_412;WeightsStore[8][413]<=Wgt_8_413;WeightsStore[8][414]<=Wgt_8_414;WeightsStore[8][415]<=Wgt_8_415;WeightsStore[8][416]<=Wgt_8_416;WeightsStore[8][417]<=Wgt_8_417;WeightsStore[8][418]<=Wgt_8_418;WeightsStore[8][419]<=Wgt_8_419;WeightsStore[8][420]<=Wgt_8_420;WeightsStore[8][421]<=Wgt_8_421;WeightsStore[8][422]<=Wgt_8_422;WeightsStore[8][423]<=Wgt_8_423;WeightsStore[8][424]<=Wgt_8_424;WeightsStore[8][425]<=Wgt_8_425;WeightsStore[8][426]<=Wgt_8_426;WeightsStore[8][427]<=Wgt_8_427;WeightsStore[8][428]<=Wgt_8_428;WeightsStore[8][429]<=Wgt_8_429;WeightsStore[8][430]<=Wgt_8_430;WeightsStore[8][431]<=Wgt_8_431;WeightsStore[8][432]<=Wgt_8_432;WeightsStore[8][433]<=Wgt_8_433;WeightsStore[8][434]<=Wgt_8_434;WeightsStore[8][435]<=Wgt_8_435;WeightsStore[8][436]<=Wgt_8_436;WeightsStore[8][437]<=Wgt_8_437;WeightsStore[8][438]<=Wgt_8_438;WeightsStore[8][439]<=Wgt_8_439;WeightsStore[8][440]<=Wgt_8_440;WeightsStore[8][441]<=Wgt_8_441;WeightsStore[8][442]<=Wgt_8_442;WeightsStore[8][443]<=Wgt_8_443;WeightsStore[8][444]<=Wgt_8_444;WeightsStore[8][445]<=Wgt_8_445;WeightsStore[8][446]<=Wgt_8_446;WeightsStore[8][447]<=Wgt_8_447;WeightsStore[8][448]<=Wgt_8_448;WeightsStore[8][449]<=Wgt_8_449;WeightsStore[8][450]<=Wgt_8_450;WeightsStore[8][451]<=Wgt_8_451;WeightsStore[8][452]<=Wgt_8_452;WeightsStore[8][453]<=Wgt_8_453;WeightsStore[8][454]<=Wgt_8_454;WeightsStore[8][455]<=Wgt_8_455;WeightsStore[8][456]<=Wgt_8_456;WeightsStore[8][457]<=Wgt_8_457;WeightsStore[8][458]<=Wgt_8_458;WeightsStore[8][459]<=Wgt_8_459;WeightsStore[8][460]<=Wgt_8_460;WeightsStore[8][461]<=Wgt_8_461;WeightsStore[8][462]<=Wgt_8_462;WeightsStore[8][463]<=Wgt_8_463;WeightsStore[8][464]<=Wgt_8_464;WeightsStore[8][465]<=Wgt_8_465;WeightsStore[8][466]<=Wgt_8_466;WeightsStore[8][467]<=Wgt_8_467;WeightsStore[8][468]<=Wgt_8_468;WeightsStore[8][469]<=Wgt_8_469;WeightsStore[8][470]<=Wgt_8_470;WeightsStore[8][471]<=Wgt_8_471;WeightsStore[8][472]<=Wgt_8_472;WeightsStore[8][473]<=Wgt_8_473;WeightsStore[8][474]<=Wgt_8_474;WeightsStore[8][475]<=Wgt_8_475;WeightsStore[8][476]<=Wgt_8_476;WeightsStore[8][477]<=Wgt_8_477;WeightsStore[8][478]<=Wgt_8_478;WeightsStore[8][479]<=Wgt_8_479;WeightsStore[8][480]<=Wgt_8_480;WeightsStore[8][481]<=Wgt_8_481;WeightsStore[8][482]<=Wgt_8_482;WeightsStore[8][483]<=Wgt_8_483;WeightsStore[8][484]<=Wgt_8_484;WeightsStore[8][485]<=Wgt_8_485;WeightsStore[8][486]<=Wgt_8_486;WeightsStore[8][487]<=Wgt_8_487;WeightsStore[8][488]<=Wgt_8_488;WeightsStore[8][489]<=Wgt_8_489;WeightsStore[8][490]<=Wgt_8_490;WeightsStore[8][491]<=Wgt_8_491;WeightsStore[8][492]<=Wgt_8_492;WeightsStore[8][493]<=Wgt_8_493;WeightsStore[8][494]<=Wgt_8_494;WeightsStore[8][495]<=Wgt_8_495;WeightsStore[8][496]<=Wgt_8_496;WeightsStore[8][497]<=Wgt_8_497;WeightsStore[8][498]<=Wgt_8_498;WeightsStore[8][499]<=Wgt_8_499;WeightsStore[8][500]<=Wgt_8_500;WeightsStore[8][501]<=Wgt_8_501;WeightsStore[8][502]<=Wgt_8_502;WeightsStore[8][503]<=Wgt_8_503;WeightsStore[8][504]<=Wgt_8_504;WeightsStore[8][505]<=Wgt_8_505;WeightsStore[8][506]<=Wgt_8_506;WeightsStore[8][507]<=Wgt_8_507;WeightsStore[8][508]<=Wgt_8_508;WeightsStore[8][509]<=Wgt_8_509;WeightsStore[8][510]<=Wgt_8_510;WeightsStore[8][511]<=Wgt_8_511;WeightsStore[8][512]<=Wgt_8_512;WeightsStore[8][513]<=Wgt_8_513;WeightsStore[8][514]<=Wgt_8_514;WeightsStore[8][515]<=Wgt_8_515;WeightsStore[8][516]<=Wgt_8_516;WeightsStore[8][517]<=Wgt_8_517;WeightsStore[8][518]<=Wgt_8_518;WeightsStore[8][519]<=Wgt_8_519;WeightsStore[8][520]<=Wgt_8_520;WeightsStore[8][521]<=Wgt_8_521;WeightsStore[8][522]<=Wgt_8_522;WeightsStore[8][523]<=Wgt_8_523;WeightsStore[8][524]<=Wgt_8_524;WeightsStore[8][525]<=Wgt_8_525;WeightsStore[8][526]<=Wgt_8_526;WeightsStore[8][527]<=Wgt_8_527;WeightsStore[8][528]<=Wgt_8_528;WeightsStore[8][529]<=Wgt_8_529;WeightsStore[8][530]<=Wgt_8_530;WeightsStore[8][531]<=Wgt_8_531;WeightsStore[8][532]<=Wgt_8_532;WeightsStore[8][533]<=Wgt_8_533;WeightsStore[8][534]<=Wgt_8_534;WeightsStore[8][535]<=Wgt_8_535;WeightsStore[8][536]<=Wgt_8_536;WeightsStore[8][537]<=Wgt_8_537;WeightsStore[8][538]<=Wgt_8_538;WeightsStore[8][539]<=Wgt_8_539;WeightsStore[8][540]<=Wgt_8_540;WeightsStore[8][541]<=Wgt_8_541;WeightsStore[8][542]<=Wgt_8_542;WeightsStore[8][543]<=Wgt_8_543;WeightsStore[8][544]<=Wgt_8_544;WeightsStore[8][545]<=Wgt_8_545;WeightsStore[8][546]<=Wgt_8_546;WeightsStore[8][547]<=Wgt_8_547;WeightsStore[8][548]<=Wgt_8_548;WeightsStore[8][549]<=Wgt_8_549;WeightsStore[8][550]<=Wgt_8_550;WeightsStore[8][551]<=Wgt_8_551;WeightsStore[8][552]<=Wgt_8_552;WeightsStore[8][553]<=Wgt_8_553;WeightsStore[8][554]<=Wgt_8_554;WeightsStore[8][555]<=Wgt_8_555;WeightsStore[8][556]<=Wgt_8_556;WeightsStore[8][557]<=Wgt_8_557;WeightsStore[8][558]<=Wgt_8_558;WeightsStore[8][559]<=Wgt_8_559;WeightsStore[8][560]<=Wgt_8_560;WeightsStore[8][561]<=Wgt_8_561;WeightsStore[8][562]<=Wgt_8_562;WeightsStore[8][563]<=Wgt_8_563;WeightsStore[8][564]<=Wgt_8_564;WeightsStore[8][565]<=Wgt_8_565;WeightsStore[8][566]<=Wgt_8_566;WeightsStore[8][567]<=Wgt_8_567;WeightsStore[8][568]<=Wgt_8_568;WeightsStore[8][569]<=Wgt_8_569;WeightsStore[8][570]<=Wgt_8_570;WeightsStore[8][571]<=Wgt_8_571;WeightsStore[8][572]<=Wgt_8_572;WeightsStore[8][573]<=Wgt_8_573;WeightsStore[8][574]<=Wgt_8_574;WeightsStore[8][575]<=Wgt_8_575;WeightsStore[8][576]<=Wgt_8_576;WeightsStore[8][577]<=Wgt_8_577;WeightsStore[8][578]<=Wgt_8_578;WeightsStore[8][579]<=Wgt_8_579;WeightsStore[8][580]<=Wgt_8_580;WeightsStore[8][581]<=Wgt_8_581;WeightsStore[8][582]<=Wgt_8_582;WeightsStore[8][583]<=Wgt_8_583;WeightsStore[8][584]<=Wgt_8_584;WeightsStore[8][585]<=Wgt_8_585;WeightsStore[8][586]<=Wgt_8_586;WeightsStore[8][587]<=Wgt_8_587;WeightsStore[8][588]<=Wgt_8_588;WeightsStore[8][589]<=Wgt_8_589;WeightsStore[8][590]<=Wgt_8_590;WeightsStore[8][591]<=Wgt_8_591;WeightsStore[8][592]<=Wgt_8_592;WeightsStore[8][593]<=Wgt_8_593;WeightsStore[8][594]<=Wgt_8_594;WeightsStore[8][595]<=Wgt_8_595;WeightsStore[8][596]<=Wgt_8_596;WeightsStore[8][597]<=Wgt_8_597;WeightsStore[8][598]<=Wgt_8_598;WeightsStore[8][599]<=Wgt_8_599;WeightsStore[8][600]<=Wgt_8_600;WeightsStore[8][601]<=Wgt_8_601;WeightsStore[8][602]<=Wgt_8_602;WeightsStore[8][603]<=Wgt_8_603;WeightsStore[8][604]<=Wgt_8_604;WeightsStore[8][605]<=Wgt_8_605;WeightsStore[8][606]<=Wgt_8_606;WeightsStore[8][607]<=Wgt_8_607;WeightsStore[8][608]<=Wgt_8_608;WeightsStore[8][609]<=Wgt_8_609;WeightsStore[8][610]<=Wgt_8_610;WeightsStore[8][611]<=Wgt_8_611;WeightsStore[8][612]<=Wgt_8_612;WeightsStore[8][613]<=Wgt_8_613;WeightsStore[8][614]<=Wgt_8_614;WeightsStore[8][615]<=Wgt_8_615;WeightsStore[8][616]<=Wgt_8_616;WeightsStore[8][617]<=Wgt_8_617;WeightsStore[8][618]<=Wgt_8_618;WeightsStore[8][619]<=Wgt_8_619;WeightsStore[8][620]<=Wgt_8_620;WeightsStore[8][621]<=Wgt_8_621;WeightsStore[8][622]<=Wgt_8_622;WeightsStore[8][623]<=Wgt_8_623;WeightsStore[8][624]<=Wgt_8_624;WeightsStore[8][625]<=Wgt_8_625;WeightsStore[8][626]<=Wgt_8_626;WeightsStore[8][627]<=Wgt_8_627;WeightsStore[8][628]<=Wgt_8_628;WeightsStore[8][629]<=Wgt_8_629;WeightsStore[8][630]<=Wgt_8_630;WeightsStore[8][631]<=Wgt_8_631;WeightsStore[8][632]<=Wgt_8_632;WeightsStore[8][633]<=Wgt_8_633;WeightsStore[8][634]<=Wgt_8_634;WeightsStore[8][635]<=Wgt_8_635;WeightsStore[8][636]<=Wgt_8_636;WeightsStore[8][637]<=Wgt_8_637;WeightsStore[8][638]<=Wgt_8_638;WeightsStore[8][639]<=Wgt_8_639;WeightsStore[8][640]<=Wgt_8_640;WeightsStore[8][641]<=Wgt_8_641;WeightsStore[8][642]<=Wgt_8_642;WeightsStore[8][643]<=Wgt_8_643;WeightsStore[8][644]<=Wgt_8_644;WeightsStore[8][645]<=Wgt_8_645;WeightsStore[8][646]<=Wgt_8_646;WeightsStore[8][647]<=Wgt_8_647;WeightsStore[8][648]<=Wgt_8_648;WeightsStore[8][649]<=Wgt_8_649;WeightsStore[8][650]<=Wgt_8_650;WeightsStore[8][651]<=Wgt_8_651;WeightsStore[8][652]<=Wgt_8_652;WeightsStore[8][653]<=Wgt_8_653;WeightsStore[8][654]<=Wgt_8_654;WeightsStore[8][655]<=Wgt_8_655;WeightsStore[8][656]<=Wgt_8_656;WeightsStore[8][657]<=Wgt_8_657;WeightsStore[8][658]<=Wgt_8_658;WeightsStore[8][659]<=Wgt_8_659;WeightsStore[8][660]<=Wgt_8_660;WeightsStore[8][661]<=Wgt_8_661;WeightsStore[8][662]<=Wgt_8_662;WeightsStore[8][663]<=Wgt_8_663;WeightsStore[8][664]<=Wgt_8_664;WeightsStore[8][665]<=Wgt_8_665;WeightsStore[8][666]<=Wgt_8_666;WeightsStore[8][667]<=Wgt_8_667;WeightsStore[8][668]<=Wgt_8_668;WeightsStore[8][669]<=Wgt_8_669;WeightsStore[8][670]<=Wgt_8_670;WeightsStore[8][671]<=Wgt_8_671;WeightsStore[8][672]<=Wgt_8_672;WeightsStore[8][673]<=Wgt_8_673;WeightsStore[8][674]<=Wgt_8_674;WeightsStore[8][675]<=Wgt_8_675;WeightsStore[8][676]<=Wgt_8_676;WeightsStore[8][677]<=Wgt_8_677;WeightsStore[8][678]<=Wgt_8_678;WeightsStore[8][679]<=Wgt_8_679;WeightsStore[8][680]<=Wgt_8_680;WeightsStore[8][681]<=Wgt_8_681;WeightsStore[8][682]<=Wgt_8_682;WeightsStore[8][683]<=Wgt_8_683;WeightsStore[8][684]<=Wgt_8_684;WeightsStore[8][685]<=Wgt_8_685;WeightsStore[8][686]<=Wgt_8_686;WeightsStore[8][687]<=Wgt_8_687;WeightsStore[8][688]<=Wgt_8_688;WeightsStore[8][689]<=Wgt_8_689;WeightsStore[8][690]<=Wgt_8_690;WeightsStore[8][691]<=Wgt_8_691;WeightsStore[8][692]<=Wgt_8_692;WeightsStore[8][693]<=Wgt_8_693;WeightsStore[8][694]<=Wgt_8_694;WeightsStore[8][695]<=Wgt_8_695;WeightsStore[8][696]<=Wgt_8_696;WeightsStore[8][697]<=Wgt_8_697;WeightsStore[8][698]<=Wgt_8_698;WeightsStore[8][699]<=Wgt_8_699;WeightsStore[8][700]<=Wgt_8_700;WeightsStore[8][701]<=Wgt_8_701;WeightsStore[8][702]<=Wgt_8_702;WeightsStore[8][703]<=Wgt_8_703;WeightsStore[8][704]<=Wgt_8_704;WeightsStore[8][705]<=Wgt_8_705;WeightsStore[8][706]<=Wgt_8_706;WeightsStore[8][707]<=Wgt_8_707;WeightsStore[8][708]<=Wgt_8_708;WeightsStore[8][709]<=Wgt_8_709;WeightsStore[8][710]<=Wgt_8_710;WeightsStore[8][711]<=Wgt_8_711;WeightsStore[8][712]<=Wgt_8_712;WeightsStore[8][713]<=Wgt_8_713;WeightsStore[8][714]<=Wgt_8_714;WeightsStore[8][715]<=Wgt_8_715;WeightsStore[8][716]<=Wgt_8_716;WeightsStore[8][717]<=Wgt_8_717;WeightsStore[8][718]<=Wgt_8_718;WeightsStore[8][719]<=Wgt_8_719;WeightsStore[8][720]<=Wgt_8_720;WeightsStore[8][721]<=Wgt_8_721;WeightsStore[8][722]<=Wgt_8_722;WeightsStore[8][723]<=Wgt_8_723;WeightsStore[8][724]<=Wgt_8_724;WeightsStore[8][725]<=Wgt_8_725;WeightsStore[8][726]<=Wgt_8_726;WeightsStore[8][727]<=Wgt_8_727;WeightsStore[8][728]<=Wgt_8_728;WeightsStore[8][729]<=Wgt_8_729;WeightsStore[8][730]<=Wgt_8_730;WeightsStore[8][731]<=Wgt_8_731;WeightsStore[8][732]<=Wgt_8_732;WeightsStore[8][733]<=Wgt_8_733;WeightsStore[8][734]<=Wgt_8_734;WeightsStore[8][735]<=Wgt_8_735;WeightsStore[8][736]<=Wgt_8_736;WeightsStore[8][737]<=Wgt_8_737;WeightsStore[8][738]<=Wgt_8_738;WeightsStore[8][739]<=Wgt_8_739;WeightsStore[8][740]<=Wgt_8_740;WeightsStore[8][741]<=Wgt_8_741;WeightsStore[8][742]<=Wgt_8_742;WeightsStore[8][743]<=Wgt_8_743;WeightsStore[8][744]<=Wgt_8_744;WeightsStore[8][745]<=Wgt_8_745;WeightsStore[8][746]<=Wgt_8_746;WeightsStore[8][747]<=Wgt_8_747;WeightsStore[8][748]<=Wgt_8_748;WeightsStore[8][749]<=Wgt_8_749;WeightsStore[8][750]<=Wgt_8_750;WeightsStore[8][751]<=Wgt_8_751;WeightsStore[8][752]<=Wgt_8_752;WeightsStore[8][753]<=Wgt_8_753;WeightsStore[8][754]<=Wgt_8_754;WeightsStore[8][755]<=Wgt_8_755;WeightsStore[8][756]<=Wgt_8_756;WeightsStore[8][757]<=Wgt_8_757;WeightsStore[8][758]<=Wgt_8_758;WeightsStore[8][759]<=Wgt_8_759;WeightsStore[8][760]<=Wgt_8_760;WeightsStore[8][761]<=Wgt_8_761;WeightsStore[8][762]<=Wgt_8_762;WeightsStore[8][763]<=Wgt_8_763;WeightsStore[8][764]<=Wgt_8_764;WeightsStore[8][765]<=Wgt_8_765;WeightsStore[8][766]<=Wgt_8_766;WeightsStore[8][767]<=Wgt_8_767;WeightsStore[8][768]<=Wgt_8_768;WeightsStore[8][769]<=Wgt_8_769;WeightsStore[8][770]<=Wgt_8_770;WeightsStore[8][771]<=Wgt_8_771;WeightsStore[8][772]<=Wgt_8_772;WeightsStore[8][773]<=Wgt_8_773;WeightsStore[8][774]<=Wgt_8_774;WeightsStore[8][775]<=Wgt_8_775;WeightsStore[8][776]<=Wgt_8_776;WeightsStore[8][777]<=Wgt_8_777;WeightsStore[8][778]<=Wgt_8_778;WeightsStore[8][779]<=Wgt_8_779;WeightsStore[8][780]<=Wgt_8_780;WeightsStore[8][781]<=Wgt_8_781;WeightsStore[8][782]<=Wgt_8_782;WeightsStore[8][783]<=Wgt_8_783;WeightsStore[8][784]<=Wgt_8_784;WeightsStore[9][0]<=Wgt_9_0;WeightsStore[9][1]<=Wgt_9_1;WeightsStore[9][2]<=Wgt_9_2;WeightsStore[9][3]<=Wgt_9_3;WeightsStore[9][4]<=Wgt_9_4;WeightsStore[9][5]<=Wgt_9_5;WeightsStore[9][6]<=Wgt_9_6;WeightsStore[9][7]<=Wgt_9_7;WeightsStore[9][8]<=Wgt_9_8;WeightsStore[9][9]<=Wgt_9_9;WeightsStore[9][10]<=Wgt_9_10;WeightsStore[9][11]<=Wgt_9_11;WeightsStore[9][12]<=Wgt_9_12;WeightsStore[9][13]<=Wgt_9_13;WeightsStore[9][14]<=Wgt_9_14;WeightsStore[9][15]<=Wgt_9_15;WeightsStore[9][16]<=Wgt_9_16;WeightsStore[9][17]<=Wgt_9_17;WeightsStore[9][18]<=Wgt_9_18;WeightsStore[9][19]<=Wgt_9_19;WeightsStore[9][20]<=Wgt_9_20;WeightsStore[9][21]<=Wgt_9_21;WeightsStore[9][22]<=Wgt_9_22;WeightsStore[9][23]<=Wgt_9_23;WeightsStore[9][24]<=Wgt_9_24;WeightsStore[9][25]<=Wgt_9_25;WeightsStore[9][26]<=Wgt_9_26;WeightsStore[9][27]<=Wgt_9_27;WeightsStore[9][28]<=Wgt_9_28;WeightsStore[9][29]<=Wgt_9_29;WeightsStore[9][30]<=Wgt_9_30;WeightsStore[9][31]<=Wgt_9_31;WeightsStore[9][32]<=Wgt_9_32;WeightsStore[9][33]<=Wgt_9_33;WeightsStore[9][34]<=Wgt_9_34;WeightsStore[9][35]<=Wgt_9_35;WeightsStore[9][36]<=Wgt_9_36;WeightsStore[9][37]<=Wgt_9_37;WeightsStore[9][38]<=Wgt_9_38;WeightsStore[9][39]<=Wgt_9_39;WeightsStore[9][40]<=Wgt_9_40;WeightsStore[9][41]<=Wgt_9_41;WeightsStore[9][42]<=Wgt_9_42;WeightsStore[9][43]<=Wgt_9_43;WeightsStore[9][44]<=Wgt_9_44;WeightsStore[9][45]<=Wgt_9_45;WeightsStore[9][46]<=Wgt_9_46;WeightsStore[9][47]<=Wgt_9_47;WeightsStore[9][48]<=Wgt_9_48;WeightsStore[9][49]<=Wgt_9_49;WeightsStore[9][50]<=Wgt_9_50;WeightsStore[9][51]<=Wgt_9_51;WeightsStore[9][52]<=Wgt_9_52;WeightsStore[9][53]<=Wgt_9_53;WeightsStore[9][54]<=Wgt_9_54;WeightsStore[9][55]<=Wgt_9_55;WeightsStore[9][56]<=Wgt_9_56;WeightsStore[9][57]<=Wgt_9_57;WeightsStore[9][58]<=Wgt_9_58;WeightsStore[9][59]<=Wgt_9_59;WeightsStore[9][60]<=Wgt_9_60;WeightsStore[9][61]<=Wgt_9_61;WeightsStore[9][62]<=Wgt_9_62;WeightsStore[9][63]<=Wgt_9_63;WeightsStore[9][64]<=Wgt_9_64;WeightsStore[9][65]<=Wgt_9_65;WeightsStore[9][66]<=Wgt_9_66;WeightsStore[9][67]<=Wgt_9_67;WeightsStore[9][68]<=Wgt_9_68;WeightsStore[9][69]<=Wgt_9_69;WeightsStore[9][70]<=Wgt_9_70;WeightsStore[9][71]<=Wgt_9_71;WeightsStore[9][72]<=Wgt_9_72;WeightsStore[9][73]<=Wgt_9_73;WeightsStore[9][74]<=Wgt_9_74;WeightsStore[9][75]<=Wgt_9_75;WeightsStore[9][76]<=Wgt_9_76;WeightsStore[9][77]<=Wgt_9_77;WeightsStore[9][78]<=Wgt_9_78;WeightsStore[9][79]<=Wgt_9_79;WeightsStore[9][80]<=Wgt_9_80;WeightsStore[9][81]<=Wgt_9_81;WeightsStore[9][82]<=Wgt_9_82;WeightsStore[9][83]<=Wgt_9_83;WeightsStore[9][84]<=Wgt_9_84;WeightsStore[9][85]<=Wgt_9_85;WeightsStore[9][86]<=Wgt_9_86;WeightsStore[9][87]<=Wgt_9_87;WeightsStore[9][88]<=Wgt_9_88;WeightsStore[9][89]<=Wgt_9_89;WeightsStore[9][90]<=Wgt_9_90;WeightsStore[9][91]<=Wgt_9_91;WeightsStore[9][92]<=Wgt_9_92;WeightsStore[9][93]<=Wgt_9_93;WeightsStore[9][94]<=Wgt_9_94;WeightsStore[9][95]<=Wgt_9_95;WeightsStore[9][96]<=Wgt_9_96;WeightsStore[9][97]<=Wgt_9_97;WeightsStore[9][98]<=Wgt_9_98;WeightsStore[9][99]<=Wgt_9_99;WeightsStore[9][100]<=Wgt_9_100;WeightsStore[9][101]<=Wgt_9_101;WeightsStore[9][102]<=Wgt_9_102;WeightsStore[9][103]<=Wgt_9_103;WeightsStore[9][104]<=Wgt_9_104;WeightsStore[9][105]<=Wgt_9_105;WeightsStore[9][106]<=Wgt_9_106;WeightsStore[9][107]<=Wgt_9_107;WeightsStore[9][108]<=Wgt_9_108;WeightsStore[9][109]<=Wgt_9_109;WeightsStore[9][110]<=Wgt_9_110;WeightsStore[9][111]<=Wgt_9_111;WeightsStore[9][112]<=Wgt_9_112;WeightsStore[9][113]<=Wgt_9_113;WeightsStore[9][114]<=Wgt_9_114;WeightsStore[9][115]<=Wgt_9_115;WeightsStore[9][116]<=Wgt_9_116;WeightsStore[9][117]<=Wgt_9_117;WeightsStore[9][118]<=Wgt_9_118;WeightsStore[9][119]<=Wgt_9_119;WeightsStore[9][120]<=Wgt_9_120;WeightsStore[9][121]<=Wgt_9_121;WeightsStore[9][122]<=Wgt_9_122;WeightsStore[9][123]<=Wgt_9_123;WeightsStore[9][124]<=Wgt_9_124;WeightsStore[9][125]<=Wgt_9_125;WeightsStore[9][126]<=Wgt_9_126;WeightsStore[9][127]<=Wgt_9_127;WeightsStore[9][128]<=Wgt_9_128;WeightsStore[9][129]<=Wgt_9_129;WeightsStore[9][130]<=Wgt_9_130;WeightsStore[9][131]<=Wgt_9_131;WeightsStore[9][132]<=Wgt_9_132;WeightsStore[9][133]<=Wgt_9_133;WeightsStore[9][134]<=Wgt_9_134;WeightsStore[9][135]<=Wgt_9_135;WeightsStore[9][136]<=Wgt_9_136;WeightsStore[9][137]<=Wgt_9_137;WeightsStore[9][138]<=Wgt_9_138;WeightsStore[9][139]<=Wgt_9_139;WeightsStore[9][140]<=Wgt_9_140;WeightsStore[9][141]<=Wgt_9_141;WeightsStore[9][142]<=Wgt_9_142;WeightsStore[9][143]<=Wgt_9_143;WeightsStore[9][144]<=Wgt_9_144;WeightsStore[9][145]<=Wgt_9_145;WeightsStore[9][146]<=Wgt_9_146;WeightsStore[9][147]<=Wgt_9_147;WeightsStore[9][148]<=Wgt_9_148;WeightsStore[9][149]<=Wgt_9_149;WeightsStore[9][150]<=Wgt_9_150;WeightsStore[9][151]<=Wgt_9_151;WeightsStore[9][152]<=Wgt_9_152;WeightsStore[9][153]<=Wgt_9_153;WeightsStore[9][154]<=Wgt_9_154;WeightsStore[9][155]<=Wgt_9_155;WeightsStore[9][156]<=Wgt_9_156;WeightsStore[9][157]<=Wgt_9_157;WeightsStore[9][158]<=Wgt_9_158;WeightsStore[9][159]<=Wgt_9_159;WeightsStore[9][160]<=Wgt_9_160;WeightsStore[9][161]<=Wgt_9_161;WeightsStore[9][162]<=Wgt_9_162;WeightsStore[9][163]<=Wgt_9_163;WeightsStore[9][164]<=Wgt_9_164;WeightsStore[9][165]<=Wgt_9_165;WeightsStore[9][166]<=Wgt_9_166;WeightsStore[9][167]<=Wgt_9_167;WeightsStore[9][168]<=Wgt_9_168;WeightsStore[9][169]<=Wgt_9_169;WeightsStore[9][170]<=Wgt_9_170;WeightsStore[9][171]<=Wgt_9_171;WeightsStore[9][172]<=Wgt_9_172;WeightsStore[9][173]<=Wgt_9_173;WeightsStore[9][174]<=Wgt_9_174;WeightsStore[9][175]<=Wgt_9_175;WeightsStore[9][176]<=Wgt_9_176;WeightsStore[9][177]<=Wgt_9_177;WeightsStore[9][178]<=Wgt_9_178;WeightsStore[9][179]<=Wgt_9_179;WeightsStore[9][180]<=Wgt_9_180;WeightsStore[9][181]<=Wgt_9_181;WeightsStore[9][182]<=Wgt_9_182;WeightsStore[9][183]<=Wgt_9_183;WeightsStore[9][184]<=Wgt_9_184;WeightsStore[9][185]<=Wgt_9_185;WeightsStore[9][186]<=Wgt_9_186;WeightsStore[9][187]<=Wgt_9_187;WeightsStore[9][188]<=Wgt_9_188;WeightsStore[9][189]<=Wgt_9_189;WeightsStore[9][190]<=Wgt_9_190;WeightsStore[9][191]<=Wgt_9_191;WeightsStore[9][192]<=Wgt_9_192;WeightsStore[9][193]<=Wgt_9_193;WeightsStore[9][194]<=Wgt_9_194;WeightsStore[9][195]<=Wgt_9_195;WeightsStore[9][196]<=Wgt_9_196;WeightsStore[9][197]<=Wgt_9_197;WeightsStore[9][198]<=Wgt_9_198;WeightsStore[9][199]<=Wgt_9_199;WeightsStore[9][200]<=Wgt_9_200;WeightsStore[9][201]<=Wgt_9_201;WeightsStore[9][202]<=Wgt_9_202;WeightsStore[9][203]<=Wgt_9_203;WeightsStore[9][204]<=Wgt_9_204;WeightsStore[9][205]<=Wgt_9_205;WeightsStore[9][206]<=Wgt_9_206;WeightsStore[9][207]<=Wgt_9_207;WeightsStore[9][208]<=Wgt_9_208;WeightsStore[9][209]<=Wgt_9_209;WeightsStore[9][210]<=Wgt_9_210;WeightsStore[9][211]<=Wgt_9_211;WeightsStore[9][212]<=Wgt_9_212;WeightsStore[9][213]<=Wgt_9_213;WeightsStore[9][214]<=Wgt_9_214;WeightsStore[9][215]<=Wgt_9_215;WeightsStore[9][216]<=Wgt_9_216;WeightsStore[9][217]<=Wgt_9_217;WeightsStore[9][218]<=Wgt_9_218;WeightsStore[9][219]<=Wgt_9_219;WeightsStore[9][220]<=Wgt_9_220;WeightsStore[9][221]<=Wgt_9_221;WeightsStore[9][222]<=Wgt_9_222;WeightsStore[9][223]<=Wgt_9_223;WeightsStore[9][224]<=Wgt_9_224;WeightsStore[9][225]<=Wgt_9_225;WeightsStore[9][226]<=Wgt_9_226;WeightsStore[9][227]<=Wgt_9_227;WeightsStore[9][228]<=Wgt_9_228;WeightsStore[9][229]<=Wgt_9_229;WeightsStore[9][230]<=Wgt_9_230;WeightsStore[9][231]<=Wgt_9_231;WeightsStore[9][232]<=Wgt_9_232;WeightsStore[9][233]<=Wgt_9_233;WeightsStore[9][234]<=Wgt_9_234;WeightsStore[9][235]<=Wgt_9_235;WeightsStore[9][236]<=Wgt_9_236;WeightsStore[9][237]<=Wgt_9_237;WeightsStore[9][238]<=Wgt_9_238;WeightsStore[9][239]<=Wgt_9_239;WeightsStore[9][240]<=Wgt_9_240;WeightsStore[9][241]<=Wgt_9_241;WeightsStore[9][242]<=Wgt_9_242;WeightsStore[9][243]<=Wgt_9_243;WeightsStore[9][244]<=Wgt_9_244;WeightsStore[9][245]<=Wgt_9_245;WeightsStore[9][246]<=Wgt_9_246;WeightsStore[9][247]<=Wgt_9_247;WeightsStore[9][248]<=Wgt_9_248;WeightsStore[9][249]<=Wgt_9_249;WeightsStore[9][250]<=Wgt_9_250;WeightsStore[9][251]<=Wgt_9_251;WeightsStore[9][252]<=Wgt_9_252;WeightsStore[9][253]<=Wgt_9_253;WeightsStore[9][254]<=Wgt_9_254;WeightsStore[9][255]<=Wgt_9_255;WeightsStore[9][256]<=Wgt_9_256;WeightsStore[9][257]<=Wgt_9_257;WeightsStore[9][258]<=Wgt_9_258;WeightsStore[9][259]<=Wgt_9_259;WeightsStore[9][260]<=Wgt_9_260;WeightsStore[9][261]<=Wgt_9_261;WeightsStore[9][262]<=Wgt_9_262;WeightsStore[9][263]<=Wgt_9_263;WeightsStore[9][264]<=Wgt_9_264;WeightsStore[9][265]<=Wgt_9_265;WeightsStore[9][266]<=Wgt_9_266;WeightsStore[9][267]<=Wgt_9_267;WeightsStore[9][268]<=Wgt_9_268;WeightsStore[9][269]<=Wgt_9_269;WeightsStore[9][270]<=Wgt_9_270;WeightsStore[9][271]<=Wgt_9_271;WeightsStore[9][272]<=Wgt_9_272;WeightsStore[9][273]<=Wgt_9_273;WeightsStore[9][274]<=Wgt_9_274;WeightsStore[9][275]<=Wgt_9_275;WeightsStore[9][276]<=Wgt_9_276;WeightsStore[9][277]<=Wgt_9_277;WeightsStore[9][278]<=Wgt_9_278;WeightsStore[9][279]<=Wgt_9_279;WeightsStore[9][280]<=Wgt_9_280;WeightsStore[9][281]<=Wgt_9_281;WeightsStore[9][282]<=Wgt_9_282;WeightsStore[9][283]<=Wgt_9_283;WeightsStore[9][284]<=Wgt_9_284;WeightsStore[9][285]<=Wgt_9_285;WeightsStore[9][286]<=Wgt_9_286;WeightsStore[9][287]<=Wgt_9_287;WeightsStore[9][288]<=Wgt_9_288;WeightsStore[9][289]<=Wgt_9_289;WeightsStore[9][290]<=Wgt_9_290;WeightsStore[9][291]<=Wgt_9_291;WeightsStore[9][292]<=Wgt_9_292;WeightsStore[9][293]<=Wgt_9_293;WeightsStore[9][294]<=Wgt_9_294;WeightsStore[9][295]<=Wgt_9_295;WeightsStore[9][296]<=Wgt_9_296;WeightsStore[9][297]<=Wgt_9_297;WeightsStore[9][298]<=Wgt_9_298;WeightsStore[9][299]<=Wgt_9_299;WeightsStore[9][300]<=Wgt_9_300;WeightsStore[9][301]<=Wgt_9_301;WeightsStore[9][302]<=Wgt_9_302;WeightsStore[9][303]<=Wgt_9_303;WeightsStore[9][304]<=Wgt_9_304;WeightsStore[9][305]<=Wgt_9_305;WeightsStore[9][306]<=Wgt_9_306;WeightsStore[9][307]<=Wgt_9_307;WeightsStore[9][308]<=Wgt_9_308;WeightsStore[9][309]<=Wgt_9_309;WeightsStore[9][310]<=Wgt_9_310;WeightsStore[9][311]<=Wgt_9_311;WeightsStore[9][312]<=Wgt_9_312;WeightsStore[9][313]<=Wgt_9_313;WeightsStore[9][314]<=Wgt_9_314;WeightsStore[9][315]<=Wgt_9_315;WeightsStore[9][316]<=Wgt_9_316;WeightsStore[9][317]<=Wgt_9_317;WeightsStore[9][318]<=Wgt_9_318;WeightsStore[9][319]<=Wgt_9_319;WeightsStore[9][320]<=Wgt_9_320;WeightsStore[9][321]<=Wgt_9_321;WeightsStore[9][322]<=Wgt_9_322;WeightsStore[9][323]<=Wgt_9_323;WeightsStore[9][324]<=Wgt_9_324;WeightsStore[9][325]<=Wgt_9_325;WeightsStore[9][326]<=Wgt_9_326;WeightsStore[9][327]<=Wgt_9_327;WeightsStore[9][328]<=Wgt_9_328;WeightsStore[9][329]<=Wgt_9_329;WeightsStore[9][330]<=Wgt_9_330;WeightsStore[9][331]<=Wgt_9_331;WeightsStore[9][332]<=Wgt_9_332;WeightsStore[9][333]<=Wgt_9_333;WeightsStore[9][334]<=Wgt_9_334;WeightsStore[9][335]<=Wgt_9_335;WeightsStore[9][336]<=Wgt_9_336;WeightsStore[9][337]<=Wgt_9_337;WeightsStore[9][338]<=Wgt_9_338;WeightsStore[9][339]<=Wgt_9_339;WeightsStore[9][340]<=Wgt_9_340;WeightsStore[9][341]<=Wgt_9_341;WeightsStore[9][342]<=Wgt_9_342;WeightsStore[9][343]<=Wgt_9_343;WeightsStore[9][344]<=Wgt_9_344;WeightsStore[9][345]<=Wgt_9_345;WeightsStore[9][346]<=Wgt_9_346;WeightsStore[9][347]<=Wgt_9_347;WeightsStore[9][348]<=Wgt_9_348;WeightsStore[9][349]<=Wgt_9_349;WeightsStore[9][350]<=Wgt_9_350;WeightsStore[9][351]<=Wgt_9_351;WeightsStore[9][352]<=Wgt_9_352;WeightsStore[9][353]<=Wgt_9_353;WeightsStore[9][354]<=Wgt_9_354;WeightsStore[9][355]<=Wgt_9_355;WeightsStore[9][356]<=Wgt_9_356;WeightsStore[9][357]<=Wgt_9_357;WeightsStore[9][358]<=Wgt_9_358;WeightsStore[9][359]<=Wgt_9_359;WeightsStore[9][360]<=Wgt_9_360;WeightsStore[9][361]<=Wgt_9_361;WeightsStore[9][362]<=Wgt_9_362;WeightsStore[9][363]<=Wgt_9_363;WeightsStore[9][364]<=Wgt_9_364;WeightsStore[9][365]<=Wgt_9_365;WeightsStore[9][366]<=Wgt_9_366;WeightsStore[9][367]<=Wgt_9_367;WeightsStore[9][368]<=Wgt_9_368;WeightsStore[9][369]<=Wgt_9_369;WeightsStore[9][370]<=Wgt_9_370;WeightsStore[9][371]<=Wgt_9_371;WeightsStore[9][372]<=Wgt_9_372;WeightsStore[9][373]<=Wgt_9_373;WeightsStore[9][374]<=Wgt_9_374;WeightsStore[9][375]<=Wgt_9_375;WeightsStore[9][376]<=Wgt_9_376;WeightsStore[9][377]<=Wgt_9_377;WeightsStore[9][378]<=Wgt_9_378;WeightsStore[9][379]<=Wgt_9_379;WeightsStore[9][380]<=Wgt_9_380;WeightsStore[9][381]<=Wgt_9_381;WeightsStore[9][382]<=Wgt_9_382;WeightsStore[9][383]<=Wgt_9_383;WeightsStore[9][384]<=Wgt_9_384;WeightsStore[9][385]<=Wgt_9_385;WeightsStore[9][386]<=Wgt_9_386;WeightsStore[9][387]<=Wgt_9_387;WeightsStore[9][388]<=Wgt_9_388;WeightsStore[9][389]<=Wgt_9_389;WeightsStore[9][390]<=Wgt_9_390;WeightsStore[9][391]<=Wgt_9_391;WeightsStore[9][392]<=Wgt_9_392;WeightsStore[9][393]<=Wgt_9_393;WeightsStore[9][394]<=Wgt_9_394;WeightsStore[9][395]<=Wgt_9_395;WeightsStore[9][396]<=Wgt_9_396;WeightsStore[9][397]<=Wgt_9_397;WeightsStore[9][398]<=Wgt_9_398;WeightsStore[9][399]<=Wgt_9_399;WeightsStore[9][400]<=Wgt_9_400;WeightsStore[9][401]<=Wgt_9_401;WeightsStore[9][402]<=Wgt_9_402;WeightsStore[9][403]<=Wgt_9_403;WeightsStore[9][404]<=Wgt_9_404;WeightsStore[9][405]<=Wgt_9_405;WeightsStore[9][406]<=Wgt_9_406;WeightsStore[9][407]<=Wgt_9_407;WeightsStore[9][408]<=Wgt_9_408;WeightsStore[9][409]<=Wgt_9_409;WeightsStore[9][410]<=Wgt_9_410;WeightsStore[9][411]<=Wgt_9_411;WeightsStore[9][412]<=Wgt_9_412;WeightsStore[9][413]<=Wgt_9_413;WeightsStore[9][414]<=Wgt_9_414;WeightsStore[9][415]<=Wgt_9_415;WeightsStore[9][416]<=Wgt_9_416;WeightsStore[9][417]<=Wgt_9_417;WeightsStore[9][418]<=Wgt_9_418;WeightsStore[9][419]<=Wgt_9_419;WeightsStore[9][420]<=Wgt_9_420;WeightsStore[9][421]<=Wgt_9_421;WeightsStore[9][422]<=Wgt_9_422;WeightsStore[9][423]<=Wgt_9_423;WeightsStore[9][424]<=Wgt_9_424;WeightsStore[9][425]<=Wgt_9_425;WeightsStore[9][426]<=Wgt_9_426;WeightsStore[9][427]<=Wgt_9_427;WeightsStore[9][428]<=Wgt_9_428;WeightsStore[9][429]<=Wgt_9_429;WeightsStore[9][430]<=Wgt_9_430;WeightsStore[9][431]<=Wgt_9_431;WeightsStore[9][432]<=Wgt_9_432;WeightsStore[9][433]<=Wgt_9_433;WeightsStore[9][434]<=Wgt_9_434;WeightsStore[9][435]<=Wgt_9_435;WeightsStore[9][436]<=Wgt_9_436;WeightsStore[9][437]<=Wgt_9_437;WeightsStore[9][438]<=Wgt_9_438;WeightsStore[9][439]<=Wgt_9_439;WeightsStore[9][440]<=Wgt_9_440;WeightsStore[9][441]<=Wgt_9_441;WeightsStore[9][442]<=Wgt_9_442;WeightsStore[9][443]<=Wgt_9_443;WeightsStore[9][444]<=Wgt_9_444;WeightsStore[9][445]<=Wgt_9_445;WeightsStore[9][446]<=Wgt_9_446;WeightsStore[9][447]<=Wgt_9_447;WeightsStore[9][448]<=Wgt_9_448;WeightsStore[9][449]<=Wgt_9_449;WeightsStore[9][450]<=Wgt_9_450;WeightsStore[9][451]<=Wgt_9_451;WeightsStore[9][452]<=Wgt_9_452;WeightsStore[9][453]<=Wgt_9_453;WeightsStore[9][454]<=Wgt_9_454;WeightsStore[9][455]<=Wgt_9_455;WeightsStore[9][456]<=Wgt_9_456;WeightsStore[9][457]<=Wgt_9_457;WeightsStore[9][458]<=Wgt_9_458;WeightsStore[9][459]<=Wgt_9_459;WeightsStore[9][460]<=Wgt_9_460;WeightsStore[9][461]<=Wgt_9_461;WeightsStore[9][462]<=Wgt_9_462;WeightsStore[9][463]<=Wgt_9_463;WeightsStore[9][464]<=Wgt_9_464;WeightsStore[9][465]<=Wgt_9_465;WeightsStore[9][466]<=Wgt_9_466;WeightsStore[9][467]<=Wgt_9_467;WeightsStore[9][468]<=Wgt_9_468;WeightsStore[9][469]<=Wgt_9_469;WeightsStore[9][470]<=Wgt_9_470;WeightsStore[9][471]<=Wgt_9_471;WeightsStore[9][472]<=Wgt_9_472;WeightsStore[9][473]<=Wgt_9_473;WeightsStore[9][474]<=Wgt_9_474;WeightsStore[9][475]<=Wgt_9_475;WeightsStore[9][476]<=Wgt_9_476;WeightsStore[9][477]<=Wgt_9_477;WeightsStore[9][478]<=Wgt_9_478;WeightsStore[9][479]<=Wgt_9_479;WeightsStore[9][480]<=Wgt_9_480;WeightsStore[9][481]<=Wgt_9_481;WeightsStore[9][482]<=Wgt_9_482;WeightsStore[9][483]<=Wgt_9_483;WeightsStore[9][484]<=Wgt_9_484;WeightsStore[9][485]<=Wgt_9_485;WeightsStore[9][486]<=Wgt_9_486;WeightsStore[9][487]<=Wgt_9_487;WeightsStore[9][488]<=Wgt_9_488;WeightsStore[9][489]<=Wgt_9_489;WeightsStore[9][490]<=Wgt_9_490;WeightsStore[9][491]<=Wgt_9_491;WeightsStore[9][492]<=Wgt_9_492;WeightsStore[9][493]<=Wgt_9_493;WeightsStore[9][494]<=Wgt_9_494;WeightsStore[9][495]<=Wgt_9_495;WeightsStore[9][496]<=Wgt_9_496;WeightsStore[9][497]<=Wgt_9_497;WeightsStore[9][498]<=Wgt_9_498;WeightsStore[9][499]<=Wgt_9_499;WeightsStore[9][500]<=Wgt_9_500;WeightsStore[9][501]<=Wgt_9_501;WeightsStore[9][502]<=Wgt_9_502;WeightsStore[9][503]<=Wgt_9_503;WeightsStore[9][504]<=Wgt_9_504;WeightsStore[9][505]<=Wgt_9_505;WeightsStore[9][506]<=Wgt_9_506;WeightsStore[9][507]<=Wgt_9_507;WeightsStore[9][508]<=Wgt_9_508;WeightsStore[9][509]<=Wgt_9_509;WeightsStore[9][510]<=Wgt_9_510;WeightsStore[9][511]<=Wgt_9_511;WeightsStore[9][512]<=Wgt_9_512;WeightsStore[9][513]<=Wgt_9_513;WeightsStore[9][514]<=Wgt_9_514;WeightsStore[9][515]<=Wgt_9_515;WeightsStore[9][516]<=Wgt_9_516;WeightsStore[9][517]<=Wgt_9_517;WeightsStore[9][518]<=Wgt_9_518;WeightsStore[9][519]<=Wgt_9_519;WeightsStore[9][520]<=Wgt_9_520;WeightsStore[9][521]<=Wgt_9_521;WeightsStore[9][522]<=Wgt_9_522;WeightsStore[9][523]<=Wgt_9_523;WeightsStore[9][524]<=Wgt_9_524;WeightsStore[9][525]<=Wgt_9_525;WeightsStore[9][526]<=Wgt_9_526;WeightsStore[9][527]<=Wgt_9_527;WeightsStore[9][528]<=Wgt_9_528;WeightsStore[9][529]<=Wgt_9_529;WeightsStore[9][530]<=Wgt_9_530;WeightsStore[9][531]<=Wgt_9_531;WeightsStore[9][532]<=Wgt_9_532;WeightsStore[9][533]<=Wgt_9_533;WeightsStore[9][534]<=Wgt_9_534;WeightsStore[9][535]<=Wgt_9_535;WeightsStore[9][536]<=Wgt_9_536;WeightsStore[9][537]<=Wgt_9_537;WeightsStore[9][538]<=Wgt_9_538;WeightsStore[9][539]<=Wgt_9_539;WeightsStore[9][540]<=Wgt_9_540;WeightsStore[9][541]<=Wgt_9_541;WeightsStore[9][542]<=Wgt_9_542;WeightsStore[9][543]<=Wgt_9_543;WeightsStore[9][544]<=Wgt_9_544;WeightsStore[9][545]<=Wgt_9_545;WeightsStore[9][546]<=Wgt_9_546;WeightsStore[9][547]<=Wgt_9_547;WeightsStore[9][548]<=Wgt_9_548;WeightsStore[9][549]<=Wgt_9_549;WeightsStore[9][550]<=Wgt_9_550;WeightsStore[9][551]<=Wgt_9_551;WeightsStore[9][552]<=Wgt_9_552;WeightsStore[9][553]<=Wgt_9_553;WeightsStore[9][554]<=Wgt_9_554;WeightsStore[9][555]<=Wgt_9_555;WeightsStore[9][556]<=Wgt_9_556;WeightsStore[9][557]<=Wgt_9_557;WeightsStore[9][558]<=Wgt_9_558;WeightsStore[9][559]<=Wgt_9_559;WeightsStore[9][560]<=Wgt_9_560;WeightsStore[9][561]<=Wgt_9_561;WeightsStore[9][562]<=Wgt_9_562;WeightsStore[9][563]<=Wgt_9_563;WeightsStore[9][564]<=Wgt_9_564;WeightsStore[9][565]<=Wgt_9_565;WeightsStore[9][566]<=Wgt_9_566;WeightsStore[9][567]<=Wgt_9_567;WeightsStore[9][568]<=Wgt_9_568;WeightsStore[9][569]<=Wgt_9_569;WeightsStore[9][570]<=Wgt_9_570;WeightsStore[9][571]<=Wgt_9_571;WeightsStore[9][572]<=Wgt_9_572;WeightsStore[9][573]<=Wgt_9_573;WeightsStore[9][574]<=Wgt_9_574;WeightsStore[9][575]<=Wgt_9_575;WeightsStore[9][576]<=Wgt_9_576;WeightsStore[9][577]<=Wgt_9_577;WeightsStore[9][578]<=Wgt_9_578;WeightsStore[9][579]<=Wgt_9_579;WeightsStore[9][580]<=Wgt_9_580;WeightsStore[9][581]<=Wgt_9_581;WeightsStore[9][582]<=Wgt_9_582;WeightsStore[9][583]<=Wgt_9_583;WeightsStore[9][584]<=Wgt_9_584;WeightsStore[9][585]<=Wgt_9_585;WeightsStore[9][586]<=Wgt_9_586;WeightsStore[9][587]<=Wgt_9_587;WeightsStore[9][588]<=Wgt_9_588;WeightsStore[9][589]<=Wgt_9_589;WeightsStore[9][590]<=Wgt_9_590;WeightsStore[9][591]<=Wgt_9_591;WeightsStore[9][592]<=Wgt_9_592;WeightsStore[9][593]<=Wgt_9_593;WeightsStore[9][594]<=Wgt_9_594;WeightsStore[9][595]<=Wgt_9_595;WeightsStore[9][596]<=Wgt_9_596;WeightsStore[9][597]<=Wgt_9_597;WeightsStore[9][598]<=Wgt_9_598;WeightsStore[9][599]<=Wgt_9_599;WeightsStore[9][600]<=Wgt_9_600;WeightsStore[9][601]<=Wgt_9_601;WeightsStore[9][602]<=Wgt_9_602;WeightsStore[9][603]<=Wgt_9_603;WeightsStore[9][604]<=Wgt_9_604;WeightsStore[9][605]<=Wgt_9_605;WeightsStore[9][606]<=Wgt_9_606;WeightsStore[9][607]<=Wgt_9_607;WeightsStore[9][608]<=Wgt_9_608;WeightsStore[9][609]<=Wgt_9_609;WeightsStore[9][610]<=Wgt_9_610;WeightsStore[9][611]<=Wgt_9_611;WeightsStore[9][612]<=Wgt_9_612;WeightsStore[9][613]<=Wgt_9_613;WeightsStore[9][614]<=Wgt_9_614;WeightsStore[9][615]<=Wgt_9_615;WeightsStore[9][616]<=Wgt_9_616;WeightsStore[9][617]<=Wgt_9_617;WeightsStore[9][618]<=Wgt_9_618;WeightsStore[9][619]<=Wgt_9_619;WeightsStore[9][620]<=Wgt_9_620;WeightsStore[9][621]<=Wgt_9_621;WeightsStore[9][622]<=Wgt_9_622;WeightsStore[9][623]<=Wgt_9_623;WeightsStore[9][624]<=Wgt_9_624;WeightsStore[9][625]<=Wgt_9_625;WeightsStore[9][626]<=Wgt_9_626;WeightsStore[9][627]<=Wgt_9_627;WeightsStore[9][628]<=Wgt_9_628;WeightsStore[9][629]<=Wgt_9_629;WeightsStore[9][630]<=Wgt_9_630;WeightsStore[9][631]<=Wgt_9_631;WeightsStore[9][632]<=Wgt_9_632;WeightsStore[9][633]<=Wgt_9_633;WeightsStore[9][634]<=Wgt_9_634;WeightsStore[9][635]<=Wgt_9_635;WeightsStore[9][636]<=Wgt_9_636;WeightsStore[9][637]<=Wgt_9_637;WeightsStore[9][638]<=Wgt_9_638;WeightsStore[9][639]<=Wgt_9_639;WeightsStore[9][640]<=Wgt_9_640;WeightsStore[9][641]<=Wgt_9_641;WeightsStore[9][642]<=Wgt_9_642;WeightsStore[9][643]<=Wgt_9_643;WeightsStore[9][644]<=Wgt_9_644;WeightsStore[9][645]<=Wgt_9_645;WeightsStore[9][646]<=Wgt_9_646;WeightsStore[9][647]<=Wgt_9_647;WeightsStore[9][648]<=Wgt_9_648;WeightsStore[9][649]<=Wgt_9_649;WeightsStore[9][650]<=Wgt_9_650;WeightsStore[9][651]<=Wgt_9_651;WeightsStore[9][652]<=Wgt_9_652;WeightsStore[9][653]<=Wgt_9_653;WeightsStore[9][654]<=Wgt_9_654;WeightsStore[9][655]<=Wgt_9_655;WeightsStore[9][656]<=Wgt_9_656;WeightsStore[9][657]<=Wgt_9_657;WeightsStore[9][658]<=Wgt_9_658;WeightsStore[9][659]<=Wgt_9_659;WeightsStore[9][660]<=Wgt_9_660;WeightsStore[9][661]<=Wgt_9_661;WeightsStore[9][662]<=Wgt_9_662;WeightsStore[9][663]<=Wgt_9_663;WeightsStore[9][664]<=Wgt_9_664;WeightsStore[9][665]<=Wgt_9_665;WeightsStore[9][666]<=Wgt_9_666;WeightsStore[9][667]<=Wgt_9_667;WeightsStore[9][668]<=Wgt_9_668;WeightsStore[9][669]<=Wgt_9_669;WeightsStore[9][670]<=Wgt_9_670;WeightsStore[9][671]<=Wgt_9_671;WeightsStore[9][672]<=Wgt_9_672;WeightsStore[9][673]<=Wgt_9_673;WeightsStore[9][674]<=Wgt_9_674;WeightsStore[9][675]<=Wgt_9_675;WeightsStore[9][676]<=Wgt_9_676;WeightsStore[9][677]<=Wgt_9_677;WeightsStore[9][678]<=Wgt_9_678;WeightsStore[9][679]<=Wgt_9_679;WeightsStore[9][680]<=Wgt_9_680;WeightsStore[9][681]<=Wgt_9_681;WeightsStore[9][682]<=Wgt_9_682;WeightsStore[9][683]<=Wgt_9_683;WeightsStore[9][684]<=Wgt_9_684;WeightsStore[9][685]<=Wgt_9_685;WeightsStore[9][686]<=Wgt_9_686;WeightsStore[9][687]<=Wgt_9_687;WeightsStore[9][688]<=Wgt_9_688;WeightsStore[9][689]<=Wgt_9_689;WeightsStore[9][690]<=Wgt_9_690;WeightsStore[9][691]<=Wgt_9_691;WeightsStore[9][692]<=Wgt_9_692;WeightsStore[9][693]<=Wgt_9_693;WeightsStore[9][694]<=Wgt_9_694;WeightsStore[9][695]<=Wgt_9_695;WeightsStore[9][696]<=Wgt_9_696;WeightsStore[9][697]<=Wgt_9_697;WeightsStore[9][698]<=Wgt_9_698;WeightsStore[9][699]<=Wgt_9_699;WeightsStore[9][700]<=Wgt_9_700;WeightsStore[9][701]<=Wgt_9_701;WeightsStore[9][702]<=Wgt_9_702;WeightsStore[9][703]<=Wgt_9_703;WeightsStore[9][704]<=Wgt_9_704;WeightsStore[9][705]<=Wgt_9_705;WeightsStore[9][706]<=Wgt_9_706;WeightsStore[9][707]<=Wgt_9_707;WeightsStore[9][708]<=Wgt_9_708;WeightsStore[9][709]<=Wgt_9_709;WeightsStore[9][710]<=Wgt_9_710;WeightsStore[9][711]<=Wgt_9_711;WeightsStore[9][712]<=Wgt_9_712;WeightsStore[9][713]<=Wgt_9_713;WeightsStore[9][714]<=Wgt_9_714;WeightsStore[9][715]<=Wgt_9_715;WeightsStore[9][716]<=Wgt_9_716;WeightsStore[9][717]<=Wgt_9_717;WeightsStore[9][718]<=Wgt_9_718;WeightsStore[9][719]<=Wgt_9_719;WeightsStore[9][720]<=Wgt_9_720;WeightsStore[9][721]<=Wgt_9_721;WeightsStore[9][722]<=Wgt_9_722;WeightsStore[9][723]<=Wgt_9_723;WeightsStore[9][724]<=Wgt_9_724;WeightsStore[9][725]<=Wgt_9_725;WeightsStore[9][726]<=Wgt_9_726;WeightsStore[9][727]<=Wgt_9_727;WeightsStore[9][728]<=Wgt_9_728;WeightsStore[9][729]<=Wgt_9_729;WeightsStore[9][730]<=Wgt_9_730;WeightsStore[9][731]<=Wgt_9_731;WeightsStore[9][732]<=Wgt_9_732;WeightsStore[9][733]<=Wgt_9_733;WeightsStore[9][734]<=Wgt_9_734;WeightsStore[9][735]<=Wgt_9_735;WeightsStore[9][736]<=Wgt_9_736;WeightsStore[9][737]<=Wgt_9_737;WeightsStore[9][738]<=Wgt_9_738;WeightsStore[9][739]<=Wgt_9_739;WeightsStore[9][740]<=Wgt_9_740;WeightsStore[9][741]<=Wgt_9_741;WeightsStore[9][742]<=Wgt_9_742;WeightsStore[9][743]<=Wgt_9_743;WeightsStore[9][744]<=Wgt_9_744;WeightsStore[9][745]<=Wgt_9_745;WeightsStore[9][746]<=Wgt_9_746;WeightsStore[9][747]<=Wgt_9_747;WeightsStore[9][748]<=Wgt_9_748;WeightsStore[9][749]<=Wgt_9_749;WeightsStore[9][750]<=Wgt_9_750;WeightsStore[9][751]<=Wgt_9_751;WeightsStore[9][752]<=Wgt_9_752;WeightsStore[9][753]<=Wgt_9_753;WeightsStore[9][754]<=Wgt_9_754;WeightsStore[9][755]<=Wgt_9_755;WeightsStore[9][756]<=Wgt_9_756;WeightsStore[9][757]<=Wgt_9_757;WeightsStore[9][758]<=Wgt_9_758;WeightsStore[9][759]<=Wgt_9_759;WeightsStore[9][760]<=Wgt_9_760;WeightsStore[9][761]<=Wgt_9_761;WeightsStore[9][762]<=Wgt_9_762;WeightsStore[9][763]<=Wgt_9_763;WeightsStore[9][764]<=Wgt_9_764;WeightsStore[9][765]<=Wgt_9_765;WeightsStore[9][766]<=Wgt_9_766;WeightsStore[9][767]<=Wgt_9_767;WeightsStore[9][768]<=Wgt_9_768;WeightsStore[9][769]<=Wgt_9_769;WeightsStore[9][770]<=Wgt_9_770;WeightsStore[9][771]<=Wgt_9_771;WeightsStore[9][772]<=Wgt_9_772;WeightsStore[9][773]<=Wgt_9_773;WeightsStore[9][774]<=Wgt_9_774;WeightsStore[9][775]<=Wgt_9_775;WeightsStore[9][776]<=Wgt_9_776;WeightsStore[9][777]<=Wgt_9_777;WeightsStore[9][778]<=Wgt_9_778;WeightsStore[9][779]<=Wgt_9_779;WeightsStore[9][780]<=Wgt_9_780;WeightsStore[9][781]<=Wgt_9_781;WeightsStore[9][782]<=Wgt_9_782;WeightsStore[9][783]<=Wgt_9_783;WeightsStore[9][784]<=Wgt_9_784;
   end
end
endmodule
