module Image_Classifier(
input clk,
input GlobalReset,
input Input_Valid,
input [18:0] Wgt_0_0,
input [18:0] Wgt_0_1,
input [18:0] Wgt_0_2,
input [18:0] Wgt_0_3,
input [18:0] Wgt_0_4,
input [18:0] Wgt_0_5,
input [18:0] Wgt_0_6,
input [18:0] Wgt_0_7,
input [18:0] Wgt_0_8,
input [18:0] Wgt_0_9,
input [18:0] Wgt_0_10,
input [18:0] Wgt_0_11,
input [18:0] Wgt_0_12,
input [18:0] Wgt_0_13,
input [18:0] Wgt_0_14,
input [18:0] Wgt_0_15,
input [18:0] Wgt_0_16,
input [18:0] Wgt_0_17,
input [18:0] Wgt_0_18,
input [18:0] Wgt_0_19,
input [18:0] Wgt_0_20,
input [18:0] Wgt_0_21,
input [18:0] Wgt_0_22,
input [18:0] Wgt_0_23,
input [18:0] Wgt_0_24,
input [18:0] Wgt_0_25,
input [18:0] Wgt_0_26,
input [18:0] Wgt_0_27,
input [18:0] Wgt_0_28,
input [18:0] Wgt_0_29,
input [18:0] Wgt_0_30,
input [18:0] Wgt_0_31,
input [18:0] Wgt_0_32,
input [18:0] Wgt_0_33,
input [18:0] Wgt_0_34,
input [18:0] Wgt_0_35,
input [18:0] Wgt_0_36,
input [18:0] Wgt_0_37,
input [18:0] Wgt_0_38,
input [18:0] Wgt_0_39,
input [18:0] Wgt_0_40,
input [18:0] Wgt_0_41,
input [18:0] Wgt_0_42,
input [18:0] Wgt_0_43,
input [18:0] Wgt_0_44,
input [18:0] Wgt_0_45,
input [18:0] Wgt_0_46,
input [18:0] Wgt_0_47,
input [18:0] Wgt_0_48,
input [18:0] Wgt_0_49,
input [18:0] Wgt_0_50,
input [18:0] Wgt_0_51,
input [18:0] Wgt_0_52,
input [18:0] Wgt_0_53,
input [18:0] Wgt_0_54,
input [18:0] Wgt_0_55,
input [18:0] Wgt_0_56,
input [18:0] Wgt_0_57,
input [18:0] Wgt_0_58,
input [18:0] Wgt_0_59,
input [18:0] Wgt_0_60,
input [18:0] Wgt_0_61,
input [18:0] Wgt_0_62,
input [18:0] Wgt_0_63,
input [18:0] Wgt_0_64,
input [18:0] Wgt_0_65,
input [18:0] Wgt_0_66,
input [18:0] Wgt_0_67,
input [18:0] Wgt_0_68,
input [18:0] Wgt_0_69,
input [18:0] Wgt_0_70,
input [18:0] Wgt_0_71,
input [18:0] Wgt_0_72,
input [18:0] Wgt_0_73,
input [18:0] Wgt_0_74,
input [18:0] Wgt_0_75,
input [18:0] Wgt_0_76,
input [18:0] Wgt_0_77,
input [18:0] Wgt_0_78,
input [18:0] Wgt_0_79,
input [18:0] Wgt_0_80,
input [18:0] Wgt_0_81,
input [18:0] Wgt_0_82,
input [18:0] Wgt_0_83,
input [18:0] Wgt_0_84,
input [18:0] Wgt_0_85,
input [18:0] Wgt_0_86,
input [18:0] Wgt_0_87,
input [18:0] Wgt_0_88,
input [18:0] Wgt_0_89,
input [18:0] Wgt_0_90,
input [18:0] Wgt_0_91,
input [18:0] Wgt_0_92,
input [18:0] Wgt_0_93,
input [18:0] Wgt_0_94,
input [18:0] Wgt_0_95,
input [18:0] Wgt_0_96,
input [18:0] Wgt_0_97,
input [18:0] Wgt_0_98,
input [18:0] Wgt_0_99,
input [18:0] Wgt_0_100,
input [18:0] Wgt_0_101,
input [18:0] Wgt_0_102,
input [18:0] Wgt_0_103,
input [18:0] Wgt_0_104,
input [18:0] Wgt_0_105,
input [18:0] Wgt_0_106,
input [18:0] Wgt_0_107,
input [18:0] Wgt_0_108,
input [18:0] Wgt_0_109,
input [18:0] Wgt_0_110,
input [18:0] Wgt_0_111,
input [18:0] Wgt_0_112,
input [18:0] Wgt_0_113,
input [18:0] Wgt_0_114,
input [18:0] Wgt_0_115,
input [18:0] Wgt_0_116,
input [18:0] Wgt_0_117,
input [18:0] Wgt_0_118,
input [18:0] Wgt_0_119,
input [18:0] Wgt_0_120,
input [18:0] Wgt_0_121,
input [18:0] Wgt_0_122,
input [18:0] Wgt_0_123,
input [18:0] Wgt_0_124,
input [18:0] Wgt_0_125,
input [18:0] Wgt_0_126,
input [18:0] Wgt_0_127,
input [18:0] Wgt_0_128,
input [18:0] Wgt_0_129,
input [18:0] Wgt_0_130,
input [18:0] Wgt_0_131,
input [18:0] Wgt_0_132,
input [18:0] Wgt_0_133,
input [18:0] Wgt_0_134,
input [18:0] Wgt_0_135,
input [18:0] Wgt_0_136,
input [18:0] Wgt_0_137,
input [18:0] Wgt_0_138,
input [18:0] Wgt_0_139,
input [18:0] Wgt_0_140,
input [18:0] Wgt_0_141,
input [18:0] Wgt_0_142,
input [18:0] Wgt_0_143,
input [18:0] Wgt_0_144,
input [18:0] Wgt_0_145,
input [18:0] Wgt_0_146,
input [18:0] Wgt_0_147,
input [18:0] Wgt_0_148,
input [18:0] Wgt_0_149,
input [18:0] Wgt_0_150,
input [18:0] Wgt_0_151,
input [18:0] Wgt_0_152,
input [18:0] Wgt_0_153,
input [18:0] Wgt_0_154,
input [18:0] Wgt_0_155,
input [18:0] Wgt_0_156,
input [18:0] Wgt_0_157,
input [18:0] Wgt_0_158,
input [18:0] Wgt_0_159,
input [18:0] Wgt_0_160,
input [18:0] Wgt_0_161,
input [18:0] Wgt_0_162,
input [18:0] Wgt_0_163,
input [18:0] Wgt_0_164,
input [18:0] Wgt_0_165,
input [18:0] Wgt_0_166,
input [18:0] Wgt_0_167,
input [18:0] Wgt_0_168,
input [18:0] Wgt_0_169,
input [18:0] Wgt_0_170,
input [18:0] Wgt_0_171,
input [18:0] Wgt_0_172,
input [18:0] Wgt_0_173,
input [18:0] Wgt_0_174,
input [18:0] Wgt_0_175,
input [18:0] Wgt_0_176,
input [18:0] Wgt_0_177,
input [18:0] Wgt_0_178,
input [18:0] Wgt_0_179,
input [18:0] Wgt_0_180,
input [18:0] Wgt_0_181,
input [18:0] Wgt_0_182,
input [18:0] Wgt_0_183,
input [18:0] Wgt_0_184,
input [18:0] Wgt_0_185,
input [18:0] Wgt_0_186,
input [18:0] Wgt_0_187,
input [18:0] Wgt_0_188,
input [18:0] Wgt_0_189,
input [18:0] Wgt_0_190,
input [18:0] Wgt_0_191,
input [18:0] Wgt_0_192,
input [18:0] Wgt_0_193,
input [18:0] Wgt_0_194,
input [18:0] Wgt_0_195,
input [18:0] Wgt_0_196,
input [18:0] Wgt_0_197,
input [18:0] Wgt_0_198,
input [18:0] Wgt_0_199,
input [18:0] Wgt_0_200,
input [18:0] Wgt_0_201,
input [18:0] Wgt_0_202,
input [18:0] Wgt_0_203,
input [18:0] Wgt_0_204,
input [18:0] Wgt_0_205,
input [18:0] Wgt_0_206,
input [18:0] Wgt_0_207,
input [18:0] Wgt_0_208,
input [18:0] Wgt_0_209,
input [18:0] Wgt_0_210,
input [18:0] Wgt_0_211,
input [18:0] Wgt_0_212,
input [18:0] Wgt_0_213,
input [18:0] Wgt_0_214,
input [18:0] Wgt_0_215,
input [18:0] Wgt_0_216,
input [18:0] Wgt_0_217,
input [18:0] Wgt_0_218,
input [18:0] Wgt_0_219,
input [18:0] Wgt_0_220,
input [18:0] Wgt_0_221,
input [18:0] Wgt_0_222,
input [18:0] Wgt_0_223,
input [18:0] Wgt_0_224,
input [18:0] Wgt_0_225,
input [18:0] Wgt_0_226,
input [18:0] Wgt_0_227,
input [18:0] Wgt_0_228,
input [18:0] Wgt_0_229,
input [18:0] Wgt_0_230,
input [18:0] Wgt_0_231,
input [18:0] Wgt_0_232,
input [18:0] Wgt_0_233,
input [18:0] Wgt_0_234,
input [18:0] Wgt_0_235,
input [18:0] Wgt_0_236,
input [18:0] Wgt_0_237,
input [18:0] Wgt_0_238,
input [18:0] Wgt_0_239,
input [18:0] Wgt_0_240,
input [18:0] Wgt_0_241,
input [18:0] Wgt_0_242,
input [18:0] Wgt_0_243,
input [18:0] Wgt_0_244,
input [18:0] Wgt_0_245,
input [18:0] Wgt_0_246,
input [18:0] Wgt_0_247,
input [18:0] Wgt_0_248,
input [18:0] Wgt_0_249,
input [18:0] Wgt_0_250,
input [18:0] Wgt_0_251,
input [18:0] Wgt_0_252,
input [18:0] Wgt_0_253,
input [18:0] Wgt_0_254,
input [18:0] Wgt_0_255,
input [18:0] Wgt_0_256,
input [18:0] Wgt_0_257,
input [18:0] Wgt_0_258,
input [18:0] Wgt_0_259,
input [18:0] Wgt_0_260,
input [18:0] Wgt_0_261,
input [18:0] Wgt_0_262,
input [18:0] Wgt_0_263,
input [18:0] Wgt_0_264,
input [18:0] Wgt_0_265,
input [18:0] Wgt_0_266,
input [18:0] Wgt_0_267,
input [18:0] Wgt_0_268,
input [18:0] Wgt_0_269,
input [18:0] Wgt_0_270,
input [18:0] Wgt_0_271,
input [18:0] Wgt_0_272,
input [18:0] Wgt_0_273,
input [18:0] Wgt_0_274,
input [18:0] Wgt_0_275,
input [18:0] Wgt_0_276,
input [18:0] Wgt_0_277,
input [18:0] Wgt_0_278,
input [18:0] Wgt_0_279,
input [18:0] Wgt_0_280,
input [18:0] Wgt_0_281,
input [18:0] Wgt_0_282,
input [18:0] Wgt_0_283,
input [18:0] Wgt_0_284,
input [18:0] Wgt_0_285,
input [18:0] Wgt_0_286,
input [18:0] Wgt_0_287,
input [18:0] Wgt_0_288,
input [18:0] Wgt_0_289,
input [18:0] Wgt_0_290,
input [18:0] Wgt_0_291,
input [18:0] Wgt_0_292,
input [18:0] Wgt_0_293,
input [18:0] Wgt_0_294,
input [18:0] Wgt_0_295,
input [18:0] Wgt_0_296,
input [18:0] Wgt_0_297,
input [18:0] Wgt_0_298,
input [18:0] Wgt_0_299,
input [18:0] Wgt_0_300,
input [18:0] Wgt_0_301,
input [18:0] Wgt_0_302,
input [18:0] Wgt_0_303,
input [18:0] Wgt_0_304,
input [18:0] Wgt_0_305,
input [18:0] Wgt_0_306,
input [18:0] Wgt_0_307,
input [18:0] Wgt_0_308,
input [18:0] Wgt_0_309,
input [18:0] Wgt_0_310,
input [18:0] Wgt_0_311,
input [18:0] Wgt_0_312,
input [18:0] Wgt_0_313,
input [18:0] Wgt_0_314,
input [18:0] Wgt_0_315,
input [18:0] Wgt_0_316,
input [18:0] Wgt_0_317,
input [18:0] Wgt_0_318,
input [18:0] Wgt_0_319,
input [18:0] Wgt_0_320,
input [18:0] Wgt_0_321,
input [18:0] Wgt_0_322,
input [18:0] Wgt_0_323,
input [18:0] Wgt_0_324,
input [18:0] Wgt_0_325,
input [18:0] Wgt_0_326,
input [18:0] Wgt_0_327,
input [18:0] Wgt_0_328,
input [18:0] Wgt_0_329,
input [18:0] Wgt_0_330,
input [18:0] Wgt_0_331,
input [18:0] Wgt_0_332,
input [18:0] Wgt_0_333,
input [18:0] Wgt_0_334,
input [18:0] Wgt_0_335,
input [18:0] Wgt_0_336,
input [18:0] Wgt_0_337,
input [18:0] Wgt_0_338,
input [18:0] Wgt_0_339,
input [18:0] Wgt_0_340,
input [18:0] Wgt_0_341,
input [18:0] Wgt_0_342,
input [18:0] Wgt_0_343,
input [18:0] Wgt_0_344,
input [18:0] Wgt_0_345,
input [18:0] Wgt_0_346,
input [18:0] Wgt_0_347,
input [18:0] Wgt_0_348,
input [18:0] Wgt_0_349,
input [18:0] Wgt_0_350,
input [18:0] Wgt_0_351,
input [18:0] Wgt_0_352,
input [18:0] Wgt_0_353,
input [18:0] Wgt_0_354,
input [18:0] Wgt_0_355,
input [18:0] Wgt_0_356,
input [18:0] Wgt_0_357,
input [18:0] Wgt_0_358,
input [18:0] Wgt_0_359,
input [18:0] Wgt_0_360,
input [18:0] Wgt_0_361,
input [18:0] Wgt_0_362,
input [18:0] Wgt_0_363,
input [18:0] Wgt_0_364,
input [18:0] Wgt_0_365,
input [18:0] Wgt_0_366,
input [18:0] Wgt_0_367,
input [18:0] Wgt_0_368,
input [18:0] Wgt_0_369,
input [18:0] Wgt_0_370,
input [18:0] Wgt_0_371,
input [18:0] Wgt_0_372,
input [18:0] Wgt_0_373,
input [18:0] Wgt_0_374,
input [18:0] Wgt_0_375,
input [18:0] Wgt_0_376,
input [18:0] Wgt_0_377,
input [18:0] Wgt_0_378,
input [18:0] Wgt_0_379,
input [18:0] Wgt_0_380,
input [18:0] Wgt_0_381,
input [18:0] Wgt_0_382,
input [18:0] Wgt_0_383,
input [18:0] Wgt_0_384,
input [18:0] Wgt_0_385,
input [18:0] Wgt_0_386,
input [18:0] Wgt_0_387,
input [18:0] Wgt_0_388,
input [18:0] Wgt_0_389,
input [18:0] Wgt_0_390,
input [18:0] Wgt_0_391,
input [18:0] Wgt_0_392,
input [18:0] Wgt_0_393,
input [18:0] Wgt_0_394,
input [18:0] Wgt_0_395,
input [18:0] Wgt_0_396,
input [18:0] Wgt_0_397,
input [18:0] Wgt_0_398,
input [18:0] Wgt_0_399,
input [18:0] Wgt_0_400,
input [18:0] Wgt_0_401,
input [18:0] Wgt_0_402,
input [18:0] Wgt_0_403,
input [18:0] Wgt_0_404,
input [18:0] Wgt_0_405,
input [18:0] Wgt_0_406,
input [18:0] Wgt_0_407,
input [18:0] Wgt_0_408,
input [18:0] Wgt_0_409,
input [18:0] Wgt_0_410,
input [18:0] Wgt_0_411,
input [18:0] Wgt_0_412,
input [18:0] Wgt_0_413,
input [18:0] Wgt_0_414,
input [18:0] Wgt_0_415,
input [18:0] Wgt_0_416,
input [18:0] Wgt_0_417,
input [18:0] Wgt_0_418,
input [18:0] Wgt_0_419,
input [18:0] Wgt_0_420,
input [18:0] Wgt_0_421,
input [18:0] Wgt_0_422,
input [18:0] Wgt_0_423,
input [18:0] Wgt_0_424,
input [18:0] Wgt_0_425,
input [18:0] Wgt_0_426,
input [18:0] Wgt_0_427,
input [18:0] Wgt_0_428,
input [18:0] Wgt_0_429,
input [18:0] Wgt_0_430,
input [18:0] Wgt_0_431,
input [18:0] Wgt_0_432,
input [18:0] Wgt_0_433,
input [18:0] Wgt_0_434,
input [18:0] Wgt_0_435,
input [18:0] Wgt_0_436,
input [18:0] Wgt_0_437,
input [18:0] Wgt_0_438,
input [18:0] Wgt_0_439,
input [18:0] Wgt_0_440,
input [18:0] Wgt_0_441,
input [18:0] Wgt_0_442,
input [18:0] Wgt_0_443,
input [18:0] Wgt_0_444,
input [18:0] Wgt_0_445,
input [18:0] Wgt_0_446,
input [18:0] Wgt_0_447,
input [18:0] Wgt_0_448,
input [18:0] Wgt_0_449,
input [18:0] Wgt_0_450,
input [18:0] Wgt_0_451,
input [18:0] Wgt_0_452,
input [18:0] Wgt_0_453,
input [18:0] Wgt_0_454,
input [18:0] Wgt_0_455,
input [18:0] Wgt_0_456,
input [18:0] Wgt_0_457,
input [18:0] Wgt_0_458,
input [18:0] Wgt_0_459,
input [18:0] Wgt_0_460,
input [18:0] Wgt_0_461,
input [18:0] Wgt_0_462,
input [18:0] Wgt_0_463,
input [18:0] Wgt_0_464,
input [18:0] Wgt_0_465,
input [18:0] Wgt_0_466,
input [18:0] Wgt_0_467,
input [18:0] Wgt_0_468,
input [18:0] Wgt_0_469,
input [18:0] Wgt_0_470,
input [18:0] Wgt_0_471,
input [18:0] Wgt_0_472,
input [18:0] Wgt_0_473,
input [18:0] Wgt_0_474,
input [18:0] Wgt_0_475,
input [18:0] Wgt_0_476,
input [18:0] Wgt_0_477,
input [18:0] Wgt_0_478,
input [18:0] Wgt_0_479,
input [18:0] Wgt_0_480,
input [18:0] Wgt_0_481,
input [18:0] Wgt_0_482,
input [18:0] Wgt_0_483,
input [18:0] Wgt_0_484,
input [18:0] Wgt_0_485,
input [18:0] Wgt_0_486,
input [18:0] Wgt_0_487,
input [18:0] Wgt_0_488,
input [18:0] Wgt_0_489,
input [18:0] Wgt_0_490,
input [18:0] Wgt_0_491,
input [18:0] Wgt_0_492,
input [18:0] Wgt_0_493,
input [18:0] Wgt_0_494,
input [18:0] Wgt_0_495,
input [18:0] Wgt_0_496,
input [18:0] Wgt_0_497,
input [18:0] Wgt_0_498,
input [18:0] Wgt_0_499,
input [18:0] Wgt_0_500,
input [18:0] Wgt_0_501,
input [18:0] Wgt_0_502,
input [18:0] Wgt_0_503,
input [18:0] Wgt_0_504,
input [18:0] Wgt_0_505,
input [18:0] Wgt_0_506,
input [18:0] Wgt_0_507,
input [18:0] Wgt_0_508,
input [18:0] Wgt_0_509,
input [18:0] Wgt_0_510,
input [18:0] Wgt_0_511,
input [18:0] Wgt_0_512,
input [18:0] Wgt_0_513,
input [18:0] Wgt_0_514,
input [18:0] Wgt_0_515,
input [18:0] Wgt_0_516,
input [18:0] Wgt_0_517,
input [18:0] Wgt_0_518,
input [18:0] Wgt_0_519,
input [18:0] Wgt_0_520,
input [18:0] Wgt_0_521,
input [18:0] Wgt_0_522,
input [18:0] Wgt_0_523,
input [18:0] Wgt_0_524,
input [18:0] Wgt_0_525,
input [18:0] Wgt_0_526,
input [18:0] Wgt_0_527,
input [18:0] Wgt_0_528,
input [18:0] Wgt_0_529,
input [18:0] Wgt_0_530,
input [18:0] Wgt_0_531,
input [18:0] Wgt_0_532,
input [18:0] Wgt_0_533,
input [18:0] Wgt_0_534,
input [18:0] Wgt_0_535,
input [18:0] Wgt_0_536,
input [18:0] Wgt_0_537,
input [18:0] Wgt_0_538,
input [18:0] Wgt_0_539,
input [18:0] Wgt_0_540,
input [18:0] Wgt_0_541,
input [18:0] Wgt_0_542,
input [18:0] Wgt_0_543,
input [18:0] Wgt_0_544,
input [18:0] Wgt_0_545,
input [18:0] Wgt_0_546,
input [18:0] Wgt_0_547,
input [18:0] Wgt_0_548,
input [18:0] Wgt_0_549,
input [18:0] Wgt_0_550,
input [18:0] Wgt_0_551,
input [18:0] Wgt_0_552,
input [18:0] Wgt_0_553,
input [18:0] Wgt_0_554,
input [18:0] Wgt_0_555,
input [18:0] Wgt_0_556,
input [18:0] Wgt_0_557,
input [18:0] Wgt_0_558,
input [18:0] Wgt_0_559,
input [18:0] Wgt_0_560,
input [18:0] Wgt_0_561,
input [18:0] Wgt_0_562,
input [18:0] Wgt_0_563,
input [18:0] Wgt_0_564,
input [18:0] Wgt_0_565,
input [18:0] Wgt_0_566,
input [18:0] Wgt_0_567,
input [18:0] Wgt_0_568,
input [18:0] Wgt_0_569,
input [18:0] Wgt_0_570,
input [18:0] Wgt_0_571,
input [18:0] Wgt_0_572,
input [18:0] Wgt_0_573,
input [18:0] Wgt_0_574,
input [18:0] Wgt_0_575,
input [18:0] Wgt_0_576,
input [18:0] Wgt_0_577,
input [18:0] Wgt_0_578,
input [18:0] Wgt_0_579,
input [18:0] Wgt_0_580,
input [18:0] Wgt_0_581,
input [18:0] Wgt_0_582,
input [18:0] Wgt_0_583,
input [18:0] Wgt_0_584,
input [18:0] Wgt_0_585,
input [18:0] Wgt_0_586,
input [18:0] Wgt_0_587,
input [18:0] Wgt_0_588,
input [18:0] Wgt_0_589,
input [18:0] Wgt_0_590,
input [18:0] Wgt_0_591,
input [18:0] Wgt_0_592,
input [18:0] Wgt_0_593,
input [18:0] Wgt_0_594,
input [18:0] Wgt_0_595,
input [18:0] Wgt_0_596,
input [18:0] Wgt_0_597,
input [18:0] Wgt_0_598,
input [18:0] Wgt_0_599,
input [18:0] Wgt_0_600,
input [18:0] Wgt_0_601,
input [18:0] Wgt_0_602,
input [18:0] Wgt_0_603,
input [18:0] Wgt_0_604,
input [18:0] Wgt_0_605,
input [18:0] Wgt_0_606,
input [18:0] Wgt_0_607,
input [18:0] Wgt_0_608,
input [18:0] Wgt_0_609,
input [18:0] Wgt_0_610,
input [18:0] Wgt_0_611,
input [18:0] Wgt_0_612,
input [18:0] Wgt_0_613,
input [18:0] Wgt_0_614,
input [18:0] Wgt_0_615,
input [18:0] Wgt_0_616,
input [18:0] Wgt_0_617,
input [18:0] Wgt_0_618,
input [18:0] Wgt_0_619,
input [18:0] Wgt_0_620,
input [18:0] Wgt_0_621,
input [18:0] Wgt_0_622,
input [18:0] Wgt_0_623,
input [18:0] Wgt_0_624,
input [18:0] Wgt_0_625,
input [18:0] Wgt_0_626,
input [18:0] Wgt_0_627,
input [18:0] Wgt_0_628,
input [18:0] Wgt_0_629,
input [18:0] Wgt_0_630,
input [18:0] Wgt_0_631,
input [18:0] Wgt_0_632,
input [18:0] Wgt_0_633,
input [18:0] Wgt_0_634,
input [18:0] Wgt_0_635,
input [18:0] Wgt_0_636,
input [18:0] Wgt_0_637,
input [18:0] Wgt_0_638,
input [18:0] Wgt_0_639,
input [18:0] Wgt_0_640,
input [18:0] Wgt_0_641,
input [18:0] Wgt_0_642,
input [18:0] Wgt_0_643,
input [18:0] Wgt_0_644,
input [18:0] Wgt_0_645,
input [18:0] Wgt_0_646,
input [18:0] Wgt_0_647,
input [18:0] Wgt_0_648,
input [18:0] Wgt_0_649,
input [18:0] Wgt_0_650,
input [18:0] Wgt_0_651,
input [18:0] Wgt_0_652,
input [18:0] Wgt_0_653,
input [18:0] Wgt_0_654,
input [18:0] Wgt_0_655,
input [18:0] Wgt_0_656,
input [18:0] Wgt_0_657,
input [18:0] Wgt_0_658,
input [18:0] Wgt_0_659,
input [18:0] Wgt_0_660,
input [18:0] Wgt_0_661,
input [18:0] Wgt_0_662,
input [18:0] Wgt_0_663,
input [18:0] Wgt_0_664,
input [18:0] Wgt_0_665,
input [18:0] Wgt_0_666,
input [18:0] Wgt_0_667,
input [18:0] Wgt_0_668,
input [18:0] Wgt_0_669,
input [18:0] Wgt_0_670,
input [18:0] Wgt_0_671,
input [18:0] Wgt_0_672,
input [18:0] Wgt_0_673,
input [18:0] Wgt_0_674,
input [18:0] Wgt_0_675,
input [18:0] Wgt_0_676,
input [18:0] Wgt_0_677,
input [18:0] Wgt_0_678,
input [18:0] Wgt_0_679,
input [18:0] Wgt_0_680,
input [18:0] Wgt_0_681,
input [18:0] Wgt_0_682,
input [18:0] Wgt_0_683,
input [18:0] Wgt_0_684,
input [18:0] Wgt_0_685,
input [18:0] Wgt_0_686,
input [18:0] Wgt_0_687,
input [18:0] Wgt_0_688,
input [18:0] Wgt_0_689,
input [18:0] Wgt_0_690,
input [18:0] Wgt_0_691,
input [18:0] Wgt_0_692,
input [18:0] Wgt_0_693,
input [18:0] Wgt_0_694,
input [18:0] Wgt_0_695,
input [18:0] Wgt_0_696,
input [18:0] Wgt_0_697,
input [18:0] Wgt_0_698,
input [18:0] Wgt_0_699,
input [18:0] Wgt_0_700,
input [18:0] Wgt_0_701,
input [18:0] Wgt_0_702,
input [18:0] Wgt_0_703,
input [18:0] Wgt_0_704,
input [18:0] Wgt_0_705,
input [18:0] Wgt_0_706,
input [18:0] Wgt_0_707,
input [18:0] Wgt_0_708,
input [18:0] Wgt_0_709,
input [18:0] Wgt_0_710,
input [18:0] Wgt_0_711,
input [18:0] Wgt_0_712,
input [18:0] Wgt_0_713,
input [18:0] Wgt_0_714,
input [18:0] Wgt_0_715,
input [18:0] Wgt_0_716,
input [18:0] Wgt_0_717,
input [18:0] Wgt_0_718,
input [18:0] Wgt_0_719,
input [18:0] Wgt_0_720,
input [18:0] Wgt_0_721,
input [18:0] Wgt_0_722,
input [18:0] Wgt_0_723,
input [18:0] Wgt_0_724,
input [18:0] Wgt_0_725,
input [18:0] Wgt_0_726,
input [18:0] Wgt_0_727,
input [18:0] Wgt_0_728,
input [18:0] Wgt_0_729,
input [18:0] Wgt_0_730,
input [18:0] Wgt_0_731,
input [18:0] Wgt_0_732,
input [18:0] Wgt_0_733,
input [18:0] Wgt_0_734,
input [18:0] Wgt_0_735,
input [18:0] Wgt_0_736,
input [18:0] Wgt_0_737,
input [18:0] Wgt_0_738,
input [18:0] Wgt_0_739,
input [18:0] Wgt_0_740,
input [18:0] Wgt_0_741,
input [18:0] Wgt_0_742,
input [18:0] Wgt_0_743,
input [18:0] Wgt_0_744,
input [18:0] Wgt_0_745,
input [18:0] Wgt_0_746,
input [18:0] Wgt_0_747,
input [18:0] Wgt_0_748,
input [18:0] Wgt_0_749,
input [18:0] Wgt_0_750,
input [18:0] Wgt_0_751,
input [18:0] Wgt_0_752,
input [18:0] Wgt_0_753,
input [18:0] Wgt_0_754,
input [18:0] Wgt_0_755,
input [18:0] Wgt_0_756,
input [18:0] Wgt_0_757,
input [18:0] Wgt_0_758,
input [18:0] Wgt_0_759,
input [18:0] Wgt_0_760,
input [18:0] Wgt_0_761,
input [18:0] Wgt_0_762,
input [18:0] Wgt_0_763,
input [18:0] Wgt_0_764,
input [18:0] Wgt_0_765,
input [18:0] Wgt_0_766,
input [18:0] Wgt_0_767,
input [18:0] Wgt_0_768,
input [18:0] Wgt_0_769,
input [18:0] Wgt_0_770,
input [18:0] Wgt_0_771,
input [18:0] Wgt_0_772,
input [18:0] Wgt_0_773,
input [18:0] Wgt_0_774,
input [18:0] Wgt_0_775,
input [18:0] Wgt_0_776,
input [18:0] Wgt_0_777,
input [18:0] Wgt_0_778,
input [18:0] Wgt_0_779,
input [18:0] Wgt_0_780,
input [18:0] Wgt_0_781,
input [18:0] Wgt_0_782,
input [18:0] Wgt_0_783,
input [18:0] Wgt_0_784,
input [18:0] Wgt_1_0,
input [18:0] Wgt_1_1,
input [18:0] Wgt_1_2,
input [18:0] Wgt_1_3,
input [18:0] Wgt_1_4,
input [18:0] Wgt_1_5,
input [18:0] Wgt_1_6,
input [18:0] Wgt_1_7,
input [18:0] Wgt_1_8,
input [18:0] Wgt_1_9,
input [18:0] Wgt_1_10,
input [18:0] Wgt_1_11,
input [18:0] Wgt_1_12,
input [18:0] Wgt_1_13,
input [18:0] Wgt_1_14,
input [18:0] Wgt_1_15,
input [18:0] Wgt_1_16,
input [18:0] Wgt_1_17,
input [18:0] Wgt_1_18,
input [18:0] Wgt_1_19,
input [18:0] Wgt_1_20,
input [18:0] Wgt_1_21,
input [18:0] Wgt_1_22,
input [18:0] Wgt_1_23,
input [18:0] Wgt_1_24,
input [18:0] Wgt_1_25,
input [18:0] Wgt_1_26,
input [18:0] Wgt_1_27,
input [18:0] Wgt_1_28,
input [18:0] Wgt_1_29,
input [18:0] Wgt_1_30,
input [18:0] Wgt_1_31,
input [18:0] Wgt_1_32,
input [18:0] Wgt_1_33,
input [18:0] Wgt_1_34,
input [18:0] Wgt_1_35,
input [18:0] Wgt_1_36,
input [18:0] Wgt_1_37,
input [18:0] Wgt_1_38,
input [18:0] Wgt_1_39,
input [18:0] Wgt_1_40,
input [18:0] Wgt_1_41,
input [18:0] Wgt_1_42,
input [18:0] Wgt_1_43,
input [18:0] Wgt_1_44,
input [18:0] Wgt_1_45,
input [18:0] Wgt_1_46,
input [18:0] Wgt_1_47,
input [18:0] Wgt_1_48,
input [18:0] Wgt_1_49,
input [18:0] Wgt_1_50,
input [18:0] Wgt_1_51,
input [18:0] Wgt_1_52,
input [18:0] Wgt_1_53,
input [18:0] Wgt_1_54,
input [18:0] Wgt_1_55,
input [18:0] Wgt_1_56,
input [18:0] Wgt_1_57,
input [18:0] Wgt_1_58,
input [18:0] Wgt_1_59,
input [18:0] Wgt_1_60,
input [18:0] Wgt_1_61,
input [18:0] Wgt_1_62,
input [18:0] Wgt_1_63,
input [18:0] Wgt_1_64,
input [18:0] Wgt_1_65,
input [18:0] Wgt_1_66,
input [18:0] Wgt_1_67,
input [18:0] Wgt_1_68,
input [18:0] Wgt_1_69,
input [18:0] Wgt_1_70,
input [18:0] Wgt_1_71,
input [18:0] Wgt_1_72,
input [18:0] Wgt_1_73,
input [18:0] Wgt_1_74,
input [18:0] Wgt_1_75,
input [18:0] Wgt_1_76,
input [18:0] Wgt_1_77,
input [18:0] Wgt_1_78,
input [18:0] Wgt_1_79,
input [18:0] Wgt_1_80,
input [18:0] Wgt_1_81,
input [18:0] Wgt_1_82,
input [18:0] Wgt_1_83,
input [18:0] Wgt_1_84,
input [18:0] Wgt_1_85,
input [18:0] Wgt_1_86,
input [18:0] Wgt_1_87,
input [18:0] Wgt_1_88,
input [18:0] Wgt_1_89,
input [18:0] Wgt_1_90,
input [18:0] Wgt_1_91,
input [18:0] Wgt_1_92,
input [18:0] Wgt_1_93,
input [18:0] Wgt_1_94,
input [18:0] Wgt_1_95,
input [18:0] Wgt_1_96,
input [18:0] Wgt_1_97,
input [18:0] Wgt_1_98,
input [18:0] Wgt_1_99,
input [18:0] Wgt_1_100,
input [18:0] Wgt_1_101,
input [18:0] Wgt_1_102,
input [18:0] Wgt_1_103,
input [18:0] Wgt_1_104,
input [18:0] Wgt_1_105,
input [18:0] Wgt_1_106,
input [18:0] Wgt_1_107,
input [18:0] Wgt_1_108,
input [18:0] Wgt_1_109,
input [18:0] Wgt_1_110,
input [18:0] Wgt_1_111,
input [18:0] Wgt_1_112,
input [18:0] Wgt_1_113,
input [18:0] Wgt_1_114,
input [18:0] Wgt_1_115,
input [18:0] Wgt_1_116,
input [18:0] Wgt_1_117,
input [18:0] Wgt_1_118,
input [18:0] Wgt_1_119,
input [18:0] Wgt_1_120,
input [18:0] Wgt_1_121,
input [18:0] Wgt_1_122,
input [18:0] Wgt_1_123,
input [18:0] Wgt_1_124,
input [18:0] Wgt_1_125,
input [18:0] Wgt_1_126,
input [18:0] Wgt_1_127,
input [18:0] Wgt_1_128,
input [18:0] Wgt_1_129,
input [18:0] Wgt_1_130,
input [18:0] Wgt_1_131,
input [18:0] Wgt_1_132,
input [18:0] Wgt_1_133,
input [18:0] Wgt_1_134,
input [18:0] Wgt_1_135,
input [18:0] Wgt_1_136,
input [18:0] Wgt_1_137,
input [18:0] Wgt_1_138,
input [18:0] Wgt_1_139,
input [18:0] Wgt_1_140,
input [18:0] Wgt_1_141,
input [18:0] Wgt_1_142,
input [18:0] Wgt_1_143,
input [18:0] Wgt_1_144,
input [18:0] Wgt_1_145,
input [18:0] Wgt_1_146,
input [18:0] Wgt_1_147,
input [18:0] Wgt_1_148,
input [18:0] Wgt_1_149,
input [18:0] Wgt_1_150,
input [18:0] Wgt_1_151,
input [18:0] Wgt_1_152,
input [18:0] Wgt_1_153,
input [18:0] Wgt_1_154,
input [18:0] Wgt_1_155,
input [18:0] Wgt_1_156,
input [18:0] Wgt_1_157,
input [18:0] Wgt_1_158,
input [18:0] Wgt_1_159,
input [18:0] Wgt_1_160,
input [18:0] Wgt_1_161,
input [18:0] Wgt_1_162,
input [18:0] Wgt_1_163,
input [18:0] Wgt_1_164,
input [18:0] Wgt_1_165,
input [18:0] Wgt_1_166,
input [18:0] Wgt_1_167,
input [18:0] Wgt_1_168,
input [18:0] Wgt_1_169,
input [18:0] Wgt_1_170,
input [18:0] Wgt_1_171,
input [18:0] Wgt_1_172,
input [18:0] Wgt_1_173,
input [18:0] Wgt_1_174,
input [18:0] Wgt_1_175,
input [18:0] Wgt_1_176,
input [18:0] Wgt_1_177,
input [18:0] Wgt_1_178,
input [18:0] Wgt_1_179,
input [18:0] Wgt_1_180,
input [18:0] Wgt_1_181,
input [18:0] Wgt_1_182,
input [18:0] Wgt_1_183,
input [18:0] Wgt_1_184,
input [18:0] Wgt_1_185,
input [18:0] Wgt_1_186,
input [18:0] Wgt_1_187,
input [18:0] Wgt_1_188,
input [18:0] Wgt_1_189,
input [18:0] Wgt_1_190,
input [18:0] Wgt_1_191,
input [18:0] Wgt_1_192,
input [18:0] Wgt_1_193,
input [18:0] Wgt_1_194,
input [18:0] Wgt_1_195,
input [18:0] Wgt_1_196,
input [18:0] Wgt_1_197,
input [18:0] Wgt_1_198,
input [18:0] Wgt_1_199,
input [18:0] Wgt_1_200,
input [18:0] Wgt_1_201,
input [18:0] Wgt_1_202,
input [18:0] Wgt_1_203,
input [18:0] Wgt_1_204,
input [18:0] Wgt_1_205,
input [18:0] Wgt_1_206,
input [18:0] Wgt_1_207,
input [18:0] Wgt_1_208,
input [18:0] Wgt_1_209,
input [18:0] Wgt_1_210,
input [18:0] Wgt_1_211,
input [18:0] Wgt_1_212,
input [18:0] Wgt_1_213,
input [18:0] Wgt_1_214,
input [18:0] Wgt_1_215,
input [18:0] Wgt_1_216,
input [18:0] Wgt_1_217,
input [18:0] Wgt_1_218,
input [18:0] Wgt_1_219,
input [18:0] Wgt_1_220,
input [18:0] Wgt_1_221,
input [18:0] Wgt_1_222,
input [18:0] Wgt_1_223,
input [18:0] Wgt_1_224,
input [18:0] Wgt_1_225,
input [18:0] Wgt_1_226,
input [18:0] Wgt_1_227,
input [18:0] Wgt_1_228,
input [18:0] Wgt_1_229,
input [18:0] Wgt_1_230,
input [18:0] Wgt_1_231,
input [18:0] Wgt_1_232,
input [18:0] Wgt_1_233,
input [18:0] Wgt_1_234,
input [18:0] Wgt_1_235,
input [18:0] Wgt_1_236,
input [18:0] Wgt_1_237,
input [18:0] Wgt_1_238,
input [18:0] Wgt_1_239,
input [18:0] Wgt_1_240,
input [18:0] Wgt_1_241,
input [18:0] Wgt_1_242,
input [18:0] Wgt_1_243,
input [18:0] Wgt_1_244,
input [18:0] Wgt_1_245,
input [18:0] Wgt_1_246,
input [18:0] Wgt_1_247,
input [18:0] Wgt_1_248,
input [18:0] Wgt_1_249,
input [18:0] Wgt_1_250,
input [18:0] Wgt_1_251,
input [18:0] Wgt_1_252,
input [18:0] Wgt_1_253,
input [18:0] Wgt_1_254,
input [18:0] Wgt_1_255,
input [18:0] Wgt_1_256,
input [18:0] Wgt_1_257,
input [18:0] Wgt_1_258,
input [18:0] Wgt_1_259,
input [18:0] Wgt_1_260,
input [18:0] Wgt_1_261,
input [18:0] Wgt_1_262,
input [18:0] Wgt_1_263,
input [18:0] Wgt_1_264,
input [18:0] Wgt_1_265,
input [18:0] Wgt_1_266,
input [18:0] Wgt_1_267,
input [18:0] Wgt_1_268,
input [18:0] Wgt_1_269,
input [18:0] Wgt_1_270,
input [18:0] Wgt_1_271,
input [18:0] Wgt_1_272,
input [18:0] Wgt_1_273,
input [18:0] Wgt_1_274,
input [18:0] Wgt_1_275,
input [18:0] Wgt_1_276,
input [18:0] Wgt_1_277,
input [18:0] Wgt_1_278,
input [18:0] Wgt_1_279,
input [18:0] Wgt_1_280,
input [18:0] Wgt_1_281,
input [18:0] Wgt_1_282,
input [18:0] Wgt_1_283,
input [18:0] Wgt_1_284,
input [18:0] Wgt_1_285,
input [18:0] Wgt_1_286,
input [18:0] Wgt_1_287,
input [18:0] Wgt_1_288,
input [18:0] Wgt_1_289,
input [18:0] Wgt_1_290,
input [18:0] Wgt_1_291,
input [18:0] Wgt_1_292,
input [18:0] Wgt_1_293,
input [18:0] Wgt_1_294,
input [18:0] Wgt_1_295,
input [18:0] Wgt_1_296,
input [18:0] Wgt_1_297,
input [18:0] Wgt_1_298,
input [18:0] Wgt_1_299,
input [18:0] Wgt_1_300,
input [18:0] Wgt_1_301,
input [18:0] Wgt_1_302,
input [18:0] Wgt_1_303,
input [18:0] Wgt_1_304,
input [18:0] Wgt_1_305,
input [18:0] Wgt_1_306,
input [18:0] Wgt_1_307,
input [18:0] Wgt_1_308,
input [18:0] Wgt_1_309,
input [18:0] Wgt_1_310,
input [18:0] Wgt_1_311,
input [18:0] Wgt_1_312,
input [18:0] Wgt_1_313,
input [18:0] Wgt_1_314,
input [18:0] Wgt_1_315,
input [18:0] Wgt_1_316,
input [18:0] Wgt_1_317,
input [18:0] Wgt_1_318,
input [18:0] Wgt_1_319,
input [18:0] Wgt_1_320,
input [18:0] Wgt_1_321,
input [18:0] Wgt_1_322,
input [18:0] Wgt_1_323,
input [18:0] Wgt_1_324,
input [18:0] Wgt_1_325,
input [18:0] Wgt_1_326,
input [18:0] Wgt_1_327,
input [18:0] Wgt_1_328,
input [18:0] Wgt_1_329,
input [18:0] Wgt_1_330,
input [18:0] Wgt_1_331,
input [18:0] Wgt_1_332,
input [18:0] Wgt_1_333,
input [18:0] Wgt_1_334,
input [18:0] Wgt_1_335,
input [18:0] Wgt_1_336,
input [18:0] Wgt_1_337,
input [18:0] Wgt_1_338,
input [18:0] Wgt_1_339,
input [18:0] Wgt_1_340,
input [18:0] Wgt_1_341,
input [18:0] Wgt_1_342,
input [18:0] Wgt_1_343,
input [18:0] Wgt_1_344,
input [18:0] Wgt_1_345,
input [18:0] Wgt_1_346,
input [18:0] Wgt_1_347,
input [18:0] Wgt_1_348,
input [18:0] Wgt_1_349,
input [18:0] Wgt_1_350,
input [18:0] Wgt_1_351,
input [18:0] Wgt_1_352,
input [18:0] Wgt_1_353,
input [18:0] Wgt_1_354,
input [18:0] Wgt_1_355,
input [18:0] Wgt_1_356,
input [18:0] Wgt_1_357,
input [18:0] Wgt_1_358,
input [18:0] Wgt_1_359,
input [18:0] Wgt_1_360,
input [18:0] Wgt_1_361,
input [18:0] Wgt_1_362,
input [18:0] Wgt_1_363,
input [18:0] Wgt_1_364,
input [18:0] Wgt_1_365,
input [18:0] Wgt_1_366,
input [18:0] Wgt_1_367,
input [18:0] Wgt_1_368,
input [18:0] Wgt_1_369,
input [18:0] Wgt_1_370,
input [18:0] Wgt_1_371,
input [18:0] Wgt_1_372,
input [18:0] Wgt_1_373,
input [18:0] Wgt_1_374,
input [18:0] Wgt_1_375,
input [18:0] Wgt_1_376,
input [18:0] Wgt_1_377,
input [18:0] Wgt_1_378,
input [18:0] Wgt_1_379,
input [18:0] Wgt_1_380,
input [18:0] Wgt_1_381,
input [18:0] Wgt_1_382,
input [18:0] Wgt_1_383,
input [18:0] Wgt_1_384,
input [18:0] Wgt_1_385,
input [18:0] Wgt_1_386,
input [18:0] Wgt_1_387,
input [18:0] Wgt_1_388,
input [18:0] Wgt_1_389,
input [18:0] Wgt_1_390,
input [18:0] Wgt_1_391,
input [18:0] Wgt_1_392,
input [18:0] Wgt_1_393,
input [18:0] Wgt_1_394,
input [18:0] Wgt_1_395,
input [18:0] Wgt_1_396,
input [18:0] Wgt_1_397,
input [18:0] Wgt_1_398,
input [18:0] Wgt_1_399,
input [18:0] Wgt_1_400,
input [18:0] Wgt_1_401,
input [18:0] Wgt_1_402,
input [18:0] Wgt_1_403,
input [18:0] Wgt_1_404,
input [18:0] Wgt_1_405,
input [18:0] Wgt_1_406,
input [18:0] Wgt_1_407,
input [18:0] Wgt_1_408,
input [18:0] Wgt_1_409,
input [18:0] Wgt_1_410,
input [18:0] Wgt_1_411,
input [18:0] Wgt_1_412,
input [18:0] Wgt_1_413,
input [18:0] Wgt_1_414,
input [18:0] Wgt_1_415,
input [18:0] Wgt_1_416,
input [18:0] Wgt_1_417,
input [18:0] Wgt_1_418,
input [18:0] Wgt_1_419,
input [18:0] Wgt_1_420,
input [18:0] Wgt_1_421,
input [18:0] Wgt_1_422,
input [18:0] Wgt_1_423,
input [18:0] Wgt_1_424,
input [18:0] Wgt_1_425,
input [18:0] Wgt_1_426,
input [18:0] Wgt_1_427,
input [18:0] Wgt_1_428,
input [18:0] Wgt_1_429,
input [18:0] Wgt_1_430,
input [18:0] Wgt_1_431,
input [18:0] Wgt_1_432,
input [18:0] Wgt_1_433,
input [18:0] Wgt_1_434,
input [18:0] Wgt_1_435,
input [18:0] Wgt_1_436,
input [18:0] Wgt_1_437,
input [18:0] Wgt_1_438,
input [18:0] Wgt_1_439,
input [18:0] Wgt_1_440,
input [18:0] Wgt_1_441,
input [18:0] Wgt_1_442,
input [18:0] Wgt_1_443,
input [18:0] Wgt_1_444,
input [18:0] Wgt_1_445,
input [18:0] Wgt_1_446,
input [18:0] Wgt_1_447,
input [18:0] Wgt_1_448,
input [18:0] Wgt_1_449,
input [18:0] Wgt_1_450,
input [18:0] Wgt_1_451,
input [18:0] Wgt_1_452,
input [18:0] Wgt_1_453,
input [18:0] Wgt_1_454,
input [18:0] Wgt_1_455,
input [18:0] Wgt_1_456,
input [18:0] Wgt_1_457,
input [18:0] Wgt_1_458,
input [18:0] Wgt_1_459,
input [18:0] Wgt_1_460,
input [18:0] Wgt_1_461,
input [18:0] Wgt_1_462,
input [18:0] Wgt_1_463,
input [18:0] Wgt_1_464,
input [18:0] Wgt_1_465,
input [18:0] Wgt_1_466,
input [18:0] Wgt_1_467,
input [18:0] Wgt_1_468,
input [18:0] Wgt_1_469,
input [18:0] Wgt_1_470,
input [18:0] Wgt_1_471,
input [18:0] Wgt_1_472,
input [18:0] Wgt_1_473,
input [18:0] Wgt_1_474,
input [18:0] Wgt_1_475,
input [18:0] Wgt_1_476,
input [18:0] Wgt_1_477,
input [18:0] Wgt_1_478,
input [18:0] Wgt_1_479,
input [18:0] Wgt_1_480,
input [18:0] Wgt_1_481,
input [18:0] Wgt_1_482,
input [18:0] Wgt_1_483,
input [18:0] Wgt_1_484,
input [18:0] Wgt_1_485,
input [18:0] Wgt_1_486,
input [18:0] Wgt_1_487,
input [18:0] Wgt_1_488,
input [18:0] Wgt_1_489,
input [18:0] Wgt_1_490,
input [18:0] Wgt_1_491,
input [18:0] Wgt_1_492,
input [18:0] Wgt_1_493,
input [18:0] Wgt_1_494,
input [18:0] Wgt_1_495,
input [18:0] Wgt_1_496,
input [18:0] Wgt_1_497,
input [18:0] Wgt_1_498,
input [18:0] Wgt_1_499,
input [18:0] Wgt_1_500,
input [18:0] Wgt_1_501,
input [18:0] Wgt_1_502,
input [18:0] Wgt_1_503,
input [18:0] Wgt_1_504,
input [18:0] Wgt_1_505,
input [18:0] Wgt_1_506,
input [18:0] Wgt_1_507,
input [18:0] Wgt_1_508,
input [18:0] Wgt_1_509,
input [18:0] Wgt_1_510,
input [18:0] Wgt_1_511,
input [18:0] Wgt_1_512,
input [18:0] Wgt_1_513,
input [18:0] Wgt_1_514,
input [18:0] Wgt_1_515,
input [18:0] Wgt_1_516,
input [18:0] Wgt_1_517,
input [18:0] Wgt_1_518,
input [18:0] Wgt_1_519,
input [18:0] Wgt_1_520,
input [18:0] Wgt_1_521,
input [18:0] Wgt_1_522,
input [18:0] Wgt_1_523,
input [18:0] Wgt_1_524,
input [18:0] Wgt_1_525,
input [18:0] Wgt_1_526,
input [18:0] Wgt_1_527,
input [18:0] Wgt_1_528,
input [18:0] Wgt_1_529,
input [18:0] Wgt_1_530,
input [18:0] Wgt_1_531,
input [18:0] Wgt_1_532,
input [18:0] Wgt_1_533,
input [18:0] Wgt_1_534,
input [18:0] Wgt_1_535,
input [18:0] Wgt_1_536,
input [18:0] Wgt_1_537,
input [18:0] Wgt_1_538,
input [18:0] Wgt_1_539,
input [18:0] Wgt_1_540,
input [18:0] Wgt_1_541,
input [18:0] Wgt_1_542,
input [18:0] Wgt_1_543,
input [18:0] Wgt_1_544,
input [18:0] Wgt_1_545,
input [18:0] Wgt_1_546,
input [18:0] Wgt_1_547,
input [18:0] Wgt_1_548,
input [18:0] Wgt_1_549,
input [18:0] Wgt_1_550,
input [18:0] Wgt_1_551,
input [18:0] Wgt_1_552,
input [18:0] Wgt_1_553,
input [18:0] Wgt_1_554,
input [18:0] Wgt_1_555,
input [18:0] Wgt_1_556,
input [18:0] Wgt_1_557,
input [18:0] Wgt_1_558,
input [18:0] Wgt_1_559,
input [18:0] Wgt_1_560,
input [18:0] Wgt_1_561,
input [18:0] Wgt_1_562,
input [18:0] Wgt_1_563,
input [18:0] Wgt_1_564,
input [18:0] Wgt_1_565,
input [18:0] Wgt_1_566,
input [18:0] Wgt_1_567,
input [18:0] Wgt_1_568,
input [18:0] Wgt_1_569,
input [18:0] Wgt_1_570,
input [18:0] Wgt_1_571,
input [18:0] Wgt_1_572,
input [18:0] Wgt_1_573,
input [18:0] Wgt_1_574,
input [18:0] Wgt_1_575,
input [18:0] Wgt_1_576,
input [18:0] Wgt_1_577,
input [18:0] Wgt_1_578,
input [18:0] Wgt_1_579,
input [18:0] Wgt_1_580,
input [18:0] Wgt_1_581,
input [18:0] Wgt_1_582,
input [18:0] Wgt_1_583,
input [18:0] Wgt_1_584,
input [18:0] Wgt_1_585,
input [18:0] Wgt_1_586,
input [18:0] Wgt_1_587,
input [18:0] Wgt_1_588,
input [18:0] Wgt_1_589,
input [18:0] Wgt_1_590,
input [18:0] Wgt_1_591,
input [18:0] Wgt_1_592,
input [18:0] Wgt_1_593,
input [18:0] Wgt_1_594,
input [18:0] Wgt_1_595,
input [18:0] Wgt_1_596,
input [18:0] Wgt_1_597,
input [18:0] Wgt_1_598,
input [18:0] Wgt_1_599,
input [18:0] Wgt_1_600,
input [18:0] Wgt_1_601,
input [18:0] Wgt_1_602,
input [18:0] Wgt_1_603,
input [18:0] Wgt_1_604,
input [18:0] Wgt_1_605,
input [18:0] Wgt_1_606,
input [18:0] Wgt_1_607,
input [18:0] Wgt_1_608,
input [18:0] Wgt_1_609,
input [18:0] Wgt_1_610,
input [18:0] Wgt_1_611,
input [18:0] Wgt_1_612,
input [18:0] Wgt_1_613,
input [18:0] Wgt_1_614,
input [18:0] Wgt_1_615,
input [18:0] Wgt_1_616,
input [18:0] Wgt_1_617,
input [18:0] Wgt_1_618,
input [18:0] Wgt_1_619,
input [18:0] Wgt_1_620,
input [18:0] Wgt_1_621,
input [18:0] Wgt_1_622,
input [18:0] Wgt_1_623,
input [18:0] Wgt_1_624,
input [18:0] Wgt_1_625,
input [18:0] Wgt_1_626,
input [18:0] Wgt_1_627,
input [18:0] Wgt_1_628,
input [18:0] Wgt_1_629,
input [18:0] Wgt_1_630,
input [18:0] Wgt_1_631,
input [18:0] Wgt_1_632,
input [18:0] Wgt_1_633,
input [18:0] Wgt_1_634,
input [18:0] Wgt_1_635,
input [18:0] Wgt_1_636,
input [18:0] Wgt_1_637,
input [18:0] Wgt_1_638,
input [18:0] Wgt_1_639,
input [18:0] Wgt_1_640,
input [18:0] Wgt_1_641,
input [18:0] Wgt_1_642,
input [18:0] Wgt_1_643,
input [18:0] Wgt_1_644,
input [18:0] Wgt_1_645,
input [18:0] Wgt_1_646,
input [18:0] Wgt_1_647,
input [18:0] Wgt_1_648,
input [18:0] Wgt_1_649,
input [18:0] Wgt_1_650,
input [18:0] Wgt_1_651,
input [18:0] Wgt_1_652,
input [18:0] Wgt_1_653,
input [18:0] Wgt_1_654,
input [18:0] Wgt_1_655,
input [18:0] Wgt_1_656,
input [18:0] Wgt_1_657,
input [18:0] Wgt_1_658,
input [18:0] Wgt_1_659,
input [18:0] Wgt_1_660,
input [18:0] Wgt_1_661,
input [18:0] Wgt_1_662,
input [18:0] Wgt_1_663,
input [18:0] Wgt_1_664,
input [18:0] Wgt_1_665,
input [18:0] Wgt_1_666,
input [18:0] Wgt_1_667,
input [18:0] Wgt_1_668,
input [18:0] Wgt_1_669,
input [18:0] Wgt_1_670,
input [18:0] Wgt_1_671,
input [18:0] Wgt_1_672,
input [18:0] Wgt_1_673,
input [18:0] Wgt_1_674,
input [18:0] Wgt_1_675,
input [18:0] Wgt_1_676,
input [18:0] Wgt_1_677,
input [18:0] Wgt_1_678,
input [18:0] Wgt_1_679,
input [18:0] Wgt_1_680,
input [18:0] Wgt_1_681,
input [18:0] Wgt_1_682,
input [18:0] Wgt_1_683,
input [18:0] Wgt_1_684,
input [18:0] Wgt_1_685,
input [18:0] Wgt_1_686,
input [18:0] Wgt_1_687,
input [18:0] Wgt_1_688,
input [18:0] Wgt_1_689,
input [18:0] Wgt_1_690,
input [18:0] Wgt_1_691,
input [18:0] Wgt_1_692,
input [18:0] Wgt_1_693,
input [18:0] Wgt_1_694,
input [18:0] Wgt_1_695,
input [18:0] Wgt_1_696,
input [18:0] Wgt_1_697,
input [18:0] Wgt_1_698,
input [18:0] Wgt_1_699,
input [18:0] Wgt_1_700,
input [18:0] Wgt_1_701,
input [18:0] Wgt_1_702,
input [18:0] Wgt_1_703,
input [18:0] Wgt_1_704,
input [18:0] Wgt_1_705,
input [18:0] Wgt_1_706,
input [18:0] Wgt_1_707,
input [18:0] Wgt_1_708,
input [18:0] Wgt_1_709,
input [18:0] Wgt_1_710,
input [18:0] Wgt_1_711,
input [18:0] Wgt_1_712,
input [18:0] Wgt_1_713,
input [18:0] Wgt_1_714,
input [18:0] Wgt_1_715,
input [18:0] Wgt_1_716,
input [18:0] Wgt_1_717,
input [18:0] Wgt_1_718,
input [18:0] Wgt_1_719,
input [18:0] Wgt_1_720,
input [18:0] Wgt_1_721,
input [18:0] Wgt_1_722,
input [18:0] Wgt_1_723,
input [18:0] Wgt_1_724,
input [18:0] Wgt_1_725,
input [18:0] Wgt_1_726,
input [18:0] Wgt_1_727,
input [18:0] Wgt_1_728,
input [18:0] Wgt_1_729,
input [18:0] Wgt_1_730,
input [18:0] Wgt_1_731,
input [18:0] Wgt_1_732,
input [18:0] Wgt_1_733,
input [18:0] Wgt_1_734,
input [18:0] Wgt_1_735,
input [18:0] Wgt_1_736,
input [18:0] Wgt_1_737,
input [18:0] Wgt_1_738,
input [18:0] Wgt_1_739,
input [18:0] Wgt_1_740,
input [18:0] Wgt_1_741,
input [18:0] Wgt_1_742,
input [18:0] Wgt_1_743,
input [18:0] Wgt_1_744,
input [18:0] Wgt_1_745,
input [18:0] Wgt_1_746,
input [18:0] Wgt_1_747,
input [18:0] Wgt_1_748,
input [18:0] Wgt_1_749,
input [18:0] Wgt_1_750,
input [18:0] Wgt_1_751,
input [18:0] Wgt_1_752,
input [18:0] Wgt_1_753,
input [18:0] Wgt_1_754,
input [18:0] Wgt_1_755,
input [18:0] Wgt_1_756,
input [18:0] Wgt_1_757,
input [18:0] Wgt_1_758,
input [18:0] Wgt_1_759,
input [18:0] Wgt_1_760,
input [18:0] Wgt_1_761,
input [18:0] Wgt_1_762,
input [18:0] Wgt_1_763,
input [18:0] Wgt_1_764,
input [18:0] Wgt_1_765,
input [18:0] Wgt_1_766,
input [18:0] Wgt_1_767,
input [18:0] Wgt_1_768,
input [18:0] Wgt_1_769,
input [18:0] Wgt_1_770,
input [18:0] Wgt_1_771,
input [18:0] Wgt_1_772,
input [18:0] Wgt_1_773,
input [18:0] Wgt_1_774,
input [18:0] Wgt_1_775,
input [18:0] Wgt_1_776,
input [18:0] Wgt_1_777,
input [18:0] Wgt_1_778,
input [18:0] Wgt_1_779,
input [18:0] Wgt_1_780,
input [18:0] Wgt_1_781,
input [18:0] Wgt_1_782,
input [18:0] Wgt_1_783,
input [18:0] Wgt_1_784,
input [18:0] Wgt_2_0,
input [18:0] Wgt_2_1,
input [18:0] Wgt_2_2,
input [18:0] Wgt_2_3,
input [18:0] Wgt_2_4,
input [18:0] Wgt_2_5,
input [18:0] Wgt_2_6,
input [18:0] Wgt_2_7,
input [18:0] Wgt_2_8,
input [18:0] Wgt_2_9,
input [18:0] Wgt_2_10,
input [18:0] Wgt_2_11,
input [18:0] Wgt_2_12,
input [18:0] Wgt_2_13,
input [18:0] Wgt_2_14,
input [18:0] Wgt_2_15,
input [18:0] Wgt_2_16,
input [18:0] Wgt_2_17,
input [18:0] Wgt_2_18,
input [18:0] Wgt_2_19,
input [18:0] Wgt_2_20,
input [18:0] Wgt_2_21,
input [18:0] Wgt_2_22,
input [18:0] Wgt_2_23,
input [18:0] Wgt_2_24,
input [18:0] Wgt_2_25,
input [18:0] Wgt_2_26,
input [18:0] Wgt_2_27,
input [18:0] Wgt_2_28,
input [18:0] Wgt_2_29,
input [18:0] Wgt_2_30,
input [18:0] Wgt_2_31,
input [18:0] Wgt_2_32,
input [18:0] Wgt_2_33,
input [18:0] Wgt_2_34,
input [18:0] Wgt_2_35,
input [18:0] Wgt_2_36,
input [18:0] Wgt_2_37,
input [18:0] Wgt_2_38,
input [18:0] Wgt_2_39,
input [18:0] Wgt_2_40,
input [18:0] Wgt_2_41,
input [18:0] Wgt_2_42,
input [18:0] Wgt_2_43,
input [18:0] Wgt_2_44,
input [18:0] Wgt_2_45,
input [18:0] Wgt_2_46,
input [18:0] Wgt_2_47,
input [18:0] Wgt_2_48,
input [18:0] Wgt_2_49,
input [18:0] Wgt_2_50,
input [18:0] Wgt_2_51,
input [18:0] Wgt_2_52,
input [18:0] Wgt_2_53,
input [18:0] Wgt_2_54,
input [18:0] Wgt_2_55,
input [18:0] Wgt_2_56,
input [18:0] Wgt_2_57,
input [18:0] Wgt_2_58,
input [18:0] Wgt_2_59,
input [18:0] Wgt_2_60,
input [18:0] Wgt_2_61,
input [18:0] Wgt_2_62,
input [18:0] Wgt_2_63,
input [18:0] Wgt_2_64,
input [18:0] Wgt_2_65,
input [18:0] Wgt_2_66,
input [18:0] Wgt_2_67,
input [18:0] Wgt_2_68,
input [18:0] Wgt_2_69,
input [18:0] Wgt_2_70,
input [18:0] Wgt_2_71,
input [18:0] Wgt_2_72,
input [18:0] Wgt_2_73,
input [18:0] Wgt_2_74,
input [18:0] Wgt_2_75,
input [18:0] Wgt_2_76,
input [18:0] Wgt_2_77,
input [18:0] Wgt_2_78,
input [18:0] Wgt_2_79,
input [18:0] Wgt_2_80,
input [18:0] Wgt_2_81,
input [18:0] Wgt_2_82,
input [18:0] Wgt_2_83,
input [18:0] Wgt_2_84,
input [18:0] Wgt_2_85,
input [18:0] Wgt_2_86,
input [18:0] Wgt_2_87,
input [18:0] Wgt_2_88,
input [18:0] Wgt_2_89,
input [18:0] Wgt_2_90,
input [18:0] Wgt_2_91,
input [18:0] Wgt_2_92,
input [18:0] Wgt_2_93,
input [18:0] Wgt_2_94,
input [18:0] Wgt_2_95,
input [18:0] Wgt_2_96,
input [18:0] Wgt_2_97,
input [18:0] Wgt_2_98,
input [18:0] Wgt_2_99,
input [18:0] Wgt_2_100,
input [18:0] Wgt_2_101,
input [18:0] Wgt_2_102,
input [18:0] Wgt_2_103,
input [18:0] Wgt_2_104,
input [18:0] Wgt_2_105,
input [18:0] Wgt_2_106,
input [18:0] Wgt_2_107,
input [18:0] Wgt_2_108,
input [18:0] Wgt_2_109,
input [18:0] Wgt_2_110,
input [18:0] Wgt_2_111,
input [18:0] Wgt_2_112,
input [18:0] Wgt_2_113,
input [18:0] Wgt_2_114,
input [18:0] Wgt_2_115,
input [18:0] Wgt_2_116,
input [18:0] Wgt_2_117,
input [18:0] Wgt_2_118,
input [18:0] Wgt_2_119,
input [18:0] Wgt_2_120,
input [18:0] Wgt_2_121,
input [18:0] Wgt_2_122,
input [18:0] Wgt_2_123,
input [18:0] Wgt_2_124,
input [18:0] Wgt_2_125,
input [18:0] Wgt_2_126,
input [18:0] Wgt_2_127,
input [18:0] Wgt_2_128,
input [18:0] Wgt_2_129,
input [18:0] Wgt_2_130,
input [18:0] Wgt_2_131,
input [18:0] Wgt_2_132,
input [18:0] Wgt_2_133,
input [18:0] Wgt_2_134,
input [18:0] Wgt_2_135,
input [18:0] Wgt_2_136,
input [18:0] Wgt_2_137,
input [18:0] Wgt_2_138,
input [18:0] Wgt_2_139,
input [18:0] Wgt_2_140,
input [18:0] Wgt_2_141,
input [18:0] Wgt_2_142,
input [18:0] Wgt_2_143,
input [18:0] Wgt_2_144,
input [18:0] Wgt_2_145,
input [18:0] Wgt_2_146,
input [18:0] Wgt_2_147,
input [18:0] Wgt_2_148,
input [18:0] Wgt_2_149,
input [18:0] Wgt_2_150,
input [18:0] Wgt_2_151,
input [18:0] Wgt_2_152,
input [18:0] Wgt_2_153,
input [18:0] Wgt_2_154,
input [18:0] Wgt_2_155,
input [18:0] Wgt_2_156,
input [18:0] Wgt_2_157,
input [18:0] Wgt_2_158,
input [18:0] Wgt_2_159,
input [18:0] Wgt_2_160,
input [18:0] Wgt_2_161,
input [18:0] Wgt_2_162,
input [18:0] Wgt_2_163,
input [18:0] Wgt_2_164,
input [18:0] Wgt_2_165,
input [18:0] Wgt_2_166,
input [18:0] Wgt_2_167,
input [18:0] Wgt_2_168,
input [18:0] Wgt_2_169,
input [18:0] Wgt_2_170,
input [18:0] Wgt_2_171,
input [18:0] Wgt_2_172,
input [18:0] Wgt_2_173,
input [18:0] Wgt_2_174,
input [18:0] Wgt_2_175,
input [18:0] Wgt_2_176,
input [18:0] Wgt_2_177,
input [18:0] Wgt_2_178,
input [18:0] Wgt_2_179,
input [18:0] Wgt_2_180,
input [18:0] Wgt_2_181,
input [18:0] Wgt_2_182,
input [18:0] Wgt_2_183,
input [18:0] Wgt_2_184,
input [18:0] Wgt_2_185,
input [18:0] Wgt_2_186,
input [18:0] Wgt_2_187,
input [18:0] Wgt_2_188,
input [18:0] Wgt_2_189,
input [18:0] Wgt_2_190,
input [18:0] Wgt_2_191,
input [18:0] Wgt_2_192,
input [18:0] Wgt_2_193,
input [18:0] Wgt_2_194,
input [18:0] Wgt_2_195,
input [18:0] Wgt_2_196,
input [18:0] Wgt_2_197,
input [18:0] Wgt_2_198,
input [18:0] Wgt_2_199,
input [18:0] Wgt_2_200,
input [18:0] Wgt_2_201,
input [18:0] Wgt_2_202,
input [18:0] Wgt_2_203,
input [18:0] Wgt_2_204,
input [18:0] Wgt_2_205,
input [18:0] Wgt_2_206,
input [18:0] Wgt_2_207,
input [18:0] Wgt_2_208,
input [18:0] Wgt_2_209,
input [18:0] Wgt_2_210,
input [18:0] Wgt_2_211,
input [18:0] Wgt_2_212,
input [18:0] Wgt_2_213,
input [18:0] Wgt_2_214,
input [18:0] Wgt_2_215,
input [18:0] Wgt_2_216,
input [18:0] Wgt_2_217,
input [18:0] Wgt_2_218,
input [18:0] Wgt_2_219,
input [18:0] Wgt_2_220,
input [18:0] Wgt_2_221,
input [18:0] Wgt_2_222,
input [18:0] Wgt_2_223,
input [18:0] Wgt_2_224,
input [18:0] Wgt_2_225,
input [18:0] Wgt_2_226,
input [18:0] Wgt_2_227,
input [18:0] Wgt_2_228,
input [18:0] Wgt_2_229,
input [18:0] Wgt_2_230,
input [18:0] Wgt_2_231,
input [18:0] Wgt_2_232,
input [18:0] Wgt_2_233,
input [18:0] Wgt_2_234,
input [18:0] Wgt_2_235,
input [18:0] Wgt_2_236,
input [18:0] Wgt_2_237,
input [18:0] Wgt_2_238,
input [18:0] Wgt_2_239,
input [18:0] Wgt_2_240,
input [18:0] Wgt_2_241,
input [18:0] Wgt_2_242,
input [18:0] Wgt_2_243,
input [18:0] Wgt_2_244,
input [18:0] Wgt_2_245,
input [18:0] Wgt_2_246,
input [18:0] Wgt_2_247,
input [18:0] Wgt_2_248,
input [18:0] Wgt_2_249,
input [18:0] Wgt_2_250,
input [18:0] Wgt_2_251,
input [18:0] Wgt_2_252,
input [18:0] Wgt_2_253,
input [18:0] Wgt_2_254,
input [18:0] Wgt_2_255,
input [18:0] Wgt_2_256,
input [18:0] Wgt_2_257,
input [18:0] Wgt_2_258,
input [18:0] Wgt_2_259,
input [18:0] Wgt_2_260,
input [18:0] Wgt_2_261,
input [18:0] Wgt_2_262,
input [18:0] Wgt_2_263,
input [18:0] Wgt_2_264,
input [18:0] Wgt_2_265,
input [18:0] Wgt_2_266,
input [18:0] Wgt_2_267,
input [18:0] Wgt_2_268,
input [18:0] Wgt_2_269,
input [18:0] Wgt_2_270,
input [18:0] Wgt_2_271,
input [18:0] Wgt_2_272,
input [18:0] Wgt_2_273,
input [18:0] Wgt_2_274,
input [18:0] Wgt_2_275,
input [18:0] Wgt_2_276,
input [18:0] Wgt_2_277,
input [18:0] Wgt_2_278,
input [18:0] Wgt_2_279,
input [18:0] Wgt_2_280,
input [18:0] Wgt_2_281,
input [18:0] Wgt_2_282,
input [18:0] Wgt_2_283,
input [18:0] Wgt_2_284,
input [18:0] Wgt_2_285,
input [18:0] Wgt_2_286,
input [18:0] Wgt_2_287,
input [18:0] Wgt_2_288,
input [18:0] Wgt_2_289,
input [18:0] Wgt_2_290,
input [18:0] Wgt_2_291,
input [18:0] Wgt_2_292,
input [18:0] Wgt_2_293,
input [18:0] Wgt_2_294,
input [18:0] Wgt_2_295,
input [18:0] Wgt_2_296,
input [18:0] Wgt_2_297,
input [18:0] Wgt_2_298,
input [18:0] Wgt_2_299,
input [18:0] Wgt_2_300,
input [18:0] Wgt_2_301,
input [18:0] Wgt_2_302,
input [18:0] Wgt_2_303,
input [18:0] Wgt_2_304,
input [18:0] Wgt_2_305,
input [18:0] Wgt_2_306,
input [18:0] Wgt_2_307,
input [18:0] Wgt_2_308,
input [18:0] Wgt_2_309,
input [18:0] Wgt_2_310,
input [18:0] Wgt_2_311,
input [18:0] Wgt_2_312,
input [18:0] Wgt_2_313,
input [18:0] Wgt_2_314,
input [18:0] Wgt_2_315,
input [18:0] Wgt_2_316,
input [18:0] Wgt_2_317,
input [18:0] Wgt_2_318,
input [18:0] Wgt_2_319,
input [18:0] Wgt_2_320,
input [18:0] Wgt_2_321,
input [18:0] Wgt_2_322,
input [18:0] Wgt_2_323,
input [18:0] Wgt_2_324,
input [18:0] Wgt_2_325,
input [18:0] Wgt_2_326,
input [18:0] Wgt_2_327,
input [18:0] Wgt_2_328,
input [18:0] Wgt_2_329,
input [18:0] Wgt_2_330,
input [18:0] Wgt_2_331,
input [18:0] Wgt_2_332,
input [18:0] Wgt_2_333,
input [18:0] Wgt_2_334,
input [18:0] Wgt_2_335,
input [18:0] Wgt_2_336,
input [18:0] Wgt_2_337,
input [18:0] Wgt_2_338,
input [18:0] Wgt_2_339,
input [18:0] Wgt_2_340,
input [18:0] Wgt_2_341,
input [18:0] Wgt_2_342,
input [18:0] Wgt_2_343,
input [18:0] Wgt_2_344,
input [18:0] Wgt_2_345,
input [18:0] Wgt_2_346,
input [18:0] Wgt_2_347,
input [18:0] Wgt_2_348,
input [18:0] Wgt_2_349,
input [18:0] Wgt_2_350,
input [18:0] Wgt_2_351,
input [18:0] Wgt_2_352,
input [18:0] Wgt_2_353,
input [18:0] Wgt_2_354,
input [18:0] Wgt_2_355,
input [18:0] Wgt_2_356,
input [18:0] Wgt_2_357,
input [18:0] Wgt_2_358,
input [18:0] Wgt_2_359,
input [18:0] Wgt_2_360,
input [18:0] Wgt_2_361,
input [18:0] Wgt_2_362,
input [18:0] Wgt_2_363,
input [18:0] Wgt_2_364,
input [18:0] Wgt_2_365,
input [18:0] Wgt_2_366,
input [18:0] Wgt_2_367,
input [18:0] Wgt_2_368,
input [18:0] Wgt_2_369,
input [18:0] Wgt_2_370,
input [18:0] Wgt_2_371,
input [18:0] Wgt_2_372,
input [18:0] Wgt_2_373,
input [18:0] Wgt_2_374,
input [18:0] Wgt_2_375,
input [18:0] Wgt_2_376,
input [18:0] Wgt_2_377,
input [18:0] Wgt_2_378,
input [18:0] Wgt_2_379,
input [18:0] Wgt_2_380,
input [18:0] Wgt_2_381,
input [18:0] Wgt_2_382,
input [18:0] Wgt_2_383,
input [18:0] Wgt_2_384,
input [18:0] Wgt_2_385,
input [18:0] Wgt_2_386,
input [18:0] Wgt_2_387,
input [18:0] Wgt_2_388,
input [18:0] Wgt_2_389,
input [18:0] Wgt_2_390,
input [18:0] Wgt_2_391,
input [18:0] Wgt_2_392,
input [18:0] Wgt_2_393,
input [18:0] Wgt_2_394,
input [18:0] Wgt_2_395,
input [18:0] Wgt_2_396,
input [18:0] Wgt_2_397,
input [18:0] Wgt_2_398,
input [18:0] Wgt_2_399,
input [18:0] Wgt_2_400,
input [18:0] Wgt_2_401,
input [18:0] Wgt_2_402,
input [18:0] Wgt_2_403,
input [18:0] Wgt_2_404,
input [18:0] Wgt_2_405,
input [18:0] Wgt_2_406,
input [18:0] Wgt_2_407,
input [18:0] Wgt_2_408,
input [18:0] Wgt_2_409,
input [18:0] Wgt_2_410,
input [18:0] Wgt_2_411,
input [18:0] Wgt_2_412,
input [18:0] Wgt_2_413,
input [18:0] Wgt_2_414,
input [18:0] Wgt_2_415,
input [18:0] Wgt_2_416,
input [18:0] Wgt_2_417,
input [18:0] Wgt_2_418,
input [18:0] Wgt_2_419,
input [18:0] Wgt_2_420,
input [18:0] Wgt_2_421,
input [18:0] Wgt_2_422,
input [18:0] Wgt_2_423,
input [18:0] Wgt_2_424,
input [18:0] Wgt_2_425,
input [18:0] Wgt_2_426,
input [18:0] Wgt_2_427,
input [18:0] Wgt_2_428,
input [18:0] Wgt_2_429,
input [18:0] Wgt_2_430,
input [18:0] Wgt_2_431,
input [18:0] Wgt_2_432,
input [18:0] Wgt_2_433,
input [18:0] Wgt_2_434,
input [18:0] Wgt_2_435,
input [18:0] Wgt_2_436,
input [18:0] Wgt_2_437,
input [18:0] Wgt_2_438,
input [18:0] Wgt_2_439,
input [18:0] Wgt_2_440,
input [18:0] Wgt_2_441,
input [18:0] Wgt_2_442,
input [18:0] Wgt_2_443,
input [18:0] Wgt_2_444,
input [18:0] Wgt_2_445,
input [18:0] Wgt_2_446,
input [18:0] Wgt_2_447,
input [18:0] Wgt_2_448,
input [18:0] Wgt_2_449,
input [18:0] Wgt_2_450,
input [18:0] Wgt_2_451,
input [18:0] Wgt_2_452,
input [18:0] Wgt_2_453,
input [18:0] Wgt_2_454,
input [18:0] Wgt_2_455,
input [18:0] Wgt_2_456,
input [18:0] Wgt_2_457,
input [18:0] Wgt_2_458,
input [18:0] Wgt_2_459,
input [18:0] Wgt_2_460,
input [18:0] Wgt_2_461,
input [18:0] Wgt_2_462,
input [18:0] Wgt_2_463,
input [18:0] Wgt_2_464,
input [18:0] Wgt_2_465,
input [18:0] Wgt_2_466,
input [18:0] Wgt_2_467,
input [18:0] Wgt_2_468,
input [18:0] Wgt_2_469,
input [18:0] Wgt_2_470,
input [18:0] Wgt_2_471,
input [18:0] Wgt_2_472,
input [18:0] Wgt_2_473,
input [18:0] Wgt_2_474,
input [18:0] Wgt_2_475,
input [18:0] Wgt_2_476,
input [18:0] Wgt_2_477,
input [18:0] Wgt_2_478,
input [18:0] Wgt_2_479,
input [18:0] Wgt_2_480,
input [18:0] Wgt_2_481,
input [18:0] Wgt_2_482,
input [18:0] Wgt_2_483,
input [18:0] Wgt_2_484,
input [18:0] Wgt_2_485,
input [18:0] Wgt_2_486,
input [18:0] Wgt_2_487,
input [18:0] Wgt_2_488,
input [18:0] Wgt_2_489,
input [18:0] Wgt_2_490,
input [18:0] Wgt_2_491,
input [18:0] Wgt_2_492,
input [18:0] Wgt_2_493,
input [18:0] Wgt_2_494,
input [18:0] Wgt_2_495,
input [18:0] Wgt_2_496,
input [18:0] Wgt_2_497,
input [18:0] Wgt_2_498,
input [18:0] Wgt_2_499,
input [18:0] Wgt_2_500,
input [18:0] Wgt_2_501,
input [18:0] Wgt_2_502,
input [18:0] Wgt_2_503,
input [18:0] Wgt_2_504,
input [18:0] Wgt_2_505,
input [18:0] Wgt_2_506,
input [18:0] Wgt_2_507,
input [18:0] Wgt_2_508,
input [18:0] Wgt_2_509,
input [18:0] Wgt_2_510,
input [18:0] Wgt_2_511,
input [18:0] Wgt_2_512,
input [18:0] Wgt_2_513,
input [18:0] Wgt_2_514,
input [18:0] Wgt_2_515,
input [18:0] Wgt_2_516,
input [18:0] Wgt_2_517,
input [18:0] Wgt_2_518,
input [18:0] Wgt_2_519,
input [18:0] Wgt_2_520,
input [18:0] Wgt_2_521,
input [18:0] Wgt_2_522,
input [18:0] Wgt_2_523,
input [18:0] Wgt_2_524,
input [18:0] Wgt_2_525,
input [18:0] Wgt_2_526,
input [18:0] Wgt_2_527,
input [18:0] Wgt_2_528,
input [18:0] Wgt_2_529,
input [18:0] Wgt_2_530,
input [18:0] Wgt_2_531,
input [18:0] Wgt_2_532,
input [18:0] Wgt_2_533,
input [18:0] Wgt_2_534,
input [18:0] Wgt_2_535,
input [18:0] Wgt_2_536,
input [18:0] Wgt_2_537,
input [18:0] Wgt_2_538,
input [18:0] Wgt_2_539,
input [18:0] Wgt_2_540,
input [18:0] Wgt_2_541,
input [18:0] Wgt_2_542,
input [18:0] Wgt_2_543,
input [18:0] Wgt_2_544,
input [18:0] Wgt_2_545,
input [18:0] Wgt_2_546,
input [18:0] Wgt_2_547,
input [18:0] Wgt_2_548,
input [18:0] Wgt_2_549,
input [18:0] Wgt_2_550,
input [18:0] Wgt_2_551,
input [18:0] Wgt_2_552,
input [18:0] Wgt_2_553,
input [18:0] Wgt_2_554,
input [18:0] Wgt_2_555,
input [18:0] Wgt_2_556,
input [18:0] Wgt_2_557,
input [18:0] Wgt_2_558,
input [18:0] Wgt_2_559,
input [18:0] Wgt_2_560,
input [18:0] Wgt_2_561,
input [18:0] Wgt_2_562,
input [18:0] Wgt_2_563,
input [18:0] Wgt_2_564,
input [18:0] Wgt_2_565,
input [18:0] Wgt_2_566,
input [18:0] Wgt_2_567,
input [18:0] Wgt_2_568,
input [18:0] Wgt_2_569,
input [18:0] Wgt_2_570,
input [18:0] Wgt_2_571,
input [18:0] Wgt_2_572,
input [18:0] Wgt_2_573,
input [18:0] Wgt_2_574,
input [18:0] Wgt_2_575,
input [18:0] Wgt_2_576,
input [18:0] Wgt_2_577,
input [18:0] Wgt_2_578,
input [18:0] Wgt_2_579,
input [18:0] Wgt_2_580,
input [18:0] Wgt_2_581,
input [18:0] Wgt_2_582,
input [18:0] Wgt_2_583,
input [18:0] Wgt_2_584,
input [18:0] Wgt_2_585,
input [18:0] Wgt_2_586,
input [18:0] Wgt_2_587,
input [18:0] Wgt_2_588,
input [18:0] Wgt_2_589,
input [18:0] Wgt_2_590,
input [18:0] Wgt_2_591,
input [18:0] Wgt_2_592,
input [18:0] Wgt_2_593,
input [18:0] Wgt_2_594,
input [18:0] Wgt_2_595,
input [18:0] Wgt_2_596,
input [18:0] Wgt_2_597,
input [18:0] Wgt_2_598,
input [18:0] Wgt_2_599,
input [18:0] Wgt_2_600,
input [18:0] Wgt_2_601,
input [18:0] Wgt_2_602,
input [18:0] Wgt_2_603,
input [18:0] Wgt_2_604,
input [18:0] Wgt_2_605,
input [18:0] Wgt_2_606,
input [18:0] Wgt_2_607,
input [18:0] Wgt_2_608,
input [18:0] Wgt_2_609,
input [18:0] Wgt_2_610,
input [18:0] Wgt_2_611,
input [18:0] Wgt_2_612,
input [18:0] Wgt_2_613,
input [18:0] Wgt_2_614,
input [18:0] Wgt_2_615,
input [18:0] Wgt_2_616,
input [18:0] Wgt_2_617,
input [18:0] Wgt_2_618,
input [18:0] Wgt_2_619,
input [18:0] Wgt_2_620,
input [18:0] Wgt_2_621,
input [18:0] Wgt_2_622,
input [18:0] Wgt_2_623,
input [18:0] Wgt_2_624,
input [18:0] Wgt_2_625,
input [18:0] Wgt_2_626,
input [18:0] Wgt_2_627,
input [18:0] Wgt_2_628,
input [18:0] Wgt_2_629,
input [18:0] Wgt_2_630,
input [18:0] Wgt_2_631,
input [18:0] Wgt_2_632,
input [18:0] Wgt_2_633,
input [18:0] Wgt_2_634,
input [18:0] Wgt_2_635,
input [18:0] Wgt_2_636,
input [18:0] Wgt_2_637,
input [18:0] Wgt_2_638,
input [18:0] Wgt_2_639,
input [18:0] Wgt_2_640,
input [18:0] Wgt_2_641,
input [18:0] Wgt_2_642,
input [18:0] Wgt_2_643,
input [18:0] Wgt_2_644,
input [18:0] Wgt_2_645,
input [18:0] Wgt_2_646,
input [18:0] Wgt_2_647,
input [18:0] Wgt_2_648,
input [18:0] Wgt_2_649,
input [18:0] Wgt_2_650,
input [18:0] Wgt_2_651,
input [18:0] Wgt_2_652,
input [18:0] Wgt_2_653,
input [18:0] Wgt_2_654,
input [18:0] Wgt_2_655,
input [18:0] Wgt_2_656,
input [18:0] Wgt_2_657,
input [18:0] Wgt_2_658,
input [18:0] Wgt_2_659,
input [18:0] Wgt_2_660,
input [18:0] Wgt_2_661,
input [18:0] Wgt_2_662,
input [18:0] Wgt_2_663,
input [18:0] Wgt_2_664,
input [18:0] Wgt_2_665,
input [18:0] Wgt_2_666,
input [18:0] Wgt_2_667,
input [18:0] Wgt_2_668,
input [18:0] Wgt_2_669,
input [18:0] Wgt_2_670,
input [18:0] Wgt_2_671,
input [18:0] Wgt_2_672,
input [18:0] Wgt_2_673,
input [18:0] Wgt_2_674,
input [18:0] Wgt_2_675,
input [18:0] Wgt_2_676,
input [18:0] Wgt_2_677,
input [18:0] Wgt_2_678,
input [18:0] Wgt_2_679,
input [18:0] Wgt_2_680,
input [18:0] Wgt_2_681,
input [18:0] Wgt_2_682,
input [18:0] Wgt_2_683,
input [18:0] Wgt_2_684,
input [18:0] Wgt_2_685,
input [18:0] Wgt_2_686,
input [18:0] Wgt_2_687,
input [18:0] Wgt_2_688,
input [18:0] Wgt_2_689,
input [18:0] Wgt_2_690,
input [18:0] Wgt_2_691,
input [18:0] Wgt_2_692,
input [18:0] Wgt_2_693,
input [18:0] Wgt_2_694,
input [18:0] Wgt_2_695,
input [18:0] Wgt_2_696,
input [18:0] Wgt_2_697,
input [18:0] Wgt_2_698,
input [18:0] Wgt_2_699,
input [18:0] Wgt_2_700,
input [18:0] Wgt_2_701,
input [18:0] Wgt_2_702,
input [18:0] Wgt_2_703,
input [18:0] Wgt_2_704,
input [18:0] Wgt_2_705,
input [18:0] Wgt_2_706,
input [18:0] Wgt_2_707,
input [18:0] Wgt_2_708,
input [18:0] Wgt_2_709,
input [18:0] Wgt_2_710,
input [18:0] Wgt_2_711,
input [18:0] Wgt_2_712,
input [18:0] Wgt_2_713,
input [18:0] Wgt_2_714,
input [18:0] Wgt_2_715,
input [18:0] Wgt_2_716,
input [18:0] Wgt_2_717,
input [18:0] Wgt_2_718,
input [18:0] Wgt_2_719,
input [18:0] Wgt_2_720,
input [18:0] Wgt_2_721,
input [18:0] Wgt_2_722,
input [18:0] Wgt_2_723,
input [18:0] Wgt_2_724,
input [18:0] Wgt_2_725,
input [18:0] Wgt_2_726,
input [18:0] Wgt_2_727,
input [18:0] Wgt_2_728,
input [18:0] Wgt_2_729,
input [18:0] Wgt_2_730,
input [18:0] Wgt_2_731,
input [18:0] Wgt_2_732,
input [18:0] Wgt_2_733,
input [18:0] Wgt_2_734,
input [18:0] Wgt_2_735,
input [18:0] Wgt_2_736,
input [18:0] Wgt_2_737,
input [18:0] Wgt_2_738,
input [18:0] Wgt_2_739,
input [18:0] Wgt_2_740,
input [18:0] Wgt_2_741,
input [18:0] Wgt_2_742,
input [18:0] Wgt_2_743,
input [18:0] Wgt_2_744,
input [18:0] Wgt_2_745,
input [18:0] Wgt_2_746,
input [18:0] Wgt_2_747,
input [18:0] Wgt_2_748,
input [18:0] Wgt_2_749,
input [18:0] Wgt_2_750,
input [18:0] Wgt_2_751,
input [18:0] Wgt_2_752,
input [18:0] Wgt_2_753,
input [18:0] Wgt_2_754,
input [18:0] Wgt_2_755,
input [18:0] Wgt_2_756,
input [18:0] Wgt_2_757,
input [18:0] Wgt_2_758,
input [18:0] Wgt_2_759,
input [18:0] Wgt_2_760,
input [18:0] Wgt_2_761,
input [18:0] Wgt_2_762,
input [18:0] Wgt_2_763,
input [18:0] Wgt_2_764,
input [18:0] Wgt_2_765,
input [18:0] Wgt_2_766,
input [18:0] Wgt_2_767,
input [18:0] Wgt_2_768,
input [18:0] Wgt_2_769,
input [18:0] Wgt_2_770,
input [18:0] Wgt_2_771,
input [18:0] Wgt_2_772,
input [18:0] Wgt_2_773,
input [18:0] Wgt_2_774,
input [18:0] Wgt_2_775,
input [18:0] Wgt_2_776,
input [18:0] Wgt_2_777,
input [18:0] Wgt_2_778,
input [18:0] Wgt_2_779,
input [18:0] Wgt_2_780,
input [18:0] Wgt_2_781,
input [18:0] Wgt_2_782,
input [18:0] Wgt_2_783,
input [18:0] Wgt_2_784,
input [18:0] Wgt_3_0,
input [18:0] Wgt_3_1,
input [18:0] Wgt_3_2,
input [18:0] Wgt_3_3,
input [18:0] Wgt_3_4,
input [18:0] Wgt_3_5,
input [18:0] Wgt_3_6,
input [18:0] Wgt_3_7,
input [18:0] Wgt_3_8,
input [18:0] Wgt_3_9,
input [18:0] Wgt_3_10,
input [18:0] Wgt_3_11,
input [18:0] Wgt_3_12,
input [18:0] Wgt_3_13,
input [18:0] Wgt_3_14,
input [18:0] Wgt_3_15,
input [18:0] Wgt_3_16,
input [18:0] Wgt_3_17,
input [18:0] Wgt_3_18,
input [18:0] Wgt_3_19,
input [18:0] Wgt_3_20,
input [18:0] Wgt_3_21,
input [18:0] Wgt_3_22,
input [18:0] Wgt_3_23,
input [18:0] Wgt_3_24,
input [18:0] Wgt_3_25,
input [18:0] Wgt_3_26,
input [18:0] Wgt_3_27,
input [18:0] Wgt_3_28,
input [18:0] Wgt_3_29,
input [18:0] Wgt_3_30,
input [18:0] Wgt_3_31,
input [18:0] Wgt_3_32,
input [18:0] Wgt_3_33,
input [18:0] Wgt_3_34,
input [18:0] Wgt_3_35,
input [18:0] Wgt_3_36,
input [18:0] Wgt_3_37,
input [18:0] Wgt_3_38,
input [18:0] Wgt_3_39,
input [18:0] Wgt_3_40,
input [18:0] Wgt_3_41,
input [18:0] Wgt_3_42,
input [18:0] Wgt_3_43,
input [18:0] Wgt_3_44,
input [18:0] Wgt_3_45,
input [18:0] Wgt_3_46,
input [18:0] Wgt_3_47,
input [18:0] Wgt_3_48,
input [18:0] Wgt_3_49,
input [18:0] Wgt_3_50,
input [18:0] Wgt_3_51,
input [18:0] Wgt_3_52,
input [18:0] Wgt_3_53,
input [18:0] Wgt_3_54,
input [18:0] Wgt_3_55,
input [18:0] Wgt_3_56,
input [18:0] Wgt_3_57,
input [18:0] Wgt_3_58,
input [18:0] Wgt_3_59,
input [18:0] Wgt_3_60,
input [18:0] Wgt_3_61,
input [18:0] Wgt_3_62,
input [18:0] Wgt_3_63,
input [18:0] Wgt_3_64,
input [18:0] Wgt_3_65,
input [18:0] Wgt_3_66,
input [18:0] Wgt_3_67,
input [18:0] Wgt_3_68,
input [18:0] Wgt_3_69,
input [18:0] Wgt_3_70,
input [18:0] Wgt_3_71,
input [18:0] Wgt_3_72,
input [18:0] Wgt_3_73,
input [18:0] Wgt_3_74,
input [18:0] Wgt_3_75,
input [18:0] Wgt_3_76,
input [18:0] Wgt_3_77,
input [18:0] Wgt_3_78,
input [18:0] Wgt_3_79,
input [18:0] Wgt_3_80,
input [18:0] Wgt_3_81,
input [18:0] Wgt_3_82,
input [18:0] Wgt_3_83,
input [18:0] Wgt_3_84,
input [18:0] Wgt_3_85,
input [18:0] Wgt_3_86,
input [18:0] Wgt_3_87,
input [18:0] Wgt_3_88,
input [18:0] Wgt_3_89,
input [18:0] Wgt_3_90,
input [18:0] Wgt_3_91,
input [18:0] Wgt_3_92,
input [18:0] Wgt_3_93,
input [18:0] Wgt_3_94,
input [18:0] Wgt_3_95,
input [18:0] Wgt_3_96,
input [18:0] Wgt_3_97,
input [18:0] Wgt_3_98,
input [18:0] Wgt_3_99,
input [18:0] Wgt_3_100,
input [18:0] Wgt_3_101,
input [18:0] Wgt_3_102,
input [18:0] Wgt_3_103,
input [18:0] Wgt_3_104,
input [18:0] Wgt_3_105,
input [18:0] Wgt_3_106,
input [18:0] Wgt_3_107,
input [18:0] Wgt_3_108,
input [18:0] Wgt_3_109,
input [18:0] Wgt_3_110,
input [18:0] Wgt_3_111,
input [18:0] Wgt_3_112,
input [18:0] Wgt_3_113,
input [18:0] Wgt_3_114,
input [18:0] Wgt_3_115,
input [18:0] Wgt_3_116,
input [18:0] Wgt_3_117,
input [18:0] Wgt_3_118,
input [18:0] Wgt_3_119,
input [18:0] Wgt_3_120,
input [18:0] Wgt_3_121,
input [18:0] Wgt_3_122,
input [18:0] Wgt_3_123,
input [18:0] Wgt_3_124,
input [18:0] Wgt_3_125,
input [18:0] Wgt_3_126,
input [18:0] Wgt_3_127,
input [18:0] Wgt_3_128,
input [18:0] Wgt_3_129,
input [18:0] Wgt_3_130,
input [18:0] Wgt_3_131,
input [18:0] Wgt_3_132,
input [18:0] Wgt_3_133,
input [18:0] Wgt_3_134,
input [18:0] Wgt_3_135,
input [18:0] Wgt_3_136,
input [18:0] Wgt_3_137,
input [18:0] Wgt_3_138,
input [18:0] Wgt_3_139,
input [18:0] Wgt_3_140,
input [18:0] Wgt_3_141,
input [18:0] Wgt_3_142,
input [18:0] Wgt_3_143,
input [18:0] Wgt_3_144,
input [18:0] Wgt_3_145,
input [18:0] Wgt_3_146,
input [18:0] Wgt_3_147,
input [18:0] Wgt_3_148,
input [18:0] Wgt_3_149,
input [18:0] Wgt_3_150,
input [18:0] Wgt_3_151,
input [18:0] Wgt_3_152,
input [18:0] Wgt_3_153,
input [18:0] Wgt_3_154,
input [18:0] Wgt_3_155,
input [18:0] Wgt_3_156,
input [18:0] Wgt_3_157,
input [18:0] Wgt_3_158,
input [18:0] Wgt_3_159,
input [18:0] Wgt_3_160,
input [18:0] Wgt_3_161,
input [18:0] Wgt_3_162,
input [18:0] Wgt_3_163,
input [18:0] Wgt_3_164,
input [18:0] Wgt_3_165,
input [18:0] Wgt_3_166,
input [18:0] Wgt_3_167,
input [18:0] Wgt_3_168,
input [18:0] Wgt_3_169,
input [18:0] Wgt_3_170,
input [18:0] Wgt_3_171,
input [18:0] Wgt_3_172,
input [18:0] Wgt_3_173,
input [18:0] Wgt_3_174,
input [18:0] Wgt_3_175,
input [18:0] Wgt_3_176,
input [18:0] Wgt_3_177,
input [18:0] Wgt_3_178,
input [18:0] Wgt_3_179,
input [18:0] Wgt_3_180,
input [18:0] Wgt_3_181,
input [18:0] Wgt_3_182,
input [18:0] Wgt_3_183,
input [18:0] Wgt_3_184,
input [18:0] Wgt_3_185,
input [18:0] Wgt_3_186,
input [18:0] Wgt_3_187,
input [18:0] Wgt_3_188,
input [18:0] Wgt_3_189,
input [18:0] Wgt_3_190,
input [18:0] Wgt_3_191,
input [18:0] Wgt_3_192,
input [18:0] Wgt_3_193,
input [18:0] Wgt_3_194,
input [18:0] Wgt_3_195,
input [18:0] Wgt_3_196,
input [18:0] Wgt_3_197,
input [18:0] Wgt_3_198,
input [18:0] Wgt_3_199,
input [18:0] Wgt_3_200,
input [18:0] Wgt_3_201,
input [18:0] Wgt_3_202,
input [18:0] Wgt_3_203,
input [18:0] Wgt_3_204,
input [18:0] Wgt_3_205,
input [18:0] Wgt_3_206,
input [18:0] Wgt_3_207,
input [18:0] Wgt_3_208,
input [18:0] Wgt_3_209,
input [18:0] Wgt_3_210,
input [18:0] Wgt_3_211,
input [18:0] Wgt_3_212,
input [18:0] Wgt_3_213,
input [18:0] Wgt_3_214,
input [18:0] Wgt_3_215,
input [18:0] Wgt_3_216,
input [18:0] Wgt_3_217,
input [18:0] Wgt_3_218,
input [18:0] Wgt_3_219,
input [18:0] Wgt_3_220,
input [18:0] Wgt_3_221,
input [18:0] Wgt_3_222,
input [18:0] Wgt_3_223,
input [18:0] Wgt_3_224,
input [18:0] Wgt_3_225,
input [18:0] Wgt_3_226,
input [18:0] Wgt_3_227,
input [18:0] Wgt_3_228,
input [18:0] Wgt_3_229,
input [18:0] Wgt_3_230,
input [18:0] Wgt_3_231,
input [18:0] Wgt_3_232,
input [18:0] Wgt_3_233,
input [18:0] Wgt_3_234,
input [18:0] Wgt_3_235,
input [18:0] Wgt_3_236,
input [18:0] Wgt_3_237,
input [18:0] Wgt_3_238,
input [18:0] Wgt_3_239,
input [18:0] Wgt_3_240,
input [18:0] Wgt_3_241,
input [18:0] Wgt_3_242,
input [18:0] Wgt_3_243,
input [18:0] Wgt_3_244,
input [18:0] Wgt_3_245,
input [18:0] Wgt_3_246,
input [18:0] Wgt_3_247,
input [18:0] Wgt_3_248,
input [18:0] Wgt_3_249,
input [18:0] Wgt_3_250,
input [18:0] Wgt_3_251,
input [18:0] Wgt_3_252,
input [18:0] Wgt_3_253,
input [18:0] Wgt_3_254,
input [18:0] Wgt_3_255,
input [18:0] Wgt_3_256,
input [18:0] Wgt_3_257,
input [18:0] Wgt_3_258,
input [18:0] Wgt_3_259,
input [18:0] Wgt_3_260,
input [18:0] Wgt_3_261,
input [18:0] Wgt_3_262,
input [18:0] Wgt_3_263,
input [18:0] Wgt_3_264,
input [18:0] Wgt_3_265,
input [18:0] Wgt_3_266,
input [18:0] Wgt_3_267,
input [18:0] Wgt_3_268,
input [18:0] Wgt_3_269,
input [18:0] Wgt_3_270,
input [18:0] Wgt_3_271,
input [18:0] Wgt_3_272,
input [18:0] Wgt_3_273,
input [18:0] Wgt_3_274,
input [18:0] Wgt_3_275,
input [18:0] Wgt_3_276,
input [18:0] Wgt_3_277,
input [18:0] Wgt_3_278,
input [18:0] Wgt_3_279,
input [18:0] Wgt_3_280,
input [18:0] Wgt_3_281,
input [18:0] Wgt_3_282,
input [18:0] Wgt_3_283,
input [18:0] Wgt_3_284,
input [18:0] Wgt_3_285,
input [18:0] Wgt_3_286,
input [18:0] Wgt_3_287,
input [18:0] Wgt_3_288,
input [18:0] Wgt_3_289,
input [18:0] Wgt_3_290,
input [18:0] Wgt_3_291,
input [18:0] Wgt_3_292,
input [18:0] Wgt_3_293,
input [18:0] Wgt_3_294,
input [18:0] Wgt_3_295,
input [18:0] Wgt_3_296,
input [18:0] Wgt_3_297,
input [18:0] Wgt_3_298,
input [18:0] Wgt_3_299,
input [18:0] Wgt_3_300,
input [18:0] Wgt_3_301,
input [18:0] Wgt_3_302,
input [18:0] Wgt_3_303,
input [18:0] Wgt_3_304,
input [18:0] Wgt_3_305,
input [18:0] Wgt_3_306,
input [18:0] Wgt_3_307,
input [18:0] Wgt_3_308,
input [18:0] Wgt_3_309,
input [18:0] Wgt_3_310,
input [18:0] Wgt_3_311,
input [18:0] Wgt_3_312,
input [18:0] Wgt_3_313,
input [18:0] Wgt_3_314,
input [18:0] Wgt_3_315,
input [18:0] Wgt_3_316,
input [18:0] Wgt_3_317,
input [18:0] Wgt_3_318,
input [18:0] Wgt_3_319,
input [18:0] Wgt_3_320,
input [18:0] Wgt_3_321,
input [18:0] Wgt_3_322,
input [18:0] Wgt_3_323,
input [18:0] Wgt_3_324,
input [18:0] Wgt_3_325,
input [18:0] Wgt_3_326,
input [18:0] Wgt_3_327,
input [18:0] Wgt_3_328,
input [18:0] Wgt_3_329,
input [18:0] Wgt_3_330,
input [18:0] Wgt_3_331,
input [18:0] Wgt_3_332,
input [18:0] Wgt_3_333,
input [18:0] Wgt_3_334,
input [18:0] Wgt_3_335,
input [18:0] Wgt_3_336,
input [18:0] Wgt_3_337,
input [18:0] Wgt_3_338,
input [18:0] Wgt_3_339,
input [18:0] Wgt_3_340,
input [18:0] Wgt_3_341,
input [18:0] Wgt_3_342,
input [18:0] Wgt_3_343,
input [18:0] Wgt_3_344,
input [18:0] Wgt_3_345,
input [18:0] Wgt_3_346,
input [18:0] Wgt_3_347,
input [18:0] Wgt_3_348,
input [18:0] Wgt_3_349,
input [18:0] Wgt_3_350,
input [18:0] Wgt_3_351,
input [18:0] Wgt_3_352,
input [18:0] Wgt_3_353,
input [18:0] Wgt_3_354,
input [18:0] Wgt_3_355,
input [18:0] Wgt_3_356,
input [18:0] Wgt_3_357,
input [18:0] Wgt_3_358,
input [18:0] Wgt_3_359,
input [18:0] Wgt_3_360,
input [18:0] Wgt_3_361,
input [18:0] Wgt_3_362,
input [18:0] Wgt_3_363,
input [18:0] Wgt_3_364,
input [18:0] Wgt_3_365,
input [18:0] Wgt_3_366,
input [18:0] Wgt_3_367,
input [18:0] Wgt_3_368,
input [18:0] Wgt_3_369,
input [18:0] Wgt_3_370,
input [18:0] Wgt_3_371,
input [18:0] Wgt_3_372,
input [18:0] Wgt_3_373,
input [18:0] Wgt_3_374,
input [18:0] Wgt_3_375,
input [18:0] Wgt_3_376,
input [18:0] Wgt_3_377,
input [18:0] Wgt_3_378,
input [18:0] Wgt_3_379,
input [18:0] Wgt_3_380,
input [18:0] Wgt_3_381,
input [18:0] Wgt_3_382,
input [18:0] Wgt_3_383,
input [18:0] Wgt_3_384,
input [18:0] Wgt_3_385,
input [18:0] Wgt_3_386,
input [18:0] Wgt_3_387,
input [18:0] Wgt_3_388,
input [18:0] Wgt_3_389,
input [18:0] Wgt_3_390,
input [18:0] Wgt_3_391,
input [18:0] Wgt_3_392,
input [18:0] Wgt_3_393,
input [18:0] Wgt_3_394,
input [18:0] Wgt_3_395,
input [18:0] Wgt_3_396,
input [18:0] Wgt_3_397,
input [18:0] Wgt_3_398,
input [18:0] Wgt_3_399,
input [18:0] Wgt_3_400,
input [18:0] Wgt_3_401,
input [18:0] Wgt_3_402,
input [18:0] Wgt_3_403,
input [18:0] Wgt_3_404,
input [18:0] Wgt_3_405,
input [18:0] Wgt_3_406,
input [18:0] Wgt_3_407,
input [18:0] Wgt_3_408,
input [18:0] Wgt_3_409,
input [18:0] Wgt_3_410,
input [18:0] Wgt_3_411,
input [18:0] Wgt_3_412,
input [18:0] Wgt_3_413,
input [18:0] Wgt_3_414,
input [18:0] Wgt_3_415,
input [18:0] Wgt_3_416,
input [18:0] Wgt_3_417,
input [18:0] Wgt_3_418,
input [18:0] Wgt_3_419,
input [18:0] Wgt_3_420,
input [18:0] Wgt_3_421,
input [18:0] Wgt_3_422,
input [18:0] Wgt_3_423,
input [18:0] Wgt_3_424,
input [18:0] Wgt_3_425,
input [18:0] Wgt_3_426,
input [18:0] Wgt_3_427,
input [18:0] Wgt_3_428,
input [18:0] Wgt_3_429,
input [18:0] Wgt_3_430,
input [18:0] Wgt_3_431,
input [18:0] Wgt_3_432,
input [18:0] Wgt_3_433,
input [18:0] Wgt_3_434,
input [18:0] Wgt_3_435,
input [18:0] Wgt_3_436,
input [18:0] Wgt_3_437,
input [18:0] Wgt_3_438,
input [18:0] Wgt_3_439,
input [18:0] Wgt_3_440,
input [18:0] Wgt_3_441,
input [18:0] Wgt_3_442,
input [18:0] Wgt_3_443,
input [18:0] Wgt_3_444,
input [18:0] Wgt_3_445,
input [18:0] Wgt_3_446,
input [18:0] Wgt_3_447,
input [18:0] Wgt_3_448,
input [18:0] Wgt_3_449,
input [18:0] Wgt_3_450,
input [18:0] Wgt_3_451,
input [18:0] Wgt_3_452,
input [18:0] Wgt_3_453,
input [18:0] Wgt_3_454,
input [18:0] Wgt_3_455,
input [18:0] Wgt_3_456,
input [18:0] Wgt_3_457,
input [18:0] Wgt_3_458,
input [18:0] Wgt_3_459,
input [18:0] Wgt_3_460,
input [18:0] Wgt_3_461,
input [18:0] Wgt_3_462,
input [18:0] Wgt_3_463,
input [18:0] Wgt_3_464,
input [18:0] Wgt_3_465,
input [18:0] Wgt_3_466,
input [18:0] Wgt_3_467,
input [18:0] Wgt_3_468,
input [18:0] Wgt_3_469,
input [18:0] Wgt_3_470,
input [18:0] Wgt_3_471,
input [18:0] Wgt_3_472,
input [18:0] Wgt_3_473,
input [18:0] Wgt_3_474,
input [18:0] Wgt_3_475,
input [18:0] Wgt_3_476,
input [18:0] Wgt_3_477,
input [18:0] Wgt_3_478,
input [18:0] Wgt_3_479,
input [18:0] Wgt_3_480,
input [18:0] Wgt_3_481,
input [18:0] Wgt_3_482,
input [18:0] Wgt_3_483,
input [18:0] Wgt_3_484,
input [18:0] Wgt_3_485,
input [18:0] Wgt_3_486,
input [18:0] Wgt_3_487,
input [18:0] Wgt_3_488,
input [18:0] Wgt_3_489,
input [18:0] Wgt_3_490,
input [18:0] Wgt_3_491,
input [18:0] Wgt_3_492,
input [18:0] Wgt_3_493,
input [18:0] Wgt_3_494,
input [18:0] Wgt_3_495,
input [18:0] Wgt_3_496,
input [18:0] Wgt_3_497,
input [18:0] Wgt_3_498,
input [18:0] Wgt_3_499,
input [18:0] Wgt_3_500,
input [18:0] Wgt_3_501,
input [18:0] Wgt_3_502,
input [18:0] Wgt_3_503,
input [18:0] Wgt_3_504,
input [18:0] Wgt_3_505,
input [18:0] Wgt_3_506,
input [18:0] Wgt_3_507,
input [18:0] Wgt_3_508,
input [18:0] Wgt_3_509,
input [18:0] Wgt_3_510,
input [18:0] Wgt_3_511,
input [18:0] Wgt_3_512,
input [18:0] Wgt_3_513,
input [18:0] Wgt_3_514,
input [18:0] Wgt_3_515,
input [18:0] Wgt_3_516,
input [18:0] Wgt_3_517,
input [18:0] Wgt_3_518,
input [18:0] Wgt_3_519,
input [18:0] Wgt_3_520,
input [18:0] Wgt_3_521,
input [18:0] Wgt_3_522,
input [18:0] Wgt_3_523,
input [18:0] Wgt_3_524,
input [18:0] Wgt_3_525,
input [18:0] Wgt_3_526,
input [18:0] Wgt_3_527,
input [18:0] Wgt_3_528,
input [18:0] Wgt_3_529,
input [18:0] Wgt_3_530,
input [18:0] Wgt_3_531,
input [18:0] Wgt_3_532,
input [18:0] Wgt_3_533,
input [18:0] Wgt_3_534,
input [18:0] Wgt_3_535,
input [18:0] Wgt_3_536,
input [18:0] Wgt_3_537,
input [18:0] Wgt_3_538,
input [18:0] Wgt_3_539,
input [18:0] Wgt_3_540,
input [18:0] Wgt_3_541,
input [18:0] Wgt_3_542,
input [18:0] Wgt_3_543,
input [18:0] Wgt_3_544,
input [18:0] Wgt_3_545,
input [18:0] Wgt_3_546,
input [18:0] Wgt_3_547,
input [18:0] Wgt_3_548,
input [18:0] Wgt_3_549,
input [18:0] Wgt_3_550,
input [18:0] Wgt_3_551,
input [18:0] Wgt_3_552,
input [18:0] Wgt_3_553,
input [18:0] Wgt_3_554,
input [18:0] Wgt_3_555,
input [18:0] Wgt_3_556,
input [18:0] Wgt_3_557,
input [18:0] Wgt_3_558,
input [18:0] Wgt_3_559,
input [18:0] Wgt_3_560,
input [18:0] Wgt_3_561,
input [18:0] Wgt_3_562,
input [18:0] Wgt_3_563,
input [18:0] Wgt_3_564,
input [18:0] Wgt_3_565,
input [18:0] Wgt_3_566,
input [18:0] Wgt_3_567,
input [18:0] Wgt_3_568,
input [18:0] Wgt_3_569,
input [18:0] Wgt_3_570,
input [18:0] Wgt_3_571,
input [18:0] Wgt_3_572,
input [18:0] Wgt_3_573,
input [18:0] Wgt_3_574,
input [18:0] Wgt_3_575,
input [18:0] Wgt_3_576,
input [18:0] Wgt_3_577,
input [18:0] Wgt_3_578,
input [18:0] Wgt_3_579,
input [18:0] Wgt_3_580,
input [18:0] Wgt_3_581,
input [18:0] Wgt_3_582,
input [18:0] Wgt_3_583,
input [18:0] Wgt_3_584,
input [18:0] Wgt_3_585,
input [18:0] Wgt_3_586,
input [18:0] Wgt_3_587,
input [18:0] Wgt_3_588,
input [18:0] Wgt_3_589,
input [18:0] Wgt_3_590,
input [18:0] Wgt_3_591,
input [18:0] Wgt_3_592,
input [18:0] Wgt_3_593,
input [18:0] Wgt_3_594,
input [18:0] Wgt_3_595,
input [18:0] Wgt_3_596,
input [18:0] Wgt_3_597,
input [18:0] Wgt_3_598,
input [18:0] Wgt_3_599,
input [18:0] Wgt_3_600,
input [18:0] Wgt_3_601,
input [18:0] Wgt_3_602,
input [18:0] Wgt_3_603,
input [18:0] Wgt_3_604,
input [18:0] Wgt_3_605,
input [18:0] Wgt_3_606,
input [18:0] Wgt_3_607,
input [18:0] Wgt_3_608,
input [18:0] Wgt_3_609,
input [18:0] Wgt_3_610,
input [18:0] Wgt_3_611,
input [18:0] Wgt_3_612,
input [18:0] Wgt_3_613,
input [18:0] Wgt_3_614,
input [18:0] Wgt_3_615,
input [18:0] Wgt_3_616,
input [18:0] Wgt_3_617,
input [18:0] Wgt_3_618,
input [18:0] Wgt_3_619,
input [18:0] Wgt_3_620,
input [18:0] Wgt_3_621,
input [18:0] Wgt_3_622,
input [18:0] Wgt_3_623,
input [18:0] Wgt_3_624,
input [18:0] Wgt_3_625,
input [18:0] Wgt_3_626,
input [18:0] Wgt_3_627,
input [18:0] Wgt_3_628,
input [18:0] Wgt_3_629,
input [18:0] Wgt_3_630,
input [18:0] Wgt_3_631,
input [18:0] Wgt_3_632,
input [18:0] Wgt_3_633,
input [18:0] Wgt_3_634,
input [18:0] Wgt_3_635,
input [18:0] Wgt_3_636,
input [18:0] Wgt_3_637,
input [18:0] Wgt_3_638,
input [18:0] Wgt_3_639,
input [18:0] Wgt_3_640,
input [18:0] Wgt_3_641,
input [18:0] Wgt_3_642,
input [18:0] Wgt_3_643,
input [18:0] Wgt_3_644,
input [18:0] Wgt_3_645,
input [18:0] Wgt_3_646,
input [18:0] Wgt_3_647,
input [18:0] Wgt_3_648,
input [18:0] Wgt_3_649,
input [18:0] Wgt_3_650,
input [18:0] Wgt_3_651,
input [18:0] Wgt_3_652,
input [18:0] Wgt_3_653,
input [18:0] Wgt_3_654,
input [18:0] Wgt_3_655,
input [18:0] Wgt_3_656,
input [18:0] Wgt_3_657,
input [18:0] Wgt_3_658,
input [18:0] Wgt_3_659,
input [18:0] Wgt_3_660,
input [18:0] Wgt_3_661,
input [18:0] Wgt_3_662,
input [18:0] Wgt_3_663,
input [18:0] Wgt_3_664,
input [18:0] Wgt_3_665,
input [18:0] Wgt_3_666,
input [18:0] Wgt_3_667,
input [18:0] Wgt_3_668,
input [18:0] Wgt_3_669,
input [18:0] Wgt_3_670,
input [18:0] Wgt_3_671,
input [18:0] Wgt_3_672,
input [18:0] Wgt_3_673,
input [18:0] Wgt_3_674,
input [18:0] Wgt_3_675,
input [18:0] Wgt_3_676,
input [18:0] Wgt_3_677,
input [18:0] Wgt_3_678,
input [18:0] Wgt_3_679,
input [18:0] Wgt_3_680,
input [18:0] Wgt_3_681,
input [18:0] Wgt_3_682,
input [18:0] Wgt_3_683,
input [18:0] Wgt_3_684,
input [18:0] Wgt_3_685,
input [18:0] Wgt_3_686,
input [18:0] Wgt_3_687,
input [18:0] Wgt_3_688,
input [18:0] Wgt_3_689,
input [18:0] Wgt_3_690,
input [18:0] Wgt_3_691,
input [18:0] Wgt_3_692,
input [18:0] Wgt_3_693,
input [18:0] Wgt_3_694,
input [18:0] Wgt_3_695,
input [18:0] Wgt_3_696,
input [18:0] Wgt_3_697,
input [18:0] Wgt_3_698,
input [18:0] Wgt_3_699,
input [18:0] Wgt_3_700,
input [18:0] Wgt_3_701,
input [18:0] Wgt_3_702,
input [18:0] Wgt_3_703,
input [18:0] Wgt_3_704,
input [18:0] Wgt_3_705,
input [18:0] Wgt_3_706,
input [18:0] Wgt_3_707,
input [18:0] Wgt_3_708,
input [18:0] Wgt_3_709,
input [18:0] Wgt_3_710,
input [18:0] Wgt_3_711,
input [18:0] Wgt_3_712,
input [18:0] Wgt_3_713,
input [18:0] Wgt_3_714,
input [18:0] Wgt_3_715,
input [18:0] Wgt_3_716,
input [18:0] Wgt_3_717,
input [18:0] Wgt_3_718,
input [18:0] Wgt_3_719,
input [18:0] Wgt_3_720,
input [18:0] Wgt_3_721,
input [18:0] Wgt_3_722,
input [18:0] Wgt_3_723,
input [18:0] Wgt_3_724,
input [18:0] Wgt_3_725,
input [18:0] Wgt_3_726,
input [18:0] Wgt_3_727,
input [18:0] Wgt_3_728,
input [18:0] Wgt_3_729,
input [18:0] Wgt_3_730,
input [18:0] Wgt_3_731,
input [18:0] Wgt_3_732,
input [18:0] Wgt_3_733,
input [18:0] Wgt_3_734,
input [18:0] Wgt_3_735,
input [18:0] Wgt_3_736,
input [18:0] Wgt_3_737,
input [18:0] Wgt_3_738,
input [18:0] Wgt_3_739,
input [18:0] Wgt_3_740,
input [18:0] Wgt_3_741,
input [18:0] Wgt_3_742,
input [18:0] Wgt_3_743,
input [18:0] Wgt_3_744,
input [18:0] Wgt_3_745,
input [18:0] Wgt_3_746,
input [18:0] Wgt_3_747,
input [18:0] Wgt_3_748,
input [18:0] Wgt_3_749,
input [18:0] Wgt_3_750,
input [18:0] Wgt_3_751,
input [18:0] Wgt_3_752,
input [18:0] Wgt_3_753,
input [18:0] Wgt_3_754,
input [18:0] Wgt_3_755,
input [18:0] Wgt_3_756,
input [18:0] Wgt_3_757,
input [18:0] Wgt_3_758,
input [18:0] Wgt_3_759,
input [18:0] Wgt_3_760,
input [18:0] Wgt_3_761,
input [18:0] Wgt_3_762,
input [18:0] Wgt_3_763,
input [18:0] Wgt_3_764,
input [18:0] Wgt_3_765,
input [18:0] Wgt_3_766,
input [18:0] Wgt_3_767,
input [18:0] Wgt_3_768,
input [18:0] Wgt_3_769,
input [18:0] Wgt_3_770,
input [18:0] Wgt_3_771,
input [18:0] Wgt_3_772,
input [18:0] Wgt_3_773,
input [18:0] Wgt_3_774,
input [18:0] Wgt_3_775,
input [18:0] Wgt_3_776,
input [18:0] Wgt_3_777,
input [18:0] Wgt_3_778,
input [18:0] Wgt_3_779,
input [18:0] Wgt_3_780,
input [18:0] Wgt_3_781,
input [18:0] Wgt_3_782,
input [18:0] Wgt_3_783,
input [18:0] Wgt_3_784,
input [18:0] Wgt_4_0,
input [18:0] Wgt_4_1,
input [18:0] Wgt_4_2,
input [18:0] Wgt_4_3,
input [18:0] Wgt_4_4,
input [18:0] Wgt_4_5,
input [18:0] Wgt_4_6,
input [18:0] Wgt_4_7,
input [18:0] Wgt_4_8,
input [18:0] Wgt_4_9,
input [18:0] Wgt_4_10,
input [18:0] Wgt_4_11,
input [18:0] Wgt_4_12,
input [18:0] Wgt_4_13,
input [18:0] Wgt_4_14,
input [18:0] Wgt_4_15,
input [18:0] Wgt_4_16,
input [18:0] Wgt_4_17,
input [18:0] Wgt_4_18,
input [18:0] Wgt_4_19,
input [18:0] Wgt_4_20,
input [18:0] Wgt_4_21,
input [18:0] Wgt_4_22,
input [18:0] Wgt_4_23,
input [18:0] Wgt_4_24,
input [18:0] Wgt_4_25,
input [18:0] Wgt_4_26,
input [18:0] Wgt_4_27,
input [18:0] Wgt_4_28,
input [18:0] Wgt_4_29,
input [18:0] Wgt_4_30,
input [18:0] Wgt_4_31,
input [18:0] Wgt_4_32,
input [18:0] Wgt_4_33,
input [18:0] Wgt_4_34,
input [18:0] Wgt_4_35,
input [18:0] Wgt_4_36,
input [18:0] Wgt_4_37,
input [18:0] Wgt_4_38,
input [18:0] Wgt_4_39,
input [18:0] Wgt_4_40,
input [18:0] Wgt_4_41,
input [18:0] Wgt_4_42,
input [18:0] Wgt_4_43,
input [18:0] Wgt_4_44,
input [18:0] Wgt_4_45,
input [18:0] Wgt_4_46,
input [18:0] Wgt_4_47,
input [18:0] Wgt_4_48,
input [18:0] Wgt_4_49,
input [18:0] Wgt_4_50,
input [18:0] Wgt_4_51,
input [18:0] Wgt_4_52,
input [18:0] Wgt_4_53,
input [18:0] Wgt_4_54,
input [18:0] Wgt_4_55,
input [18:0] Wgt_4_56,
input [18:0] Wgt_4_57,
input [18:0] Wgt_4_58,
input [18:0] Wgt_4_59,
input [18:0] Wgt_4_60,
input [18:0] Wgt_4_61,
input [18:0] Wgt_4_62,
input [18:0] Wgt_4_63,
input [18:0] Wgt_4_64,
input [18:0] Wgt_4_65,
input [18:0] Wgt_4_66,
input [18:0] Wgt_4_67,
input [18:0] Wgt_4_68,
input [18:0] Wgt_4_69,
input [18:0] Wgt_4_70,
input [18:0] Wgt_4_71,
input [18:0] Wgt_4_72,
input [18:0] Wgt_4_73,
input [18:0] Wgt_4_74,
input [18:0] Wgt_4_75,
input [18:0] Wgt_4_76,
input [18:0] Wgt_4_77,
input [18:0] Wgt_4_78,
input [18:0] Wgt_4_79,
input [18:0] Wgt_4_80,
input [18:0] Wgt_4_81,
input [18:0] Wgt_4_82,
input [18:0] Wgt_4_83,
input [18:0] Wgt_4_84,
input [18:0] Wgt_4_85,
input [18:0] Wgt_4_86,
input [18:0] Wgt_4_87,
input [18:0] Wgt_4_88,
input [18:0] Wgt_4_89,
input [18:0] Wgt_4_90,
input [18:0] Wgt_4_91,
input [18:0] Wgt_4_92,
input [18:0] Wgt_4_93,
input [18:0] Wgt_4_94,
input [18:0] Wgt_4_95,
input [18:0] Wgt_4_96,
input [18:0] Wgt_4_97,
input [18:0] Wgt_4_98,
input [18:0] Wgt_4_99,
input [18:0] Wgt_4_100,
input [18:0] Wgt_4_101,
input [18:0] Wgt_4_102,
input [18:0] Wgt_4_103,
input [18:0] Wgt_4_104,
input [18:0] Wgt_4_105,
input [18:0] Wgt_4_106,
input [18:0] Wgt_4_107,
input [18:0] Wgt_4_108,
input [18:0] Wgt_4_109,
input [18:0] Wgt_4_110,
input [18:0] Wgt_4_111,
input [18:0] Wgt_4_112,
input [18:0] Wgt_4_113,
input [18:0] Wgt_4_114,
input [18:0] Wgt_4_115,
input [18:0] Wgt_4_116,
input [18:0] Wgt_4_117,
input [18:0] Wgt_4_118,
input [18:0] Wgt_4_119,
input [18:0] Wgt_4_120,
input [18:0] Wgt_4_121,
input [18:0] Wgt_4_122,
input [18:0] Wgt_4_123,
input [18:0] Wgt_4_124,
input [18:0] Wgt_4_125,
input [18:0] Wgt_4_126,
input [18:0] Wgt_4_127,
input [18:0] Wgt_4_128,
input [18:0] Wgt_4_129,
input [18:0] Wgt_4_130,
input [18:0] Wgt_4_131,
input [18:0] Wgt_4_132,
input [18:0] Wgt_4_133,
input [18:0] Wgt_4_134,
input [18:0] Wgt_4_135,
input [18:0] Wgt_4_136,
input [18:0] Wgt_4_137,
input [18:0] Wgt_4_138,
input [18:0] Wgt_4_139,
input [18:0] Wgt_4_140,
input [18:0] Wgt_4_141,
input [18:0] Wgt_4_142,
input [18:0] Wgt_4_143,
input [18:0] Wgt_4_144,
input [18:0] Wgt_4_145,
input [18:0] Wgt_4_146,
input [18:0] Wgt_4_147,
input [18:0] Wgt_4_148,
input [18:0] Wgt_4_149,
input [18:0] Wgt_4_150,
input [18:0] Wgt_4_151,
input [18:0] Wgt_4_152,
input [18:0] Wgt_4_153,
input [18:0] Wgt_4_154,
input [18:0] Wgt_4_155,
input [18:0] Wgt_4_156,
input [18:0] Wgt_4_157,
input [18:0] Wgt_4_158,
input [18:0] Wgt_4_159,
input [18:0] Wgt_4_160,
input [18:0] Wgt_4_161,
input [18:0] Wgt_4_162,
input [18:0] Wgt_4_163,
input [18:0] Wgt_4_164,
input [18:0] Wgt_4_165,
input [18:0] Wgt_4_166,
input [18:0] Wgt_4_167,
input [18:0] Wgt_4_168,
input [18:0] Wgt_4_169,
input [18:0] Wgt_4_170,
input [18:0] Wgt_4_171,
input [18:0] Wgt_4_172,
input [18:0] Wgt_4_173,
input [18:0] Wgt_4_174,
input [18:0] Wgt_4_175,
input [18:0] Wgt_4_176,
input [18:0] Wgt_4_177,
input [18:0] Wgt_4_178,
input [18:0] Wgt_4_179,
input [18:0] Wgt_4_180,
input [18:0] Wgt_4_181,
input [18:0] Wgt_4_182,
input [18:0] Wgt_4_183,
input [18:0] Wgt_4_184,
input [18:0] Wgt_4_185,
input [18:0] Wgt_4_186,
input [18:0] Wgt_4_187,
input [18:0] Wgt_4_188,
input [18:0] Wgt_4_189,
input [18:0] Wgt_4_190,
input [18:0] Wgt_4_191,
input [18:0] Wgt_4_192,
input [18:0] Wgt_4_193,
input [18:0] Wgt_4_194,
input [18:0] Wgt_4_195,
input [18:0] Wgt_4_196,
input [18:0] Wgt_4_197,
input [18:0] Wgt_4_198,
input [18:0] Wgt_4_199,
input [18:0] Wgt_4_200,
input [18:0] Wgt_4_201,
input [18:0] Wgt_4_202,
input [18:0] Wgt_4_203,
input [18:0] Wgt_4_204,
input [18:0] Wgt_4_205,
input [18:0] Wgt_4_206,
input [18:0] Wgt_4_207,
input [18:0] Wgt_4_208,
input [18:0] Wgt_4_209,
input [18:0] Wgt_4_210,
input [18:0] Wgt_4_211,
input [18:0] Wgt_4_212,
input [18:0] Wgt_4_213,
input [18:0] Wgt_4_214,
input [18:0] Wgt_4_215,
input [18:0] Wgt_4_216,
input [18:0] Wgt_4_217,
input [18:0] Wgt_4_218,
input [18:0] Wgt_4_219,
input [18:0] Wgt_4_220,
input [18:0] Wgt_4_221,
input [18:0] Wgt_4_222,
input [18:0] Wgt_4_223,
input [18:0] Wgt_4_224,
input [18:0] Wgt_4_225,
input [18:0] Wgt_4_226,
input [18:0] Wgt_4_227,
input [18:0] Wgt_4_228,
input [18:0] Wgt_4_229,
input [18:0] Wgt_4_230,
input [18:0] Wgt_4_231,
input [18:0] Wgt_4_232,
input [18:0] Wgt_4_233,
input [18:0] Wgt_4_234,
input [18:0] Wgt_4_235,
input [18:0] Wgt_4_236,
input [18:0] Wgt_4_237,
input [18:0] Wgt_4_238,
input [18:0] Wgt_4_239,
input [18:0] Wgt_4_240,
input [18:0] Wgt_4_241,
input [18:0] Wgt_4_242,
input [18:0] Wgt_4_243,
input [18:0] Wgt_4_244,
input [18:0] Wgt_4_245,
input [18:0] Wgt_4_246,
input [18:0] Wgt_4_247,
input [18:0] Wgt_4_248,
input [18:0] Wgt_4_249,
input [18:0] Wgt_4_250,
input [18:0] Wgt_4_251,
input [18:0] Wgt_4_252,
input [18:0] Wgt_4_253,
input [18:0] Wgt_4_254,
input [18:0] Wgt_4_255,
input [18:0] Wgt_4_256,
input [18:0] Wgt_4_257,
input [18:0] Wgt_4_258,
input [18:0] Wgt_4_259,
input [18:0] Wgt_4_260,
input [18:0] Wgt_4_261,
input [18:0] Wgt_4_262,
input [18:0] Wgt_4_263,
input [18:0] Wgt_4_264,
input [18:0] Wgt_4_265,
input [18:0] Wgt_4_266,
input [18:0] Wgt_4_267,
input [18:0] Wgt_4_268,
input [18:0] Wgt_4_269,
input [18:0] Wgt_4_270,
input [18:0] Wgt_4_271,
input [18:0] Wgt_4_272,
input [18:0] Wgt_4_273,
input [18:0] Wgt_4_274,
input [18:0] Wgt_4_275,
input [18:0] Wgt_4_276,
input [18:0] Wgt_4_277,
input [18:0] Wgt_4_278,
input [18:0] Wgt_4_279,
input [18:0] Wgt_4_280,
input [18:0] Wgt_4_281,
input [18:0] Wgt_4_282,
input [18:0] Wgt_4_283,
input [18:0] Wgt_4_284,
input [18:0] Wgt_4_285,
input [18:0] Wgt_4_286,
input [18:0] Wgt_4_287,
input [18:0] Wgt_4_288,
input [18:0] Wgt_4_289,
input [18:0] Wgt_4_290,
input [18:0] Wgt_4_291,
input [18:0] Wgt_4_292,
input [18:0] Wgt_4_293,
input [18:0] Wgt_4_294,
input [18:0] Wgt_4_295,
input [18:0] Wgt_4_296,
input [18:0] Wgt_4_297,
input [18:0] Wgt_4_298,
input [18:0] Wgt_4_299,
input [18:0] Wgt_4_300,
input [18:0] Wgt_4_301,
input [18:0] Wgt_4_302,
input [18:0] Wgt_4_303,
input [18:0] Wgt_4_304,
input [18:0] Wgt_4_305,
input [18:0] Wgt_4_306,
input [18:0] Wgt_4_307,
input [18:0] Wgt_4_308,
input [18:0] Wgt_4_309,
input [18:0] Wgt_4_310,
input [18:0] Wgt_4_311,
input [18:0] Wgt_4_312,
input [18:0] Wgt_4_313,
input [18:0] Wgt_4_314,
input [18:0] Wgt_4_315,
input [18:0] Wgt_4_316,
input [18:0] Wgt_4_317,
input [18:0] Wgt_4_318,
input [18:0] Wgt_4_319,
input [18:0] Wgt_4_320,
input [18:0] Wgt_4_321,
input [18:0] Wgt_4_322,
input [18:0] Wgt_4_323,
input [18:0] Wgt_4_324,
input [18:0] Wgt_4_325,
input [18:0] Wgt_4_326,
input [18:0] Wgt_4_327,
input [18:0] Wgt_4_328,
input [18:0] Wgt_4_329,
input [18:0] Wgt_4_330,
input [18:0] Wgt_4_331,
input [18:0] Wgt_4_332,
input [18:0] Wgt_4_333,
input [18:0] Wgt_4_334,
input [18:0] Wgt_4_335,
input [18:0] Wgt_4_336,
input [18:0] Wgt_4_337,
input [18:0] Wgt_4_338,
input [18:0] Wgt_4_339,
input [18:0] Wgt_4_340,
input [18:0] Wgt_4_341,
input [18:0] Wgt_4_342,
input [18:0] Wgt_4_343,
input [18:0] Wgt_4_344,
input [18:0] Wgt_4_345,
input [18:0] Wgt_4_346,
input [18:0] Wgt_4_347,
input [18:0] Wgt_4_348,
input [18:0] Wgt_4_349,
input [18:0] Wgt_4_350,
input [18:0] Wgt_4_351,
input [18:0] Wgt_4_352,
input [18:0] Wgt_4_353,
input [18:0] Wgt_4_354,
input [18:0] Wgt_4_355,
input [18:0] Wgt_4_356,
input [18:0] Wgt_4_357,
input [18:0] Wgt_4_358,
input [18:0] Wgt_4_359,
input [18:0] Wgt_4_360,
input [18:0] Wgt_4_361,
input [18:0] Wgt_4_362,
input [18:0] Wgt_4_363,
input [18:0] Wgt_4_364,
input [18:0] Wgt_4_365,
input [18:0] Wgt_4_366,
input [18:0] Wgt_4_367,
input [18:0] Wgt_4_368,
input [18:0] Wgt_4_369,
input [18:0] Wgt_4_370,
input [18:0] Wgt_4_371,
input [18:0] Wgt_4_372,
input [18:0] Wgt_4_373,
input [18:0] Wgt_4_374,
input [18:0] Wgt_4_375,
input [18:0] Wgt_4_376,
input [18:0] Wgt_4_377,
input [18:0] Wgt_4_378,
input [18:0] Wgt_4_379,
input [18:0] Wgt_4_380,
input [18:0] Wgt_4_381,
input [18:0] Wgt_4_382,
input [18:0] Wgt_4_383,
input [18:0] Wgt_4_384,
input [18:0] Wgt_4_385,
input [18:0] Wgt_4_386,
input [18:0] Wgt_4_387,
input [18:0] Wgt_4_388,
input [18:0] Wgt_4_389,
input [18:0] Wgt_4_390,
input [18:0] Wgt_4_391,
input [18:0] Wgt_4_392,
input [18:0] Wgt_4_393,
input [18:0] Wgt_4_394,
input [18:0] Wgt_4_395,
input [18:0] Wgt_4_396,
input [18:0] Wgt_4_397,
input [18:0] Wgt_4_398,
input [18:0] Wgt_4_399,
input [18:0] Wgt_4_400,
input [18:0] Wgt_4_401,
input [18:0] Wgt_4_402,
input [18:0] Wgt_4_403,
input [18:0] Wgt_4_404,
input [18:0] Wgt_4_405,
input [18:0] Wgt_4_406,
input [18:0] Wgt_4_407,
input [18:0] Wgt_4_408,
input [18:0] Wgt_4_409,
input [18:0] Wgt_4_410,
input [18:0] Wgt_4_411,
input [18:0] Wgt_4_412,
input [18:0] Wgt_4_413,
input [18:0] Wgt_4_414,
input [18:0] Wgt_4_415,
input [18:0] Wgt_4_416,
input [18:0] Wgt_4_417,
input [18:0] Wgt_4_418,
input [18:0] Wgt_4_419,
input [18:0] Wgt_4_420,
input [18:0] Wgt_4_421,
input [18:0] Wgt_4_422,
input [18:0] Wgt_4_423,
input [18:0] Wgt_4_424,
input [18:0] Wgt_4_425,
input [18:0] Wgt_4_426,
input [18:0] Wgt_4_427,
input [18:0] Wgt_4_428,
input [18:0] Wgt_4_429,
input [18:0] Wgt_4_430,
input [18:0] Wgt_4_431,
input [18:0] Wgt_4_432,
input [18:0] Wgt_4_433,
input [18:0] Wgt_4_434,
input [18:0] Wgt_4_435,
input [18:0] Wgt_4_436,
input [18:0] Wgt_4_437,
input [18:0] Wgt_4_438,
input [18:0] Wgt_4_439,
input [18:0] Wgt_4_440,
input [18:0] Wgt_4_441,
input [18:0] Wgt_4_442,
input [18:0] Wgt_4_443,
input [18:0] Wgt_4_444,
input [18:0] Wgt_4_445,
input [18:0] Wgt_4_446,
input [18:0] Wgt_4_447,
input [18:0] Wgt_4_448,
input [18:0] Wgt_4_449,
input [18:0] Wgt_4_450,
input [18:0] Wgt_4_451,
input [18:0] Wgt_4_452,
input [18:0] Wgt_4_453,
input [18:0] Wgt_4_454,
input [18:0] Wgt_4_455,
input [18:0] Wgt_4_456,
input [18:0] Wgt_4_457,
input [18:0] Wgt_4_458,
input [18:0] Wgt_4_459,
input [18:0] Wgt_4_460,
input [18:0] Wgt_4_461,
input [18:0] Wgt_4_462,
input [18:0] Wgt_4_463,
input [18:0] Wgt_4_464,
input [18:0] Wgt_4_465,
input [18:0] Wgt_4_466,
input [18:0] Wgt_4_467,
input [18:0] Wgt_4_468,
input [18:0] Wgt_4_469,
input [18:0] Wgt_4_470,
input [18:0] Wgt_4_471,
input [18:0] Wgt_4_472,
input [18:0] Wgt_4_473,
input [18:0] Wgt_4_474,
input [18:0] Wgt_4_475,
input [18:0] Wgt_4_476,
input [18:0] Wgt_4_477,
input [18:0] Wgt_4_478,
input [18:0] Wgt_4_479,
input [18:0] Wgt_4_480,
input [18:0] Wgt_4_481,
input [18:0] Wgt_4_482,
input [18:0] Wgt_4_483,
input [18:0] Wgt_4_484,
input [18:0] Wgt_4_485,
input [18:0] Wgt_4_486,
input [18:0] Wgt_4_487,
input [18:0] Wgt_4_488,
input [18:0] Wgt_4_489,
input [18:0] Wgt_4_490,
input [18:0] Wgt_4_491,
input [18:0] Wgt_4_492,
input [18:0] Wgt_4_493,
input [18:0] Wgt_4_494,
input [18:0] Wgt_4_495,
input [18:0] Wgt_4_496,
input [18:0] Wgt_4_497,
input [18:0] Wgt_4_498,
input [18:0] Wgt_4_499,
input [18:0] Wgt_4_500,
input [18:0] Wgt_4_501,
input [18:0] Wgt_4_502,
input [18:0] Wgt_4_503,
input [18:0] Wgt_4_504,
input [18:0] Wgt_4_505,
input [18:0] Wgt_4_506,
input [18:0] Wgt_4_507,
input [18:0] Wgt_4_508,
input [18:0] Wgt_4_509,
input [18:0] Wgt_4_510,
input [18:0] Wgt_4_511,
input [18:0] Wgt_4_512,
input [18:0] Wgt_4_513,
input [18:0] Wgt_4_514,
input [18:0] Wgt_4_515,
input [18:0] Wgt_4_516,
input [18:0] Wgt_4_517,
input [18:0] Wgt_4_518,
input [18:0] Wgt_4_519,
input [18:0] Wgt_4_520,
input [18:0] Wgt_4_521,
input [18:0] Wgt_4_522,
input [18:0] Wgt_4_523,
input [18:0] Wgt_4_524,
input [18:0] Wgt_4_525,
input [18:0] Wgt_4_526,
input [18:0] Wgt_4_527,
input [18:0] Wgt_4_528,
input [18:0] Wgt_4_529,
input [18:0] Wgt_4_530,
input [18:0] Wgt_4_531,
input [18:0] Wgt_4_532,
input [18:0] Wgt_4_533,
input [18:0] Wgt_4_534,
input [18:0] Wgt_4_535,
input [18:0] Wgt_4_536,
input [18:0] Wgt_4_537,
input [18:0] Wgt_4_538,
input [18:0] Wgt_4_539,
input [18:0] Wgt_4_540,
input [18:0] Wgt_4_541,
input [18:0] Wgt_4_542,
input [18:0] Wgt_4_543,
input [18:0] Wgt_4_544,
input [18:0] Wgt_4_545,
input [18:0] Wgt_4_546,
input [18:0] Wgt_4_547,
input [18:0] Wgt_4_548,
input [18:0] Wgt_4_549,
input [18:0] Wgt_4_550,
input [18:0] Wgt_4_551,
input [18:0] Wgt_4_552,
input [18:0] Wgt_4_553,
input [18:0] Wgt_4_554,
input [18:0] Wgt_4_555,
input [18:0] Wgt_4_556,
input [18:0] Wgt_4_557,
input [18:0] Wgt_4_558,
input [18:0] Wgt_4_559,
input [18:0] Wgt_4_560,
input [18:0] Wgt_4_561,
input [18:0] Wgt_4_562,
input [18:0] Wgt_4_563,
input [18:0] Wgt_4_564,
input [18:0] Wgt_4_565,
input [18:0] Wgt_4_566,
input [18:0] Wgt_4_567,
input [18:0] Wgt_4_568,
input [18:0] Wgt_4_569,
input [18:0] Wgt_4_570,
input [18:0] Wgt_4_571,
input [18:0] Wgt_4_572,
input [18:0] Wgt_4_573,
input [18:0] Wgt_4_574,
input [18:0] Wgt_4_575,
input [18:0] Wgt_4_576,
input [18:0] Wgt_4_577,
input [18:0] Wgt_4_578,
input [18:0] Wgt_4_579,
input [18:0] Wgt_4_580,
input [18:0] Wgt_4_581,
input [18:0] Wgt_4_582,
input [18:0] Wgt_4_583,
input [18:0] Wgt_4_584,
input [18:0] Wgt_4_585,
input [18:0] Wgt_4_586,
input [18:0] Wgt_4_587,
input [18:0] Wgt_4_588,
input [18:0] Wgt_4_589,
input [18:0] Wgt_4_590,
input [18:0] Wgt_4_591,
input [18:0] Wgt_4_592,
input [18:0] Wgt_4_593,
input [18:0] Wgt_4_594,
input [18:0] Wgt_4_595,
input [18:0] Wgt_4_596,
input [18:0] Wgt_4_597,
input [18:0] Wgt_4_598,
input [18:0] Wgt_4_599,
input [18:0] Wgt_4_600,
input [18:0] Wgt_4_601,
input [18:0] Wgt_4_602,
input [18:0] Wgt_4_603,
input [18:0] Wgt_4_604,
input [18:0] Wgt_4_605,
input [18:0] Wgt_4_606,
input [18:0] Wgt_4_607,
input [18:0] Wgt_4_608,
input [18:0] Wgt_4_609,
input [18:0] Wgt_4_610,
input [18:0] Wgt_4_611,
input [18:0] Wgt_4_612,
input [18:0] Wgt_4_613,
input [18:0] Wgt_4_614,
input [18:0] Wgt_4_615,
input [18:0] Wgt_4_616,
input [18:0] Wgt_4_617,
input [18:0] Wgt_4_618,
input [18:0] Wgt_4_619,
input [18:0] Wgt_4_620,
input [18:0] Wgt_4_621,
input [18:0] Wgt_4_622,
input [18:0] Wgt_4_623,
input [18:0] Wgt_4_624,
input [18:0] Wgt_4_625,
input [18:0] Wgt_4_626,
input [18:0] Wgt_4_627,
input [18:0] Wgt_4_628,
input [18:0] Wgt_4_629,
input [18:0] Wgt_4_630,
input [18:0] Wgt_4_631,
input [18:0] Wgt_4_632,
input [18:0] Wgt_4_633,
input [18:0] Wgt_4_634,
input [18:0] Wgt_4_635,
input [18:0] Wgt_4_636,
input [18:0] Wgt_4_637,
input [18:0] Wgt_4_638,
input [18:0] Wgt_4_639,
input [18:0] Wgt_4_640,
input [18:0] Wgt_4_641,
input [18:0] Wgt_4_642,
input [18:0] Wgt_4_643,
input [18:0] Wgt_4_644,
input [18:0] Wgt_4_645,
input [18:0] Wgt_4_646,
input [18:0] Wgt_4_647,
input [18:0] Wgt_4_648,
input [18:0] Wgt_4_649,
input [18:0] Wgt_4_650,
input [18:0] Wgt_4_651,
input [18:0] Wgt_4_652,
input [18:0] Wgt_4_653,
input [18:0] Wgt_4_654,
input [18:0] Wgt_4_655,
input [18:0] Wgt_4_656,
input [18:0] Wgt_4_657,
input [18:0] Wgt_4_658,
input [18:0] Wgt_4_659,
input [18:0] Wgt_4_660,
input [18:0] Wgt_4_661,
input [18:0] Wgt_4_662,
input [18:0] Wgt_4_663,
input [18:0] Wgt_4_664,
input [18:0] Wgt_4_665,
input [18:0] Wgt_4_666,
input [18:0] Wgt_4_667,
input [18:0] Wgt_4_668,
input [18:0] Wgt_4_669,
input [18:0] Wgt_4_670,
input [18:0] Wgt_4_671,
input [18:0] Wgt_4_672,
input [18:0] Wgt_4_673,
input [18:0] Wgt_4_674,
input [18:0] Wgt_4_675,
input [18:0] Wgt_4_676,
input [18:0] Wgt_4_677,
input [18:0] Wgt_4_678,
input [18:0] Wgt_4_679,
input [18:0] Wgt_4_680,
input [18:0] Wgt_4_681,
input [18:0] Wgt_4_682,
input [18:0] Wgt_4_683,
input [18:0] Wgt_4_684,
input [18:0] Wgt_4_685,
input [18:0] Wgt_4_686,
input [18:0] Wgt_4_687,
input [18:0] Wgt_4_688,
input [18:0] Wgt_4_689,
input [18:0] Wgt_4_690,
input [18:0] Wgt_4_691,
input [18:0] Wgt_4_692,
input [18:0] Wgt_4_693,
input [18:0] Wgt_4_694,
input [18:0] Wgt_4_695,
input [18:0] Wgt_4_696,
input [18:0] Wgt_4_697,
input [18:0] Wgt_4_698,
input [18:0] Wgt_4_699,
input [18:0] Wgt_4_700,
input [18:0] Wgt_4_701,
input [18:0] Wgt_4_702,
input [18:0] Wgt_4_703,
input [18:0] Wgt_4_704,
input [18:0] Wgt_4_705,
input [18:0] Wgt_4_706,
input [18:0] Wgt_4_707,
input [18:0] Wgt_4_708,
input [18:0] Wgt_4_709,
input [18:0] Wgt_4_710,
input [18:0] Wgt_4_711,
input [18:0] Wgt_4_712,
input [18:0] Wgt_4_713,
input [18:0] Wgt_4_714,
input [18:0] Wgt_4_715,
input [18:0] Wgt_4_716,
input [18:0] Wgt_4_717,
input [18:0] Wgt_4_718,
input [18:0] Wgt_4_719,
input [18:0] Wgt_4_720,
input [18:0] Wgt_4_721,
input [18:0] Wgt_4_722,
input [18:0] Wgt_4_723,
input [18:0] Wgt_4_724,
input [18:0] Wgt_4_725,
input [18:0] Wgt_4_726,
input [18:0] Wgt_4_727,
input [18:0] Wgt_4_728,
input [18:0] Wgt_4_729,
input [18:0] Wgt_4_730,
input [18:0] Wgt_4_731,
input [18:0] Wgt_4_732,
input [18:0] Wgt_4_733,
input [18:0] Wgt_4_734,
input [18:0] Wgt_4_735,
input [18:0] Wgt_4_736,
input [18:0] Wgt_4_737,
input [18:0] Wgt_4_738,
input [18:0] Wgt_4_739,
input [18:0] Wgt_4_740,
input [18:0] Wgt_4_741,
input [18:0] Wgt_4_742,
input [18:0] Wgt_4_743,
input [18:0] Wgt_4_744,
input [18:0] Wgt_4_745,
input [18:0] Wgt_4_746,
input [18:0] Wgt_4_747,
input [18:0] Wgt_4_748,
input [18:0] Wgt_4_749,
input [18:0] Wgt_4_750,
input [18:0] Wgt_4_751,
input [18:0] Wgt_4_752,
input [18:0] Wgt_4_753,
input [18:0] Wgt_4_754,
input [18:0] Wgt_4_755,
input [18:0] Wgt_4_756,
input [18:0] Wgt_4_757,
input [18:0] Wgt_4_758,
input [18:0] Wgt_4_759,
input [18:0] Wgt_4_760,
input [18:0] Wgt_4_761,
input [18:0] Wgt_4_762,
input [18:0] Wgt_4_763,
input [18:0] Wgt_4_764,
input [18:0] Wgt_4_765,
input [18:0] Wgt_4_766,
input [18:0] Wgt_4_767,
input [18:0] Wgt_4_768,
input [18:0] Wgt_4_769,
input [18:0] Wgt_4_770,
input [18:0] Wgt_4_771,
input [18:0] Wgt_4_772,
input [18:0] Wgt_4_773,
input [18:0] Wgt_4_774,
input [18:0] Wgt_4_775,
input [18:0] Wgt_4_776,
input [18:0] Wgt_4_777,
input [18:0] Wgt_4_778,
input [18:0] Wgt_4_779,
input [18:0] Wgt_4_780,
input [18:0] Wgt_4_781,
input [18:0] Wgt_4_782,
input [18:0] Wgt_4_783,
input [18:0] Wgt_4_784,
input [18:0] Wgt_5_0,
input [18:0] Wgt_5_1,
input [18:0] Wgt_5_2,
input [18:0] Wgt_5_3,
input [18:0] Wgt_5_4,
input [18:0] Wgt_5_5,
input [18:0] Wgt_5_6,
input [18:0] Wgt_5_7,
input [18:0] Wgt_5_8,
input [18:0] Wgt_5_9,
input [18:0] Wgt_5_10,
input [18:0] Wgt_5_11,
input [18:0] Wgt_5_12,
input [18:0] Wgt_5_13,
input [18:0] Wgt_5_14,
input [18:0] Wgt_5_15,
input [18:0] Wgt_5_16,
input [18:0] Wgt_5_17,
input [18:0] Wgt_5_18,
input [18:0] Wgt_5_19,
input [18:0] Wgt_5_20,
input [18:0] Wgt_5_21,
input [18:0] Wgt_5_22,
input [18:0] Wgt_5_23,
input [18:0] Wgt_5_24,
input [18:0] Wgt_5_25,
input [18:0] Wgt_5_26,
input [18:0] Wgt_5_27,
input [18:0] Wgt_5_28,
input [18:0] Wgt_5_29,
input [18:0] Wgt_5_30,
input [18:0] Wgt_5_31,
input [18:0] Wgt_5_32,
input [18:0] Wgt_5_33,
input [18:0] Wgt_5_34,
input [18:0] Wgt_5_35,
input [18:0] Wgt_5_36,
input [18:0] Wgt_5_37,
input [18:0] Wgt_5_38,
input [18:0] Wgt_5_39,
input [18:0] Wgt_5_40,
input [18:0] Wgt_5_41,
input [18:0] Wgt_5_42,
input [18:0] Wgt_5_43,
input [18:0] Wgt_5_44,
input [18:0] Wgt_5_45,
input [18:0] Wgt_5_46,
input [18:0] Wgt_5_47,
input [18:0] Wgt_5_48,
input [18:0] Wgt_5_49,
input [18:0] Wgt_5_50,
input [18:0] Wgt_5_51,
input [18:0] Wgt_5_52,
input [18:0] Wgt_5_53,
input [18:0] Wgt_5_54,
input [18:0] Wgt_5_55,
input [18:0] Wgt_5_56,
input [18:0] Wgt_5_57,
input [18:0] Wgt_5_58,
input [18:0] Wgt_5_59,
input [18:0] Wgt_5_60,
input [18:0] Wgt_5_61,
input [18:0] Wgt_5_62,
input [18:0] Wgt_5_63,
input [18:0] Wgt_5_64,
input [18:0] Wgt_5_65,
input [18:0] Wgt_5_66,
input [18:0] Wgt_5_67,
input [18:0] Wgt_5_68,
input [18:0] Wgt_5_69,
input [18:0] Wgt_5_70,
input [18:0] Wgt_5_71,
input [18:0] Wgt_5_72,
input [18:0] Wgt_5_73,
input [18:0] Wgt_5_74,
input [18:0] Wgt_5_75,
input [18:0] Wgt_5_76,
input [18:0] Wgt_5_77,
input [18:0] Wgt_5_78,
input [18:0] Wgt_5_79,
input [18:0] Wgt_5_80,
input [18:0] Wgt_5_81,
input [18:0] Wgt_5_82,
input [18:0] Wgt_5_83,
input [18:0] Wgt_5_84,
input [18:0] Wgt_5_85,
input [18:0] Wgt_5_86,
input [18:0] Wgt_5_87,
input [18:0] Wgt_5_88,
input [18:0] Wgt_5_89,
input [18:0] Wgt_5_90,
input [18:0] Wgt_5_91,
input [18:0] Wgt_5_92,
input [18:0] Wgt_5_93,
input [18:0] Wgt_5_94,
input [18:0] Wgt_5_95,
input [18:0] Wgt_5_96,
input [18:0] Wgt_5_97,
input [18:0] Wgt_5_98,
input [18:0] Wgt_5_99,
input [18:0] Wgt_5_100,
input [18:0] Wgt_5_101,
input [18:0] Wgt_5_102,
input [18:0] Wgt_5_103,
input [18:0] Wgt_5_104,
input [18:0] Wgt_5_105,
input [18:0] Wgt_5_106,
input [18:0] Wgt_5_107,
input [18:0] Wgt_5_108,
input [18:0] Wgt_5_109,
input [18:0] Wgt_5_110,
input [18:0] Wgt_5_111,
input [18:0] Wgt_5_112,
input [18:0] Wgt_5_113,
input [18:0] Wgt_5_114,
input [18:0] Wgt_5_115,
input [18:0] Wgt_5_116,
input [18:0] Wgt_5_117,
input [18:0] Wgt_5_118,
input [18:0] Wgt_5_119,
input [18:0] Wgt_5_120,
input [18:0] Wgt_5_121,
input [18:0] Wgt_5_122,
input [18:0] Wgt_5_123,
input [18:0] Wgt_5_124,
input [18:0] Wgt_5_125,
input [18:0] Wgt_5_126,
input [18:0] Wgt_5_127,
input [18:0] Wgt_5_128,
input [18:0] Wgt_5_129,
input [18:0] Wgt_5_130,
input [18:0] Wgt_5_131,
input [18:0] Wgt_5_132,
input [18:0] Wgt_5_133,
input [18:0] Wgt_5_134,
input [18:0] Wgt_5_135,
input [18:0] Wgt_5_136,
input [18:0] Wgt_5_137,
input [18:0] Wgt_5_138,
input [18:0] Wgt_5_139,
input [18:0] Wgt_5_140,
input [18:0] Wgt_5_141,
input [18:0] Wgt_5_142,
input [18:0] Wgt_5_143,
input [18:0] Wgt_5_144,
input [18:0] Wgt_5_145,
input [18:0] Wgt_5_146,
input [18:0] Wgt_5_147,
input [18:0] Wgt_5_148,
input [18:0] Wgt_5_149,
input [18:0] Wgt_5_150,
input [18:0] Wgt_5_151,
input [18:0] Wgt_5_152,
input [18:0] Wgt_5_153,
input [18:0] Wgt_5_154,
input [18:0] Wgt_5_155,
input [18:0] Wgt_5_156,
input [18:0] Wgt_5_157,
input [18:0] Wgt_5_158,
input [18:0] Wgt_5_159,
input [18:0] Wgt_5_160,
input [18:0] Wgt_5_161,
input [18:0] Wgt_5_162,
input [18:0] Wgt_5_163,
input [18:0] Wgt_5_164,
input [18:0] Wgt_5_165,
input [18:0] Wgt_5_166,
input [18:0] Wgt_5_167,
input [18:0] Wgt_5_168,
input [18:0] Wgt_5_169,
input [18:0] Wgt_5_170,
input [18:0] Wgt_5_171,
input [18:0] Wgt_5_172,
input [18:0] Wgt_5_173,
input [18:0] Wgt_5_174,
input [18:0] Wgt_5_175,
input [18:0] Wgt_5_176,
input [18:0] Wgt_5_177,
input [18:0] Wgt_5_178,
input [18:0] Wgt_5_179,
input [18:0] Wgt_5_180,
input [18:0] Wgt_5_181,
input [18:0] Wgt_5_182,
input [18:0] Wgt_5_183,
input [18:0] Wgt_5_184,
input [18:0] Wgt_5_185,
input [18:0] Wgt_5_186,
input [18:0] Wgt_5_187,
input [18:0] Wgt_5_188,
input [18:0] Wgt_5_189,
input [18:0] Wgt_5_190,
input [18:0] Wgt_5_191,
input [18:0] Wgt_5_192,
input [18:0] Wgt_5_193,
input [18:0] Wgt_5_194,
input [18:0] Wgt_5_195,
input [18:0] Wgt_5_196,
input [18:0] Wgt_5_197,
input [18:0] Wgt_5_198,
input [18:0] Wgt_5_199,
input [18:0] Wgt_5_200,
input [18:0] Wgt_5_201,
input [18:0] Wgt_5_202,
input [18:0] Wgt_5_203,
input [18:0] Wgt_5_204,
input [18:0] Wgt_5_205,
input [18:0] Wgt_5_206,
input [18:0] Wgt_5_207,
input [18:0] Wgt_5_208,
input [18:0] Wgt_5_209,
input [18:0] Wgt_5_210,
input [18:0] Wgt_5_211,
input [18:0] Wgt_5_212,
input [18:0] Wgt_5_213,
input [18:0] Wgt_5_214,
input [18:0] Wgt_5_215,
input [18:0] Wgt_5_216,
input [18:0] Wgt_5_217,
input [18:0] Wgt_5_218,
input [18:0] Wgt_5_219,
input [18:0] Wgt_5_220,
input [18:0] Wgt_5_221,
input [18:0] Wgt_5_222,
input [18:0] Wgt_5_223,
input [18:0] Wgt_5_224,
input [18:0] Wgt_5_225,
input [18:0] Wgt_5_226,
input [18:0] Wgt_5_227,
input [18:0] Wgt_5_228,
input [18:0] Wgt_5_229,
input [18:0] Wgt_5_230,
input [18:0] Wgt_5_231,
input [18:0] Wgt_5_232,
input [18:0] Wgt_5_233,
input [18:0] Wgt_5_234,
input [18:0] Wgt_5_235,
input [18:0] Wgt_5_236,
input [18:0] Wgt_5_237,
input [18:0] Wgt_5_238,
input [18:0] Wgt_5_239,
input [18:0] Wgt_5_240,
input [18:0] Wgt_5_241,
input [18:0] Wgt_5_242,
input [18:0] Wgt_5_243,
input [18:0] Wgt_5_244,
input [18:0] Wgt_5_245,
input [18:0] Wgt_5_246,
input [18:0] Wgt_5_247,
input [18:0] Wgt_5_248,
input [18:0] Wgt_5_249,
input [18:0] Wgt_5_250,
input [18:0] Wgt_5_251,
input [18:0] Wgt_5_252,
input [18:0] Wgt_5_253,
input [18:0] Wgt_5_254,
input [18:0] Wgt_5_255,
input [18:0] Wgt_5_256,
input [18:0] Wgt_5_257,
input [18:0] Wgt_5_258,
input [18:0] Wgt_5_259,
input [18:0] Wgt_5_260,
input [18:0] Wgt_5_261,
input [18:0] Wgt_5_262,
input [18:0] Wgt_5_263,
input [18:0] Wgt_5_264,
input [18:0] Wgt_5_265,
input [18:0] Wgt_5_266,
input [18:0] Wgt_5_267,
input [18:0] Wgt_5_268,
input [18:0] Wgt_5_269,
input [18:0] Wgt_5_270,
input [18:0] Wgt_5_271,
input [18:0] Wgt_5_272,
input [18:0] Wgt_5_273,
input [18:0] Wgt_5_274,
input [18:0] Wgt_5_275,
input [18:0] Wgt_5_276,
input [18:0] Wgt_5_277,
input [18:0] Wgt_5_278,
input [18:0] Wgt_5_279,
input [18:0] Wgt_5_280,
input [18:0] Wgt_5_281,
input [18:0] Wgt_5_282,
input [18:0] Wgt_5_283,
input [18:0] Wgt_5_284,
input [18:0] Wgt_5_285,
input [18:0] Wgt_5_286,
input [18:0] Wgt_5_287,
input [18:0] Wgt_5_288,
input [18:0] Wgt_5_289,
input [18:0] Wgt_5_290,
input [18:0] Wgt_5_291,
input [18:0] Wgt_5_292,
input [18:0] Wgt_5_293,
input [18:0] Wgt_5_294,
input [18:0] Wgt_5_295,
input [18:0] Wgt_5_296,
input [18:0] Wgt_5_297,
input [18:0] Wgt_5_298,
input [18:0] Wgt_5_299,
input [18:0] Wgt_5_300,
input [18:0] Wgt_5_301,
input [18:0] Wgt_5_302,
input [18:0] Wgt_5_303,
input [18:0] Wgt_5_304,
input [18:0] Wgt_5_305,
input [18:0] Wgt_5_306,
input [18:0] Wgt_5_307,
input [18:0] Wgt_5_308,
input [18:0] Wgt_5_309,
input [18:0] Wgt_5_310,
input [18:0] Wgt_5_311,
input [18:0] Wgt_5_312,
input [18:0] Wgt_5_313,
input [18:0] Wgt_5_314,
input [18:0] Wgt_5_315,
input [18:0] Wgt_5_316,
input [18:0] Wgt_5_317,
input [18:0] Wgt_5_318,
input [18:0] Wgt_5_319,
input [18:0] Wgt_5_320,
input [18:0] Wgt_5_321,
input [18:0] Wgt_5_322,
input [18:0] Wgt_5_323,
input [18:0] Wgt_5_324,
input [18:0] Wgt_5_325,
input [18:0] Wgt_5_326,
input [18:0] Wgt_5_327,
input [18:0] Wgt_5_328,
input [18:0] Wgt_5_329,
input [18:0] Wgt_5_330,
input [18:0] Wgt_5_331,
input [18:0] Wgt_5_332,
input [18:0] Wgt_5_333,
input [18:0] Wgt_5_334,
input [18:0] Wgt_5_335,
input [18:0] Wgt_5_336,
input [18:0] Wgt_5_337,
input [18:0] Wgt_5_338,
input [18:0] Wgt_5_339,
input [18:0] Wgt_5_340,
input [18:0] Wgt_5_341,
input [18:0] Wgt_5_342,
input [18:0] Wgt_5_343,
input [18:0] Wgt_5_344,
input [18:0] Wgt_5_345,
input [18:0] Wgt_5_346,
input [18:0] Wgt_5_347,
input [18:0] Wgt_5_348,
input [18:0] Wgt_5_349,
input [18:0] Wgt_5_350,
input [18:0] Wgt_5_351,
input [18:0] Wgt_5_352,
input [18:0] Wgt_5_353,
input [18:0] Wgt_5_354,
input [18:0] Wgt_5_355,
input [18:0] Wgt_5_356,
input [18:0] Wgt_5_357,
input [18:0] Wgt_5_358,
input [18:0] Wgt_5_359,
input [18:0] Wgt_5_360,
input [18:0] Wgt_5_361,
input [18:0] Wgt_5_362,
input [18:0] Wgt_5_363,
input [18:0] Wgt_5_364,
input [18:0] Wgt_5_365,
input [18:0] Wgt_5_366,
input [18:0] Wgt_5_367,
input [18:0] Wgt_5_368,
input [18:0] Wgt_5_369,
input [18:0] Wgt_5_370,
input [18:0] Wgt_5_371,
input [18:0] Wgt_5_372,
input [18:0] Wgt_5_373,
input [18:0] Wgt_5_374,
input [18:0] Wgt_5_375,
input [18:0] Wgt_5_376,
input [18:0] Wgt_5_377,
input [18:0] Wgt_5_378,
input [18:0] Wgt_5_379,
input [18:0] Wgt_5_380,
input [18:0] Wgt_5_381,
input [18:0] Wgt_5_382,
input [18:0] Wgt_5_383,
input [18:0] Wgt_5_384,
input [18:0] Wgt_5_385,
input [18:0] Wgt_5_386,
input [18:0] Wgt_5_387,
input [18:0] Wgt_5_388,
input [18:0] Wgt_5_389,
input [18:0] Wgt_5_390,
input [18:0] Wgt_5_391,
input [18:0] Wgt_5_392,
input [18:0] Wgt_5_393,
input [18:0] Wgt_5_394,
input [18:0] Wgt_5_395,
input [18:0] Wgt_5_396,
input [18:0] Wgt_5_397,
input [18:0] Wgt_5_398,
input [18:0] Wgt_5_399,
input [18:0] Wgt_5_400,
input [18:0] Wgt_5_401,
input [18:0] Wgt_5_402,
input [18:0] Wgt_5_403,
input [18:0] Wgt_5_404,
input [18:0] Wgt_5_405,
input [18:0] Wgt_5_406,
input [18:0] Wgt_5_407,
input [18:0] Wgt_5_408,
input [18:0] Wgt_5_409,
input [18:0] Wgt_5_410,
input [18:0] Wgt_5_411,
input [18:0] Wgt_5_412,
input [18:0] Wgt_5_413,
input [18:0] Wgt_5_414,
input [18:0] Wgt_5_415,
input [18:0] Wgt_5_416,
input [18:0] Wgt_5_417,
input [18:0] Wgt_5_418,
input [18:0] Wgt_5_419,
input [18:0] Wgt_5_420,
input [18:0] Wgt_5_421,
input [18:0] Wgt_5_422,
input [18:0] Wgt_5_423,
input [18:0] Wgt_5_424,
input [18:0] Wgt_5_425,
input [18:0] Wgt_5_426,
input [18:0] Wgt_5_427,
input [18:0] Wgt_5_428,
input [18:0] Wgt_5_429,
input [18:0] Wgt_5_430,
input [18:0] Wgt_5_431,
input [18:0] Wgt_5_432,
input [18:0] Wgt_5_433,
input [18:0] Wgt_5_434,
input [18:0] Wgt_5_435,
input [18:0] Wgt_5_436,
input [18:0] Wgt_5_437,
input [18:0] Wgt_5_438,
input [18:0] Wgt_5_439,
input [18:0] Wgt_5_440,
input [18:0] Wgt_5_441,
input [18:0] Wgt_5_442,
input [18:0] Wgt_5_443,
input [18:0] Wgt_5_444,
input [18:0] Wgt_5_445,
input [18:0] Wgt_5_446,
input [18:0] Wgt_5_447,
input [18:0] Wgt_5_448,
input [18:0] Wgt_5_449,
input [18:0] Wgt_5_450,
input [18:0] Wgt_5_451,
input [18:0] Wgt_5_452,
input [18:0] Wgt_5_453,
input [18:0] Wgt_5_454,
input [18:0] Wgt_5_455,
input [18:0] Wgt_5_456,
input [18:0] Wgt_5_457,
input [18:0] Wgt_5_458,
input [18:0] Wgt_5_459,
input [18:0] Wgt_5_460,
input [18:0] Wgt_5_461,
input [18:0] Wgt_5_462,
input [18:0] Wgt_5_463,
input [18:0] Wgt_5_464,
input [18:0] Wgt_5_465,
input [18:0] Wgt_5_466,
input [18:0] Wgt_5_467,
input [18:0] Wgt_5_468,
input [18:0] Wgt_5_469,
input [18:0] Wgt_5_470,
input [18:0] Wgt_5_471,
input [18:0] Wgt_5_472,
input [18:0] Wgt_5_473,
input [18:0] Wgt_5_474,
input [18:0] Wgt_5_475,
input [18:0] Wgt_5_476,
input [18:0] Wgt_5_477,
input [18:0] Wgt_5_478,
input [18:0] Wgt_5_479,
input [18:0] Wgt_5_480,
input [18:0] Wgt_5_481,
input [18:0] Wgt_5_482,
input [18:0] Wgt_5_483,
input [18:0] Wgt_5_484,
input [18:0] Wgt_5_485,
input [18:0] Wgt_5_486,
input [18:0] Wgt_5_487,
input [18:0] Wgt_5_488,
input [18:0] Wgt_5_489,
input [18:0] Wgt_5_490,
input [18:0] Wgt_5_491,
input [18:0] Wgt_5_492,
input [18:0] Wgt_5_493,
input [18:0] Wgt_5_494,
input [18:0] Wgt_5_495,
input [18:0] Wgt_5_496,
input [18:0] Wgt_5_497,
input [18:0] Wgt_5_498,
input [18:0] Wgt_5_499,
input [18:0] Wgt_5_500,
input [18:0] Wgt_5_501,
input [18:0] Wgt_5_502,
input [18:0] Wgt_5_503,
input [18:0] Wgt_5_504,
input [18:0] Wgt_5_505,
input [18:0] Wgt_5_506,
input [18:0] Wgt_5_507,
input [18:0] Wgt_5_508,
input [18:0] Wgt_5_509,
input [18:0] Wgt_5_510,
input [18:0] Wgt_5_511,
input [18:0] Wgt_5_512,
input [18:0] Wgt_5_513,
input [18:0] Wgt_5_514,
input [18:0] Wgt_5_515,
input [18:0] Wgt_5_516,
input [18:0] Wgt_5_517,
input [18:0] Wgt_5_518,
input [18:0] Wgt_5_519,
input [18:0] Wgt_5_520,
input [18:0] Wgt_5_521,
input [18:0] Wgt_5_522,
input [18:0] Wgt_5_523,
input [18:0] Wgt_5_524,
input [18:0] Wgt_5_525,
input [18:0] Wgt_5_526,
input [18:0] Wgt_5_527,
input [18:0] Wgt_5_528,
input [18:0] Wgt_5_529,
input [18:0] Wgt_5_530,
input [18:0] Wgt_5_531,
input [18:0] Wgt_5_532,
input [18:0] Wgt_5_533,
input [18:0] Wgt_5_534,
input [18:0] Wgt_5_535,
input [18:0] Wgt_5_536,
input [18:0] Wgt_5_537,
input [18:0] Wgt_5_538,
input [18:0] Wgt_5_539,
input [18:0] Wgt_5_540,
input [18:0] Wgt_5_541,
input [18:0] Wgt_5_542,
input [18:0] Wgt_5_543,
input [18:0] Wgt_5_544,
input [18:0] Wgt_5_545,
input [18:0] Wgt_5_546,
input [18:0] Wgt_5_547,
input [18:0] Wgt_5_548,
input [18:0] Wgt_5_549,
input [18:0] Wgt_5_550,
input [18:0] Wgt_5_551,
input [18:0] Wgt_5_552,
input [18:0] Wgt_5_553,
input [18:0] Wgt_5_554,
input [18:0] Wgt_5_555,
input [18:0] Wgt_5_556,
input [18:0] Wgt_5_557,
input [18:0] Wgt_5_558,
input [18:0] Wgt_5_559,
input [18:0] Wgt_5_560,
input [18:0] Wgt_5_561,
input [18:0] Wgt_5_562,
input [18:0] Wgt_5_563,
input [18:0] Wgt_5_564,
input [18:0] Wgt_5_565,
input [18:0] Wgt_5_566,
input [18:0] Wgt_5_567,
input [18:0] Wgt_5_568,
input [18:0] Wgt_5_569,
input [18:0] Wgt_5_570,
input [18:0] Wgt_5_571,
input [18:0] Wgt_5_572,
input [18:0] Wgt_5_573,
input [18:0] Wgt_5_574,
input [18:0] Wgt_5_575,
input [18:0] Wgt_5_576,
input [18:0] Wgt_5_577,
input [18:0] Wgt_5_578,
input [18:0] Wgt_5_579,
input [18:0] Wgt_5_580,
input [18:0] Wgt_5_581,
input [18:0] Wgt_5_582,
input [18:0] Wgt_5_583,
input [18:0] Wgt_5_584,
input [18:0] Wgt_5_585,
input [18:0] Wgt_5_586,
input [18:0] Wgt_5_587,
input [18:0] Wgt_5_588,
input [18:0] Wgt_5_589,
input [18:0] Wgt_5_590,
input [18:0] Wgt_5_591,
input [18:0] Wgt_5_592,
input [18:0] Wgt_5_593,
input [18:0] Wgt_5_594,
input [18:0] Wgt_5_595,
input [18:0] Wgt_5_596,
input [18:0] Wgt_5_597,
input [18:0] Wgt_5_598,
input [18:0] Wgt_5_599,
input [18:0] Wgt_5_600,
input [18:0] Wgt_5_601,
input [18:0] Wgt_5_602,
input [18:0] Wgt_5_603,
input [18:0] Wgt_5_604,
input [18:0] Wgt_5_605,
input [18:0] Wgt_5_606,
input [18:0] Wgt_5_607,
input [18:0] Wgt_5_608,
input [18:0] Wgt_5_609,
input [18:0] Wgt_5_610,
input [18:0] Wgt_5_611,
input [18:0] Wgt_5_612,
input [18:0] Wgt_5_613,
input [18:0] Wgt_5_614,
input [18:0] Wgt_5_615,
input [18:0] Wgt_5_616,
input [18:0] Wgt_5_617,
input [18:0] Wgt_5_618,
input [18:0] Wgt_5_619,
input [18:0] Wgt_5_620,
input [18:0] Wgt_5_621,
input [18:0] Wgt_5_622,
input [18:0] Wgt_5_623,
input [18:0] Wgt_5_624,
input [18:0] Wgt_5_625,
input [18:0] Wgt_5_626,
input [18:0] Wgt_5_627,
input [18:0] Wgt_5_628,
input [18:0] Wgt_5_629,
input [18:0] Wgt_5_630,
input [18:0] Wgt_5_631,
input [18:0] Wgt_5_632,
input [18:0] Wgt_5_633,
input [18:0] Wgt_5_634,
input [18:0] Wgt_5_635,
input [18:0] Wgt_5_636,
input [18:0] Wgt_5_637,
input [18:0] Wgt_5_638,
input [18:0] Wgt_5_639,
input [18:0] Wgt_5_640,
input [18:0] Wgt_5_641,
input [18:0] Wgt_5_642,
input [18:0] Wgt_5_643,
input [18:0] Wgt_5_644,
input [18:0] Wgt_5_645,
input [18:0] Wgt_5_646,
input [18:0] Wgt_5_647,
input [18:0] Wgt_5_648,
input [18:0] Wgt_5_649,
input [18:0] Wgt_5_650,
input [18:0] Wgt_5_651,
input [18:0] Wgt_5_652,
input [18:0] Wgt_5_653,
input [18:0] Wgt_5_654,
input [18:0] Wgt_5_655,
input [18:0] Wgt_5_656,
input [18:0] Wgt_5_657,
input [18:0] Wgt_5_658,
input [18:0] Wgt_5_659,
input [18:0] Wgt_5_660,
input [18:0] Wgt_5_661,
input [18:0] Wgt_5_662,
input [18:0] Wgt_5_663,
input [18:0] Wgt_5_664,
input [18:0] Wgt_5_665,
input [18:0] Wgt_5_666,
input [18:0] Wgt_5_667,
input [18:0] Wgt_5_668,
input [18:0] Wgt_5_669,
input [18:0] Wgt_5_670,
input [18:0] Wgt_5_671,
input [18:0] Wgt_5_672,
input [18:0] Wgt_5_673,
input [18:0] Wgt_5_674,
input [18:0] Wgt_5_675,
input [18:0] Wgt_5_676,
input [18:0] Wgt_5_677,
input [18:0] Wgt_5_678,
input [18:0] Wgt_5_679,
input [18:0] Wgt_5_680,
input [18:0] Wgt_5_681,
input [18:0] Wgt_5_682,
input [18:0] Wgt_5_683,
input [18:0] Wgt_5_684,
input [18:0] Wgt_5_685,
input [18:0] Wgt_5_686,
input [18:0] Wgt_5_687,
input [18:0] Wgt_5_688,
input [18:0] Wgt_5_689,
input [18:0] Wgt_5_690,
input [18:0] Wgt_5_691,
input [18:0] Wgt_5_692,
input [18:0] Wgt_5_693,
input [18:0] Wgt_5_694,
input [18:0] Wgt_5_695,
input [18:0] Wgt_5_696,
input [18:0] Wgt_5_697,
input [18:0] Wgt_5_698,
input [18:0] Wgt_5_699,
input [18:0] Wgt_5_700,
input [18:0] Wgt_5_701,
input [18:0] Wgt_5_702,
input [18:0] Wgt_5_703,
input [18:0] Wgt_5_704,
input [18:0] Wgt_5_705,
input [18:0] Wgt_5_706,
input [18:0] Wgt_5_707,
input [18:0] Wgt_5_708,
input [18:0] Wgt_5_709,
input [18:0] Wgt_5_710,
input [18:0] Wgt_5_711,
input [18:0] Wgt_5_712,
input [18:0] Wgt_5_713,
input [18:0] Wgt_5_714,
input [18:0] Wgt_5_715,
input [18:0] Wgt_5_716,
input [18:0] Wgt_5_717,
input [18:0] Wgt_5_718,
input [18:0] Wgt_5_719,
input [18:0] Wgt_5_720,
input [18:0] Wgt_5_721,
input [18:0] Wgt_5_722,
input [18:0] Wgt_5_723,
input [18:0] Wgt_5_724,
input [18:0] Wgt_5_725,
input [18:0] Wgt_5_726,
input [18:0] Wgt_5_727,
input [18:0] Wgt_5_728,
input [18:0] Wgt_5_729,
input [18:0] Wgt_5_730,
input [18:0] Wgt_5_731,
input [18:0] Wgt_5_732,
input [18:0] Wgt_5_733,
input [18:0] Wgt_5_734,
input [18:0] Wgt_5_735,
input [18:0] Wgt_5_736,
input [18:0] Wgt_5_737,
input [18:0] Wgt_5_738,
input [18:0] Wgt_5_739,
input [18:0] Wgt_5_740,
input [18:0] Wgt_5_741,
input [18:0] Wgt_5_742,
input [18:0] Wgt_5_743,
input [18:0] Wgt_5_744,
input [18:0] Wgt_5_745,
input [18:0] Wgt_5_746,
input [18:0] Wgt_5_747,
input [18:0] Wgt_5_748,
input [18:0] Wgt_5_749,
input [18:0] Wgt_5_750,
input [18:0] Wgt_5_751,
input [18:0] Wgt_5_752,
input [18:0] Wgt_5_753,
input [18:0] Wgt_5_754,
input [18:0] Wgt_5_755,
input [18:0] Wgt_5_756,
input [18:0] Wgt_5_757,
input [18:0] Wgt_5_758,
input [18:0] Wgt_5_759,
input [18:0] Wgt_5_760,
input [18:0] Wgt_5_761,
input [18:0] Wgt_5_762,
input [18:0] Wgt_5_763,
input [18:0] Wgt_5_764,
input [18:0] Wgt_5_765,
input [18:0] Wgt_5_766,
input [18:0] Wgt_5_767,
input [18:0] Wgt_5_768,
input [18:0] Wgt_5_769,
input [18:0] Wgt_5_770,
input [18:0] Wgt_5_771,
input [18:0] Wgt_5_772,
input [18:0] Wgt_5_773,
input [18:0] Wgt_5_774,
input [18:0] Wgt_5_775,
input [18:0] Wgt_5_776,
input [18:0] Wgt_5_777,
input [18:0] Wgt_5_778,
input [18:0] Wgt_5_779,
input [18:0] Wgt_5_780,
input [18:0] Wgt_5_781,
input [18:0] Wgt_5_782,
input [18:0] Wgt_5_783,
input [18:0] Wgt_5_784,
input [18:0] Wgt_6_0,
input [18:0] Wgt_6_1,
input [18:0] Wgt_6_2,
input [18:0] Wgt_6_3,
input [18:0] Wgt_6_4,
input [18:0] Wgt_6_5,
input [18:0] Wgt_6_6,
input [18:0] Wgt_6_7,
input [18:0] Wgt_6_8,
input [18:0] Wgt_6_9,
input [18:0] Wgt_6_10,
input [18:0] Wgt_6_11,
input [18:0] Wgt_6_12,
input [18:0] Wgt_6_13,
input [18:0] Wgt_6_14,
input [18:0] Wgt_6_15,
input [18:0] Wgt_6_16,
input [18:0] Wgt_6_17,
input [18:0] Wgt_6_18,
input [18:0] Wgt_6_19,
input [18:0] Wgt_6_20,
input [18:0] Wgt_6_21,
input [18:0] Wgt_6_22,
input [18:0] Wgt_6_23,
input [18:0] Wgt_6_24,
input [18:0] Wgt_6_25,
input [18:0] Wgt_6_26,
input [18:0] Wgt_6_27,
input [18:0] Wgt_6_28,
input [18:0] Wgt_6_29,
input [18:0] Wgt_6_30,
input [18:0] Wgt_6_31,
input [18:0] Wgt_6_32,
input [18:0] Wgt_6_33,
input [18:0] Wgt_6_34,
input [18:0] Wgt_6_35,
input [18:0] Wgt_6_36,
input [18:0] Wgt_6_37,
input [18:0] Wgt_6_38,
input [18:0] Wgt_6_39,
input [18:0] Wgt_6_40,
input [18:0] Wgt_6_41,
input [18:0] Wgt_6_42,
input [18:0] Wgt_6_43,
input [18:0] Wgt_6_44,
input [18:0] Wgt_6_45,
input [18:0] Wgt_6_46,
input [18:0] Wgt_6_47,
input [18:0] Wgt_6_48,
input [18:0] Wgt_6_49,
input [18:0] Wgt_6_50,
input [18:0] Wgt_6_51,
input [18:0] Wgt_6_52,
input [18:0] Wgt_6_53,
input [18:0] Wgt_6_54,
input [18:0] Wgt_6_55,
input [18:0] Wgt_6_56,
input [18:0] Wgt_6_57,
input [18:0] Wgt_6_58,
input [18:0] Wgt_6_59,
input [18:0] Wgt_6_60,
input [18:0] Wgt_6_61,
input [18:0] Wgt_6_62,
input [18:0] Wgt_6_63,
input [18:0] Wgt_6_64,
input [18:0] Wgt_6_65,
input [18:0] Wgt_6_66,
input [18:0] Wgt_6_67,
input [18:0] Wgt_6_68,
input [18:0] Wgt_6_69,
input [18:0] Wgt_6_70,
input [18:0] Wgt_6_71,
input [18:0] Wgt_6_72,
input [18:0] Wgt_6_73,
input [18:0] Wgt_6_74,
input [18:0] Wgt_6_75,
input [18:0] Wgt_6_76,
input [18:0] Wgt_6_77,
input [18:0] Wgt_6_78,
input [18:0] Wgt_6_79,
input [18:0] Wgt_6_80,
input [18:0] Wgt_6_81,
input [18:0] Wgt_6_82,
input [18:0] Wgt_6_83,
input [18:0] Wgt_6_84,
input [18:0] Wgt_6_85,
input [18:0] Wgt_6_86,
input [18:0] Wgt_6_87,
input [18:0] Wgt_6_88,
input [18:0] Wgt_6_89,
input [18:0] Wgt_6_90,
input [18:0] Wgt_6_91,
input [18:0] Wgt_6_92,
input [18:0] Wgt_6_93,
input [18:0] Wgt_6_94,
input [18:0] Wgt_6_95,
input [18:0] Wgt_6_96,
input [18:0] Wgt_6_97,
input [18:0] Wgt_6_98,
input [18:0] Wgt_6_99,
input [18:0] Wgt_6_100,
input [18:0] Wgt_6_101,
input [18:0] Wgt_6_102,
input [18:0] Wgt_6_103,
input [18:0] Wgt_6_104,
input [18:0] Wgt_6_105,
input [18:0] Wgt_6_106,
input [18:0] Wgt_6_107,
input [18:0] Wgt_6_108,
input [18:0] Wgt_6_109,
input [18:0] Wgt_6_110,
input [18:0] Wgt_6_111,
input [18:0] Wgt_6_112,
input [18:0] Wgt_6_113,
input [18:0] Wgt_6_114,
input [18:0] Wgt_6_115,
input [18:0] Wgt_6_116,
input [18:0] Wgt_6_117,
input [18:0] Wgt_6_118,
input [18:0] Wgt_6_119,
input [18:0] Wgt_6_120,
input [18:0] Wgt_6_121,
input [18:0] Wgt_6_122,
input [18:0] Wgt_6_123,
input [18:0] Wgt_6_124,
input [18:0] Wgt_6_125,
input [18:0] Wgt_6_126,
input [18:0] Wgt_6_127,
input [18:0] Wgt_6_128,
input [18:0] Wgt_6_129,
input [18:0] Wgt_6_130,
input [18:0] Wgt_6_131,
input [18:0] Wgt_6_132,
input [18:0] Wgt_6_133,
input [18:0] Wgt_6_134,
input [18:0] Wgt_6_135,
input [18:0] Wgt_6_136,
input [18:0] Wgt_6_137,
input [18:0] Wgt_6_138,
input [18:0] Wgt_6_139,
input [18:0] Wgt_6_140,
input [18:0] Wgt_6_141,
input [18:0] Wgt_6_142,
input [18:0] Wgt_6_143,
input [18:0] Wgt_6_144,
input [18:0] Wgt_6_145,
input [18:0] Wgt_6_146,
input [18:0] Wgt_6_147,
input [18:0] Wgt_6_148,
input [18:0] Wgt_6_149,
input [18:0] Wgt_6_150,
input [18:0] Wgt_6_151,
input [18:0] Wgt_6_152,
input [18:0] Wgt_6_153,
input [18:0] Wgt_6_154,
input [18:0] Wgt_6_155,
input [18:0] Wgt_6_156,
input [18:0] Wgt_6_157,
input [18:0] Wgt_6_158,
input [18:0] Wgt_6_159,
input [18:0] Wgt_6_160,
input [18:0] Wgt_6_161,
input [18:0] Wgt_6_162,
input [18:0] Wgt_6_163,
input [18:0] Wgt_6_164,
input [18:0] Wgt_6_165,
input [18:0] Wgt_6_166,
input [18:0] Wgt_6_167,
input [18:0] Wgt_6_168,
input [18:0] Wgt_6_169,
input [18:0] Wgt_6_170,
input [18:0] Wgt_6_171,
input [18:0] Wgt_6_172,
input [18:0] Wgt_6_173,
input [18:0] Wgt_6_174,
input [18:0] Wgt_6_175,
input [18:0] Wgt_6_176,
input [18:0] Wgt_6_177,
input [18:0] Wgt_6_178,
input [18:0] Wgt_6_179,
input [18:0] Wgt_6_180,
input [18:0] Wgt_6_181,
input [18:0] Wgt_6_182,
input [18:0] Wgt_6_183,
input [18:0] Wgt_6_184,
input [18:0] Wgt_6_185,
input [18:0] Wgt_6_186,
input [18:0] Wgt_6_187,
input [18:0] Wgt_6_188,
input [18:0] Wgt_6_189,
input [18:0] Wgt_6_190,
input [18:0] Wgt_6_191,
input [18:0] Wgt_6_192,
input [18:0] Wgt_6_193,
input [18:0] Wgt_6_194,
input [18:0] Wgt_6_195,
input [18:0] Wgt_6_196,
input [18:0] Wgt_6_197,
input [18:0] Wgt_6_198,
input [18:0] Wgt_6_199,
input [18:0] Wgt_6_200,
input [18:0] Wgt_6_201,
input [18:0] Wgt_6_202,
input [18:0] Wgt_6_203,
input [18:0] Wgt_6_204,
input [18:0] Wgt_6_205,
input [18:0] Wgt_6_206,
input [18:0] Wgt_6_207,
input [18:0] Wgt_6_208,
input [18:0] Wgt_6_209,
input [18:0] Wgt_6_210,
input [18:0] Wgt_6_211,
input [18:0] Wgt_6_212,
input [18:0] Wgt_6_213,
input [18:0] Wgt_6_214,
input [18:0] Wgt_6_215,
input [18:0] Wgt_6_216,
input [18:0] Wgt_6_217,
input [18:0] Wgt_6_218,
input [18:0] Wgt_6_219,
input [18:0] Wgt_6_220,
input [18:0] Wgt_6_221,
input [18:0] Wgt_6_222,
input [18:0] Wgt_6_223,
input [18:0] Wgt_6_224,
input [18:0] Wgt_6_225,
input [18:0] Wgt_6_226,
input [18:0] Wgt_6_227,
input [18:0] Wgt_6_228,
input [18:0] Wgt_6_229,
input [18:0] Wgt_6_230,
input [18:0] Wgt_6_231,
input [18:0] Wgt_6_232,
input [18:0] Wgt_6_233,
input [18:0] Wgt_6_234,
input [18:0] Wgt_6_235,
input [18:0] Wgt_6_236,
input [18:0] Wgt_6_237,
input [18:0] Wgt_6_238,
input [18:0] Wgt_6_239,
input [18:0] Wgt_6_240,
input [18:0] Wgt_6_241,
input [18:0] Wgt_6_242,
input [18:0] Wgt_6_243,
input [18:0] Wgt_6_244,
input [18:0] Wgt_6_245,
input [18:0] Wgt_6_246,
input [18:0] Wgt_6_247,
input [18:0] Wgt_6_248,
input [18:0] Wgt_6_249,
input [18:0] Wgt_6_250,
input [18:0] Wgt_6_251,
input [18:0] Wgt_6_252,
input [18:0] Wgt_6_253,
input [18:0] Wgt_6_254,
input [18:0] Wgt_6_255,
input [18:0] Wgt_6_256,
input [18:0] Wgt_6_257,
input [18:0] Wgt_6_258,
input [18:0] Wgt_6_259,
input [18:0] Wgt_6_260,
input [18:0] Wgt_6_261,
input [18:0] Wgt_6_262,
input [18:0] Wgt_6_263,
input [18:0] Wgt_6_264,
input [18:0] Wgt_6_265,
input [18:0] Wgt_6_266,
input [18:0] Wgt_6_267,
input [18:0] Wgt_6_268,
input [18:0] Wgt_6_269,
input [18:0] Wgt_6_270,
input [18:0] Wgt_6_271,
input [18:0] Wgt_6_272,
input [18:0] Wgt_6_273,
input [18:0] Wgt_6_274,
input [18:0] Wgt_6_275,
input [18:0] Wgt_6_276,
input [18:0] Wgt_6_277,
input [18:0] Wgt_6_278,
input [18:0] Wgt_6_279,
input [18:0] Wgt_6_280,
input [18:0] Wgt_6_281,
input [18:0] Wgt_6_282,
input [18:0] Wgt_6_283,
input [18:0] Wgt_6_284,
input [18:0] Wgt_6_285,
input [18:0] Wgt_6_286,
input [18:0] Wgt_6_287,
input [18:0] Wgt_6_288,
input [18:0] Wgt_6_289,
input [18:0] Wgt_6_290,
input [18:0] Wgt_6_291,
input [18:0] Wgt_6_292,
input [18:0] Wgt_6_293,
input [18:0] Wgt_6_294,
input [18:0] Wgt_6_295,
input [18:0] Wgt_6_296,
input [18:0] Wgt_6_297,
input [18:0] Wgt_6_298,
input [18:0] Wgt_6_299,
input [18:0] Wgt_6_300,
input [18:0] Wgt_6_301,
input [18:0] Wgt_6_302,
input [18:0] Wgt_6_303,
input [18:0] Wgt_6_304,
input [18:0] Wgt_6_305,
input [18:0] Wgt_6_306,
input [18:0] Wgt_6_307,
input [18:0] Wgt_6_308,
input [18:0] Wgt_6_309,
input [18:0] Wgt_6_310,
input [18:0] Wgt_6_311,
input [18:0] Wgt_6_312,
input [18:0] Wgt_6_313,
input [18:0] Wgt_6_314,
input [18:0] Wgt_6_315,
input [18:0] Wgt_6_316,
input [18:0] Wgt_6_317,
input [18:0] Wgt_6_318,
input [18:0] Wgt_6_319,
input [18:0] Wgt_6_320,
input [18:0] Wgt_6_321,
input [18:0] Wgt_6_322,
input [18:0] Wgt_6_323,
input [18:0] Wgt_6_324,
input [18:0] Wgt_6_325,
input [18:0] Wgt_6_326,
input [18:0] Wgt_6_327,
input [18:0] Wgt_6_328,
input [18:0] Wgt_6_329,
input [18:0] Wgt_6_330,
input [18:0] Wgt_6_331,
input [18:0] Wgt_6_332,
input [18:0] Wgt_6_333,
input [18:0] Wgt_6_334,
input [18:0] Wgt_6_335,
input [18:0] Wgt_6_336,
input [18:0] Wgt_6_337,
input [18:0] Wgt_6_338,
input [18:0] Wgt_6_339,
input [18:0] Wgt_6_340,
input [18:0] Wgt_6_341,
input [18:0] Wgt_6_342,
input [18:0] Wgt_6_343,
input [18:0] Wgt_6_344,
input [18:0] Wgt_6_345,
input [18:0] Wgt_6_346,
input [18:0] Wgt_6_347,
input [18:0] Wgt_6_348,
input [18:0] Wgt_6_349,
input [18:0] Wgt_6_350,
input [18:0] Wgt_6_351,
input [18:0] Wgt_6_352,
input [18:0] Wgt_6_353,
input [18:0] Wgt_6_354,
input [18:0] Wgt_6_355,
input [18:0] Wgt_6_356,
input [18:0] Wgt_6_357,
input [18:0] Wgt_6_358,
input [18:0] Wgt_6_359,
input [18:0] Wgt_6_360,
input [18:0] Wgt_6_361,
input [18:0] Wgt_6_362,
input [18:0] Wgt_6_363,
input [18:0] Wgt_6_364,
input [18:0] Wgt_6_365,
input [18:0] Wgt_6_366,
input [18:0] Wgt_6_367,
input [18:0] Wgt_6_368,
input [18:0] Wgt_6_369,
input [18:0] Wgt_6_370,
input [18:0] Wgt_6_371,
input [18:0] Wgt_6_372,
input [18:0] Wgt_6_373,
input [18:0] Wgt_6_374,
input [18:0] Wgt_6_375,
input [18:0] Wgt_6_376,
input [18:0] Wgt_6_377,
input [18:0] Wgt_6_378,
input [18:0] Wgt_6_379,
input [18:0] Wgt_6_380,
input [18:0] Wgt_6_381,
input [18:0] Wgt_6_382,
input [18:0] Wgt_6_383,
input [18:0] Wgt_6_384,
input [18:0] Wgt_6_385,
input [18:0] Wgt_6_386,
input [18:0] Wgt_6_387,
input [18:0] Wgt_6_388,
input [18:0] Wgt_6_389,
input [18:0] Wgt_6_390,
input [18:0] Wgt_6_391,
input [18:0] Wgt_6_392,
input [18:0] Wgt_6_393,
input [18:0] Wgt_6_394,
input [18:0] Wgt_6_395,
input [18:0] Wgt_6_396,
input [18:0] Wgt_6_397,
input [18:0] Wgt_6_398,
input [18:0] Wgt_6_399,
input [18:0] Wgt_6_400,
input [18:0] Wgt_6_401,
input [18:0] Wgt_6_402,
input [18:0] Wgt_6_403,
input [18:0] Wgt_6_404,
input [18:0] Wgt_6_405,
input [18:0] Wgt_6_406,
input [18:0] Wgt_6_407,
input [18:0] Wgt_6_408,
input [18:0] Wgt_6_409,
input [18:0] Wgt_6_410,
input [18:0] Wgt_6_411,
input [18:0] Wgt_6_412,
input [18:0] Wgt_6_413,
input [18:0] Wgt_6_414,
input [18:0] Wgt_6_415,
input [18:0] Wgt_6_416,
input [18:0] Wgt_6_417,
input [18:0] Wgt_6_418,
input [18:0] Wgt_6_419,
input [18:0] Wgt_6_420,
input [18:0] Wgt_6_421,
input [18:0] Wgt_6_422,
input [18:0] Wgt_6_423,
input [18:0] Wgt_6_424,
input [18:0] Wgt_6_425,
input [18:0] Wgt_6_426,
input [18:0] Wgt_6_427,
input [18:0] Wgt_6_428,
input [18:0] Wgt_6_429,
input [18:0] Wgt_6_430,
input [18:0] Wgt_6_431,
input [18:0] Wgt_6_432,
input [18:0] Wgt_6_433,
input [18:0] Wgt_6_434,
input [18:0] Wgt_6_435,
input [18:0] Wgt_6_436,
input [18:0] Wgt_6_437,
input [18:0] Wgt_6_438,
input [18:0] Wgt_6_439,
input [18:0] Wgt_6_440,
input [18:0] Wgt_6_441,
input [18:0] Wgt_6_442,
input [18:0] Wgt_6_443,
input [18:0] Wgt_6_444,
input [18:0] Wgt_6_445,
input [18:0] Wgt_6_446,
input [18:0] Wgt_6_447,
input [18:0] Wgt_6_448,
input [18:0] Wgt_6_449,
input [18:0] Wgt_6_450,
input [18:0] Wgt_6_451,
input [18:0] Wgt_6_452,
input [18:0] Wgt_6_453,
input [18:0] Wgt_6_454,
input [18:0] Wgt_6_455,
input [18:0] Wgt_6_456,
input [18:0] Wgt_6_457,
input [18:0] Wgt_6_458,
input [18:0] Wgt_6_459,
input [18:0] Wgt_6_460,
input [18:0] Wgt_6_461,
input [18:0] Wgt_6_462,
input [18:0] Wgt_6_463,
input [18:0] Wgt_6_464,
input [18:0] Wgt_6_465,
input [18:0] Wgt_6_466,
input [18:0] Wgt_6_467,
input [18:0] Wgt_6_468,
input [18:0] Wgt_6_469,
input [18:0] Wgt_6_470,
input [18:0] Wgt_6_471,
input [18:0] Wgt_6_472,
input [18:0] Wgt_6_473,
input [18:0] Wgt_6_474,
input [18:0] Wgt_6_475,
input [18:0] Wgt_6_476,
input [18:0] Wgt_6_477,
input [18:0] Wgt_6_478,
input [18:0] Wgt_6_479,
input [18:0] Wgt_6_480,
input [18:0] Wgt_6_481,
input [18:0] Wgt_6_482,
input [18:0] Wgt_6_483,
input [18:0] Wgt_6_484,
input [18:0] Wgt_6_485,
input [18:0] Wgt_6_486,
input [18:0] Wgt_6_487,
input [18:0] Wgt_6_488,
input [18:0] Wgt_6_489,
input [18:0] Wgt_6_490,
input [18:0] Wgt_6_491,
input [18:0] Wgt_6_492,
input [18:0] Wgt_6_493,
input [18:0] Wgt_6_494,
input [18:0] Wgt_6_495,
input [18:0] Wgt_6_496,
input [18:0] Wgt_6_497,
input [18:0] Wgt_6_498,
input [18:0] Wgt_6_499,
input [18:0] Wgt_6_500,
input [18:0] Wgt_6_501,
input [18:0] Wgt_6_502,
input [18:0] Wgt_6_503,
input [18:0] Wgt_6_504,
input [18:0] Wgt_6_505,
input [18:0] Wgt_6_506,
input [18:0] Wgt_6_507,
input [18:0] Wgt_6_508,
input [18:0] Wgt_6_509,
input [18:0] Wgt_6_510,
input [18:0] Wgt_6_511,
input [18:0] Wgt_6_512,
input [18:0] Wgt_6_513,
input [18:0] Wgt_6_514,
input [18:0] Wgt_6_515,
input [18:0] Wgt_6_516,
input [18:0] Wgt_6_517,
input [18:0] Wgt_6_518,
input [18:0] Wgt_6_519,
input [18:0] Wgt_6_520,
input [18:0] Wgt_6_521,
input [18:0] Wgt_6_522,
input [18:0] Wgt_6_523,
input [18:0] Wgt_6_524,
input [18:0] Wgt_6_525,
input [18:0] Wgt_6_526,
input [18:0] Wgt_6_527,
input [18:0] Wgt_6_528,
input [18:0] Wgt_6_529,
input [18:0] Wgt_6_530,
input [18:0] Wgt_6_531,
input [18:0] Wgt_6_532,
input [18:0] Wgt_6_533,
input [18:0] Wgt_6_534,
input [18:0] Wgt_6_535,
input [18:0] Wgt_6_536,
input [18:0] Wgt_6_537,
input [18:0] Wgt_6_538,
input [18:0] Wgt_6_539,
input [18:0] Wgt_6_540,
input [18:0] Wgt_6_541,
input [18:0] Wgt_6_542,
input [18:0] Wgt_6_543,
input [18:0] Wgt_6_544,
input [18:0] Wgt_6_545,
input [18:0] Wgt_6_546,
input [18:0] Wgt_6_547,
input [18:0] Wgt_6_548,
input [18:0] Wgt_6_549,
input [18:0] Wgt_6_550,
input [18:0] Wgt_6_551,
input [18:0] Wgt_6_552,
input [18:0] Wgt_6_553,
input [18:0] Wgt_6_554,
input [18:0] Wgt_6_555,
input [18:0] Wgt_6_556,
input [18:0] Wgt_6_557,
input [18:0] Wgt_6_558,
input [18:0] Wgt_6_559,
input [18:0] Wgt_6_560,
input [18:0] Wgt_6_561,
input [18:0] Wgt_6_562,
input [18:0] Wgt_6_563,
input [18:0] Wgt_6_564,
input [18:0] Wgt_6_565,
input [18:0] Wgt_6_566,
input [18:0] Wgt_6_567,
input [18:0] Wgt_6_568,
input [18:0] Wgt_6_569,
input [18:0] Wgt_6_570,
input [18:0] Wgt_6_571,
input [18:0] Wgt_6_572,
input [18:0] Wgt_6_573,
input [18:0] Wgt_6_574,
input [18:0] Wgt_6_575,
input [18:0] Wgt_6_576,
input [18:0] Wgt_6_577,
input [18:0] Wgt_6_578,
input [18:0] Wgt_6_579,
input [18:0] Wgt_6_580,
input [18:0] Wgt_6_581,
input [18:0] Wgt_6_582,
input [18:0] Wgt_6_583,
input [18:0] Wgt_6_584,
input [18:0] Wgt_6_585,
input [18:0] Wgt_6_586,
input [18:0] Wgt_6_587,
input [18:0] Wgt_6_588,
input [18:0] Wgt_6_589,
input [18:0] Wgt_6_590,
input [18:0] Wgt_6_591,
input [18:0] Wgt_6_592,
input [18:0] Wgt_6_593,
input [18:0] Wgt_6_594,
input [18:0] Wgt_6_595,
input [18:0] Wgt_6_596,
input [18:0] Wgt_6_597,
input [18:0] Wgt_6_598,
input [18:0] Wgt_6_599,
input [18:0] Wgt_6_600,
input [18:0] Wgt_6_601,
input [18:0] Wgt_6_602,
input [18:0] Wgt_6_603,
input [18:0] Wgt_6_604,
input [18:0] Wgt_6_605,
input [18:0] Wgt_6_606,
input [18:0] Wgt_6_607,
input [18:0] Wgt_6_608,
input [18:0] Wgt_6_609,
input [18:0] Wgt_6_610,
input [18:0] Wgt_6_611,
input [18:0] Wgt_6_612,
input [18:0] Wgt_6_613,
input [18:0] Wgt_6_614,
input [18:0] Wgt_6_615,
input [18:0] Wgt_6_616,
input [18:0] Wgt_6_617,
input [18:0] Wgt_6_618,
input [18:0] Wgt_6_619,
input [18:0] Wgt_6_620,
input [18:0] Wgt_6_621,
input [18:0] Wgt_6_622,
input [18:0] Wgt_6_623,
input [18:0] Wgt_6_624,
input [18:0] Wgt_6_625,
input [18:0] Wgt_6_626,
input [18:0] Wgt_6_627,
input [18:0] Wgt_6_628,
input [18:0] Wgt_6_629,
input [18:0] Wgt_6_630,
input [18:0] Wgt_6_631,
input [18:0] Wgt_6_632,
input [18:0] Wgt_6_633,
input [18:0] Wgt_6_634,
input [18:0] Wgt_6_635,
input [18:0] Wgt_6_636,
input [18:0] Wgt_6_637,
input [18:0] Wgt_6_638,
input [18:0] Wgt_6_639,
input [18:0] Wgt_6_640,
input [18:0] Wgt_6_641,
input [18:0] Wgt_6_642,
input [18:0] Wgt_6_643,
input [18:0] Wgt_6_644,
input [18:0] Wgt_6_645,
input [18:0] Wgt_6_646,
input [18:0] Wgt_6_647,
input [18:0] Wgt_6_648,
input [18:0] Wgt_6_649,
input [18:0] Wgt_6_650,
input [18:0] Wgt_6_651,
input [18:0] Wgt_6_652,
input [18:0] Wgt_6_653,
input [18:0] Wgt_6_654,
input [18:0] Wgt_6_655,
input [18:0] Wgt_6_656,
input [18:0] Wgt_6_657,
input [18:0] Wgt_6_658,
input [18:0] Wgt_6_659,
input [18:0] Wgt_6_660,
input [18:0] Wgt_6_661,
input [18:0] Wgt_6_662,
input [18:0] Wgt_6_663,
input [18:0] Wgt_6_664,
input [18:0] Wgt_6_665,
input [18:0] Wgt_6_666,
input [18:0] Wgt_6_667,
input [18:0] Wgt_6_668,
input [18:0] Wgt_6_669,
input [18:0] Wgt_6_670,
input [18:0] Wgt_6_671,
input [18:0] Wgt_6_672,
input [18:0] Wgt_6_673,
input [18:0] Wgt_6_674,
input [18:0] Wgt_6_675,
input [18:0] Wgt_6_676,
input [18:0] Wgt_6_677,
input [18:0] Wgt_6_678,
input [18:0] Wgt_6_679,
input [18:0] Wgt_6_680,
input [18:0] Wgt_6_681,
input [18:0] Wgt_6_682,
input [18:0] Wgt_6_683,
input [18:0] Wgt_6_684,
input [18:0] Wgt_6_685,
input [18:0] Wgt_6_686,
input [18:0] Wgt_6_687,
input [18:0] Wgt_6_688,
input [18:0] Wgt_6_689,
input [18:0] Wgt_6_690,
input [18:0] Wgt_6_691,
input [18:0] Wgt_6_692,
input [18:0] Wgt_6_693,
input [18:0] Wgt_6_694,
input [18:0] Wgt_6_695,
input [18:0] Wgt_6_696,
input [18:0] Wgt_6_697,
input [18:0] Wgt_6_698,
input [18:0] Wgt_6_699,
input [18:0] Wgt_6_700,
input [18:0] Wgt_6_701,
input [18:0] Wgt_6_702,
input [18:0] Wgt_6_703,
input [18:0] Wgt_6_704,
input [18:0] Wgt_6_705,
input [18:0] Wgt_6_706,
input [18:0] Wgt_6_707,
input [18:0] Wgt_6_708,
input [18:0] Wgt_6_709,
input [18:0] Wgt_6_710,
input [18:0] Wgt_6_711,
input [18:0] Wgt_6_712,
input [18:0] Wgt_6_713,
input [18:0] Wgt_6_714,
input [18:0] Wgt_6_715,
input [18:0] Wgt_6_716,
input [18:0] Wgt_6_717,
input [18:0] Wgt_6_718,
input [18:0] Wgt_6_719,
input [18:0] Wgt_6_720,
input [18:0] Wgt_6_721,
input [18:0] Wgt_6_722,
input [18:0] Wgt_6_723,
input [18:0] Wgt_6_724,
input [18:0] Wgt_6_725,
input [18:0] Wgt_6_726,
input [18:0] Wgt_6_727,
input [18:0] Wgt_6_728,
input [18:0] Wgt_6_729,
input [18:0] Wgt_6_730,
input [18:0] Wgt_6_731,
input [18:0] Wgt_6_732,
input [18:0] Wgt_6_733,
input [18:0] Wgt_6_734,
input [18:0] Wgt_6_735,
input [18:0] Wgt_6_736,
input [18:0] Wgt_6_737,
input [18:0] Wgt_6_738,
input [18:0] Wgt_6_739,
input [18:0] Wgt_6_740,
input [18:0] Wgt_6_741,
input [18:0] Wgt_6_742,
input [18:0] Wgt_6_743,
input [18:0] Wgt_6_744,
input [18:0] Wgt_6_745,
input [18:0] Wgt_6_746,
input [18:0] Wgt_6_747,
input [18:0] Wgt_6_748,
input [18:0] Wgt_6_749,
input [18:0] Wgt_6_750,
input [18:0] Wgt_6_751,
input [18:0] Wgt_6_752,
input [18:0] Wgt_6_753,
input [18:0] Wgt_6_754,
input [18:0] Wgt_6_755,
input [18:0] Wgt_6_756,
input [18:0] Wgt_6_757,
input [18:0] Wgt_6_758,
input [18:0] Wgt_6_759,
input [18:0] Wgt_6_760,
input [18:0] Wgt_6_761,
input [18:0] Wgt_6_762,
input [18:0] Wgt_6_763,
input [18:0] Wgt_6_764,
input [18:0] Wgt_6_765,
input [18:0] Wgt_6_766,
input [18:0] Wgt_6_767,
input [18:0] Wgt_6_768,
input [18:0] Wgt_6_769,
input [18:0] Wgt_6_770,
input [18:0] Wgt_6_771,
input [18:0] Wgt_6_772,
input [18:0] Wgt_6_773,
input [18:0] Wgt_6_774,
input [18:0] Wgt_6_775,
input [18:0] Wgt_6_776,
input [18:0] Wgt_6_777,
input [18:0] Wgt_6_778,
input [18:0] Wgt_6_779,
input [18:0] Wgt_6_780,
input [18:0] Wgt_6_781,
input [18:0] Wgt_6_782,
input [18:0] Wgt_6_783,
input [18:0] Wgt_6_784,
input [18:0] Wgt_7_0,
input [18:0] Wgt_7_1,
input [18:0] Wgt_7_2,
input [18:0] Wgt_7_3,
input [18:0] Wgt_7_4,
input [18:0] Wgt_7_5,
input [18:0] Wgt_7_6,
input [18:0] Wgt_7_7,
input [18:0] Wgt_7_8,
input [18:0] Wgt_7_9,
input [18:0] Wgt_7_10,
input [18:0] Wgt_7_11,
input [18:0] Wgt_7_12,
input [18:0] Wgt_7_13,
input [18:0] Wgt_7_14,
input [18:0] Wgt_7_15,
input [18:0] Wgt_7_16,
input [18:0] Wgt_7_17,
input [18:0] Wgt_7_18,
input [18:0] Wgt_7_19,
input [18:0] Wgt_7_20,
input [18:0] Wgt_7_21,
input [18:0] Wgt_7_22,
input [18:0] Wgt_7_23,
input [18:0] Wgt_7_24,
input [18:0] Wgt_7_25,
input [18:0] Wgt_7_26,
input [18:0] Wgt_7_27,
input [18:0] Wgt_7_28,
input [18:0] Wgt_7_29,
input [18:0] Wgt_7_30,
input [18:0] Wgt_7_31,
input [18:0] Wgt_7_32,
input [18:0] Wgt_7_33,
input [18:0] Wgt_7_34,
input [18:0] Wgt_7_35,
input [18:0] Wgt_7_36,
input [18:0] Wgt_7_37,
input [18:0] Wgt_7_38,
input [18:0] Wgt_7_39,
input [18:0] Wgt_7_40,
input [18:0] Wgt_7_41,
input [18:0] Wgt_7_42,
input [18:0] Wgt_7_43,
input [18:0] Wgt_7_44,
input [18:0] Wgt_7_45,
input [18:0] Wgt_7_46,
input [18:0] Wgt_7_47,
input [18:0] Wgt_7_48,
input [18:0] Wgt_7_49,
input [18:0] Wgt_7_50,
input [18:0] Wgt_7_51,
input [18:0] Wgt_7_52,
input [18:0] Wgt_7_53,
input [18:0] Wgt_7_54,
input [18:0] Wgt_7_55,
input [18:0] Wgt_7_56,
input [18:0] Wgt_7_57,
input [18:0] Wgt_7_58,
input [18:0] Wgt_7_59,
input [18:0] Wgt_7_60,
input [18:0] Wgt_7_61,
input [18:0] Wgt_7_62,
input [18:0] Wgt_7_63,
input [18:0] Wgt_7_64,
input [18:0] Wgt_7_65,
input [18:0] Wgt_7_66,
input [18:0] Wgt_7_67,
input [18:0] Wgt_7_68,
input [18:0] Wgt_7_69,
input [18:0] Wgt_7_70,
input [18:0] Wgt_7_71,
input [18:0] Wgt_7_72,
input [18:0] Wgt_7_73,
input [18:0] Wgt_7_74,
input [18:0] Wgt_7_75,
input [18:0] Wgt_7_76,
input [18:0] Wgt_7_77,
input [18:0] Wgt_7_78,
input [18:0] Wgt_7_79,
input [18:0] Wgt_7_80,
input [18:0] Wgt_7_81,
input [18:0] Wgt_7_82,
input [18:0] Wgt_7_83,
input [18:0] Wgt_7_84,
input [18:0] Wgt_7_85,
input [18:0] Wgt_7_86,
input [18:0] Wgt_7_87,
input [18:0] Wgt_7_88,
input [18:0] Wgt_7_89,
input [18:0] Wgt_7_90,
input [18:0] Wgt_7_91,
input [18:0] Wgt_7_92,
input [18:0] Wgt_7_93,
input [18:0] Wgt_7_94,
input [18:0] Wgt_7_95,
input [18:0] Wgt_7_96,
input [18:0] Wgt_7_97,
input [18:0] Wgt_7_98,
input [18:0] Wgt_7_99,
input [18:0] Wgt_7_100,
input [18:0] Wgt_7_101,
input [18:0] Wgt_7_102,
input [18:0] Wgt_7_103,
input [18:0] Wgt_7_104,
input [18:0] Wgt_7_105,
input [18:0] Wgt_7_106,
input [18:0] Wgt_7_107,
input [18:0] Wgt_7_108,
input [18:0] Wgt_7_109,
input [18:0] Wgt_7_110,
input [18:0] Wgt_7_111,
input [18:0] Wgt_7_112,
input [18:0] Wgt_7_113,
input [18:0] Wgt_7_114,
input [18:0] Wgt_7_115,
input [18:0] Wgt_7_116,
input [18:0] Wgt_7_117,
input [18:0] Wgt_7_118,
input [18:0] Wgt_7_119,
input [18:0] Wgt_7_120,
input [18:0] Wgt_7_121,
input [18:0] Wgt_7_122,
input [18:0] Wgt_7_123,
input [18:0] Wgt_7_124,
input [18:0] Wgt_7_125,
input [18:0] Wgt_7_126,
input [18:0] Wgt_7_127,
input [18:0] Wgt_7_128,
input [18:0] Wgt_7_129,
input [18:0] Wgt_7_130,
input [18:0] Wgt_7_131,
input [18:0] Wgt_7_132,
input [18:0] Wgt_7_133,
input [18:0] Wgt_7_134,
input [18:0] Wgt_7_135,
input [18:0] Wgt_7_136,
input [18:0] Wgt_7_137,
input [18:0] Wgt_7_138,
input [18:0] Wgt_7_139,
input [18:0] Wgt_7_140,
input [18:0] Wgt_7_141,
input [18:0] Wgt_7_142,
input [18:0] Wgt_7_143,
input [18:0] Wgt_7_144,
input [18:0] Wgt_7_145,
input [18:0] Wgt_7_146,
input [18:0] Wgt_7_147,
input [18:0] Wgt_7_148,
input [18:0] Wgt_7_149,
input [18:0] Wgt_7_150,
input [18:0] Wgt_7_151,
input [18:0] Wgt_7_152,
input [18:0] Wgt_7_153,
input [18:0] Wgt_7_154,
input [18:0] Wgt_7_155,
input [18:0] Wgt_7_156,
input [18:0] Wgt_7_157,
input [18:0] Wgt_7_158,
input [18:0] Wgt_7_159,
input [18:0] Wgt_7_160,
input [18:0] Wgt_7_161,
input [18:0] Wgt_7_162,
input [18:0] Wgt_7_163,
input [18:0] Wgt_7_164,
input [18:0] Wgt_7_165,
input [18:0] Wgt_7_166,
input [18:0] Wgt_7_167,
input [18:0] Wgt_7_168,
input [18:0] Wgt_7_169,
input [18:0] Wgt_7_170,
input [18:0] Wgt_7_171,
input [18:0] Wgt_7_172,
input [18:0] Wgt_7_173,
input [18:0] Wgt_7_174,
input [18:0] Wgt_7_175,
input [18:0] Wgt_7_176,
input [18:0] Wgt_7_177,
input [18:0] Wgt_7_178,
input [18:0] Wgt_7_179,
input [18:0] Wgt_7_180,
input [18:0] Wgt_7_181,
input [18:0] Wgt_7_182,
input [18:0] Wgt_7_183,
input [18:0] Wgt_7_184,
input [18:0] Wgt_7_185,
input [18:0] Wgt_7_186,
input [18:0] Wgt_7_187,
input [18:0] Wgt_7_188,
input [18:0] Wgt_7_189,
input [18:0] Wgt_7_190,
input [18:0] Wgt_7_191,
input [18:0] Wgt_7_192,
input [18:0] Wgt_7_193,
input [18:0] Wgt_7_194,
input [18:0] Wgt_7_195,
input [18:0] Wgt_7_196,
input [18:0] Wgt_7_197,
input [18:0] Wgt_7_198,
input [18:0] Wgt_7_199,
input [18:0] Wgt_7_200,
input [18:0] Wgt_7_201,
input [18:0] Wgt_7_202,
input [18:0] Wgt_7_203,
input [18:0] Wgt_7_204,
input [18:0] Wgt_7_205,
input [18:0] Wgt_7_206,
input [18:0] Wgt_7_207,
input [18:0] Wgt_7_208,
input [18:0] Wgt_7_209,
input [18:0] Wgt_7_210,
input [18:0] Wgt_7_211,
input [18:0] Wgt_7_212,
input [18:0] Wgt_7_213,
input [18:0] Wgt_7_214,
input [18:0] Wgt_7_215,
input [18:0] Wgt_7_216,
input [18:0] Wgt_7_217,
input [18:0] Wgt_7_218,
input [18:0] Wgt_7_219,
input [18:0] Wgt_7_220,
input [18:0] Wgt_7_221,
input [18:0] Wgt_7_222,
input [18:0] Wgt_7_223,
input [18:0] Wgt_7_224,
input [18:0] Wgt_7_225,
input [18:0] Wgt_7_226,
input [18:0] Wgt_7_227,
input [18:0] Wgt_7_228,
input [18:0] Wgt_7_229,
input [18:0] Wgt_7_230,
input [18:0] Wgt_7_231,
input [18:0] Wgt_7_232,
input [18:0] Wgt_7_233,
input [18:0] Wgt_7_234,
input [18:0] Wgt_7_235,
input [18:0] Wgt_7_236,
input [18:0] Wgt_7_237,
input [18:0] Wgt_7_238,
input [18:0] Wgt_7_239,
input [18:0] Wgt_7_240,
input [18:0] Wgt_7_241,
input [18:0] Wgt_7_242,
input [18:0] Wgt_7_243,
input [18:0] Wgt_7_244,
input [18:0] Wgt_7_245,
input [18:0] Wgt_7_246,
input [18:0] Wgt_7_247,
input [18:0] Wgt_7_248,
input [18:0] Wgt_7_249,
input [18:0] Wgt_7_250,
input [18:0] Wgt_7_251,
input [18:0] Wgt_7_252,
input [18:0] Wgt_7_253,
input [18:0] Wgt_7_254,
input [18:0] Wgt_7_255,
input [18:0] Wgt_7_256,
input [18:0] Wgt_7_257,
input [18:0] Wgt_7_258,
input [18:0] Wgt_7_259,
input [18:0] Wgt_7_260,
input [18:0] Wgt_7_261,
input [18:0] Wgt_7_262,
input [18:0] Wgt_7_263,
input [18:0] Wgt_7_264,
input [18:0] Wgt_7_265,
input [18:0] Wgt_7_266,
input [18:0] Wgt_7_267,
input [18:0] Wgt_7_268,
input [18:0] Wgt_7_269,
input [18:0] Wgt_7_270,
input [18:0] Wgt_7_271,
input [18:0] Wgt_7_272,
input [18:0] Wgt_7_273,
input [18:0] Wgt_7_274,
input [18:0] Wgt_7_275,
input [18:0] Wgt_7_276,
input [18:0] Wgt_7_277,
input [18:0] Wgt_7_278,
input [18:0] Wgt_7_279,
input [18:0] Wgt_7_280,
input [18:0] Wgt_7_281,
input [18:0] Wgt_7_282,
input [18:0] Wgt_7_283,
input [18:0] Wgt_7_284,
input [18:0] Wgt_7_285,
input [18:0] Wgt_7_286,
input [18:0] Wgt_7_287,
input [18:0] Wgt_7_288,
input [18:0] Wgt_7_289,
input [18:0] Wgt_7_290,
input [18:0] Wgt_7_291,
input [18:0] Wgt_7_292,
input [18:0] Wgt_7_293,
input [18:0] Wgt_7_294,
input [18:0] Wgt_7_295,
input [18:0] Wgt_7_296,
input [18:0] Wgt_7_297,
input [18:0] Wgt_7_298,
input [18:0] Wgt_7_299,
input [18:0] Wgt_7_300,
input [18:0] Wgt_7_301,
input [18:0] Wgt_7_302,
input [18:0] Wgt_7_303,
input [18:0] Wgt_7_304,
input [18:0] Wgt_7_305,
input [18:0] Wgt_7_306,
input [18:0] Wgt_7_307,
input [18:0] Wgt_7_308,
input [18:0] Wgt_7_309,
input [18:0] Wgt_7_310,
input [18:0] Wgt_7_311,
input [18:0] Wgt_7_312,
input [18:0] Wgt_7_313,
input [18:0] Wgt_7_314,
input [18:0] Wgt_7_315,
input [18:0] Wgt_7_316,
input [18:0] Wgt_7_317,
input [18:0] Wgt_7_318,
input [18:0] Wgt_7_319,
input [18:0] Wgt_7_320,
input [18:0] Wgt_7_321,
input [18:0] Wgt_7_322,
input [18:0] Wgt_7_323,
input [18:0] Wgt_7_324,
input [18:0] Wgt_7_325,
input [18:0] Wgt_7_326,
input [18:0] Wgt_7_327,
input [18:0] Wgt_7_328,
input [18:0] Wgt_7_329,
input [18:0] Wgt_7_330,
input [18:0] Wgt_7_331,
input [18:0] Wgt_7_332,
input [18:0] Wgt_7_333,
input [18:0] Wgt_7_334,
input [18:0] Wgt_7_335,
input [18:0] Wgt_7_336,
input [18:0] Wgt_7_337,
input [18:0] Wgt_7_338,
input [18:0] Wgt_7_339,
input [18:0] Wgt_7_340,
input [18:0] Wgt_7_341,
input [18:0] Wgt_7_342,
input [18:0] Wgt_7_343,
input [18:0] Wgt_7_344,
input [18:0] Wgt_7_345,
input [18:0] Wgt_7_346,
input [18:0] Wgt_7_347,
input [18:0] Wgt_7_348,
input [18:0] Wgt_7_349,
input [18:0] Wgt_7_350,
input [18:0] Wgt_7_351,
input [18:0] Wgt_7_352,
input [18:0] Wgt_7_353,
input [18:0] Wgt_7_354,
input [18:0] Wgt_7_355,
input [18:0] Wgt_7_356,
input [18:0] Wgt_7_357,
input [18:0] Wgt_7_358,
input [18:0] Wgt_7_359,
input [18:0] Wgt_7_360,
input [18:0] Wgt_7_361,
input [18:0] Wgt_7_362,
input [18:0] Wgt_7_363,
input [18:0] Wgt_7_364,
input [18:0] Wgt_7_365,
input [18:0] Wgt_7_366,
input [18:0] Wgt_7_367,
input [18:0] Wgt_7_368,
input [18:0] Wgt_7_369,
input [18:0] Wgt_7_370,
input [18:0] Wgt_7_371,
input [18:0] Wgt_7_372,
input [18:0] Wgt_7_373,
input [18:0] Wgt_7_374,
input [18:0] Wgt_7_375,
input [18:0] Wgt_7_376,
input [18:0] Wgt_7_377,
input [18:0] Wgt_7_378,
input [18:0] Wgt_7_379,
input [18:0] Wgt_7_380,
input [18:0] Wgt_7_381,
input [18:0] Wgt_7_382,
input [18:0] Wgt_7_383,
input [18:0] Wgt_7_384,
input [18:0] Wgt_7_385,
input [18:0] Wgt_7_386,
input [18:0] Wgt_7_387,
input [18:0] Wgt_7_388,
input [18:0] Wgt_7_389,
input [18:0] Wgt_7_390,
input [18:0] Wgt_7_391,
input [18:0] Wgt_7_392,
input [18:0] Wgt_7_393,
input [18:0] Wgt_7_394,
input [18:0] Wgt_7_395,
input [18:0] Wgt_7_396,
input [18:0] Wgt_7_397,
input [18:0] Wgt_7_398,
input [18:0] Wgt_7_399,
input [18:0] Wgt_7_400,
input [18:0] Wgt_7_401,
input [18:0] Wgt_7_402,
input [18:0] Wgt_7_403,
input [18:0] Wgt_7_404,
input [18:0] Wgt_7_405,
input [18:0] Wgt_7_406,
input [18:0] Wgt_7_407,
input [18:0] Wgt_7_408,
input [18:0] Wgt_7_409,
input [18:0] Wgt_7_410,
input [18:0] Wgt_7_411,
input [18:0] Wgt_7_412,
input [18:0] Wgt_7_413,
input [18:0] Wgt_7_414,
input [18:0] Wgt_7_415,
input [18:0] Wgt_7_416,
input [18:0] Wgt_7_417,
input [18:0] Wgt_7_418,
input [18:0] Wgt_7_419,
input [18:0] Wgt_7_420,
input [18:0] Wgt_7_421,
input [18:0] Wgt_7_422,
input [18:0] Wgt_7_423,
input [18:0] Wgt_7_424,
input [18:0] Wgt_7_425,
input [18:0] Wgt_7_426,
input [18:0] Wgt_7_427,
input [18:0] Wgt_7_428,
input [18:0] Wgt_7_429,
input [18:0] Wgt_7_430,
input [18:0] Wgt_7_431,
input [18:0] Wgt_7_432,
input [18:0] Wgt_7_433,
input [18:0] Wgt_7_434,
input [18:0] Wgt_7_435,
input [18:0] Wgt_7_436,
input [18:0] Wgt_7_437,
input [18:0] Wgt_7_438,
input [18:0] Wgt_7_439,
input [18:0] Wgt_7_440,
input [18:0] Wgt_7_441,
input [18:0] Wgt_7_442,
input [18:0] Wgt_7_443,
input [18:0] Wgt_7_444,
input [18:0] Wgt_7_445,
input [18:0] Wgt_7_446,
input [18:0] Wgt_7_447,
input [18:0] Wgt_7_448,
input [18:0] Wgt_7_449,
input [18:0] Wgt_7_450,
input [18:0] Wgt_7_451,
input [18:0] Wgt_7_452,
input [18:0] Wgt_7_453,
input [18:0] Wgt_7_454,
input [18:0] Wgt_7_455,
input [18:0] Wgt_7_456,
input [18:0] Wgt_7_457,
input [18:0] Wgt_7_458,
input [18:0] Wgt_7_459,
input [18:0] Wgt_7_460,
input [18:0] Wgt_7_461,
input [18:0] Wgt_7_462,
input [18:0] Wgt_7_463,
input [18:0] Wgt_7_464,
input [18:0] Wgt_7_465,
input [18:0] Wgt_7_466,
input [18:0] Wgt_7_467,
input [18:0] Wgt_7_468,
input [18:0] Wgt_7_469,
input [18:0] Wgt_7_470,
input [18:0] Wgt_7_471,
input [18:0] Wgt_7_472,
input [18:0] Wgt_7_473,
input [18:0] Wgt_7_474,
input [18:0] Wgt_7_475,
input [18:0] Wgt_7_476,
input [18:0] Wgt_7_477,
input [18:0] Wgt_7_478,
input [18:0] Wgt_7_479,
input [18:0] Wgt_7_480,
input [18:0] Wgt_7_481,
input [18:0] Wgt_7_482,
input [18:0] Wgt_7_483,
input [18:0] Wgt_7_484,
input [18:0] Wgt_7_485,
input [18:0] Wgt_7_486,
input [18:0] Wgt_7_487,
input [18:0] Wgt_7_488,
input [18:0] Wgt_7_489,
input [18:0] Wgt_7_490,
input [18:0] Wgt_7_491,
input [18:0] Wgt_7_492,
input [18:0] Wgt_7_493,
input [18:0] Wgt_7_494,
input [18:0] Wgt_7_495,
input [18:0] Wgt_7_496,
input [18:0] Wgt_7_497,
input [18:0] Wgt_7_498,
input [18:0] Wgt_7_499,
input [18:0] Wgt_7_500,
input [18:0] Wgt_7_501,
input [18:0] Wgt_7_502,
input [18:0] Wgt_7_503,
input [18:0] Wgt_7_504,
input [18:0] Wgt_7_505,
input [18:0] Wgt_7_506,
input [18:0] Wgt_7_507,
input [18:0] Wgt_7_508,
input [18:0] Wgt_7_509,
input [18:0] Wgt_7_510,
input [18:0] Wgt_7_511,
input [18:0] Wgt_7_512,
input [18:0] Wgt_7_513,
input [18:0] Wgt_7_514,
input [18:0] Wgt_7_515,
input [18:0] Wgt_7_516,
input [18:0] Wgt_7_517,
input [18:0] Wgt_7_518,
input [18:0] Wgt_7_519,
input [18:0] Wgt_7_520,
input [18:0] Wgt_7_521,
input [18:0] Wgt_7_522,
input [18:0] Wgt_7_523,
input [18:0] Wgt_7_524,
input [18:0] Wgt_7_525,
input [18:0] Wgt_7_526,
input [18:0] Wgt_7_527,
input [18:0] Wgt_7_528,
input [18:0] Wgt_7_529,
input [18:0] Wgt_7_530,
input [18:0] Wgt_7_531,
input [18:0] Wgt_7_532,
input [18:0] Wgt_7_533,
input [18:0] Wgt_7_534,
input [18:0] Wgt_7_535,
input [18:0] Wgt_7_536,
input [18:0] Wgt_7_537,
input [18:0] Wgt_7_538,
input [18:0] Wgt_7_539,
input [18:0] Wgt_7_540,
input [18:0] Wgt_7_541,
input [18:0] Wgt_7_542,
input [18:0] Wgt_7_543,
input [18:0] Wgt_7_544,
input [18:0] Wgt_7_545,
input [18:0] Wgt_7_546,
input [18:0] Wgt_7_547,
input [18:0] Wgt_7_548,
input [18:0] Wgt_7_549,
input [18:0] Wgt_7_550,
input [18:0] Wgt_7_551,
input [18:0] Wgt_7_552,
input [18:0] Wgt_7_553,
input [18:0] Wgt_7_554,
input [18:0] Wgt_7_555,
input [18:0] Wgt_7_556,
input [18:0] Wgt_7_557,
input [18:0] Wgt_7_558,
input [18:0] Wgt_7_559,
input [18:0] Wgt_7_560,
input [18:0] Wgt_7_561,
input [18:0] Wgt_7_562,
input [18:0] Wgt_7_563,
input [18:0] Wgt_7_564,
input [18:0] Wgt_7_565,
input [18:0] Wgt_7_566,
input [18:0] Wgt_7_567,
input [18:0] Wgt_7_568,
input [18:0] Wgt_7_569,
input [18:0] Wgt_7_570,
input [18:0] Wgt_7_571,
input [18:0] Wgt_7_572,
input [18:0] Wgt_7_573,
input [18:0] Wgt_7_574,
input [18:0] Wgt_7_575,
input [18:0] Wgt_7_576,
input [18:0] Wgt_7_577,
input [18:0] Wgt_7_578,
input [18:0] Wgt_7_579,
input [18:0] Wgt_7_580,
input [18:0] Wgt_7_581,
input [18:0] Wgt_7_582,
input [18:0] Wgt_7_583,
input [18:0] Wgt_7_584,
input [18:0] Wgt_7_585,
input [18:0] Wgt_7_586,
input [18:0] Wgt_7_587,
input [18:0] Wgt_7_588,
input [18:0] Wgt_7_589,
input [18:0] Wgt_7_590,
input [18:0] Wgt_7_591,
input [18:0] Wgt_7_592,
input [18:0] Wgt_7_593,
input [18:0] Wgt_7_594,
input [18:0] Wgt_7_595,
input [18:0] Wgt_7_596,
input [18:0] Wgt_7_597,
input [18:0] Wgt_7_598,
input [18:0] Wgt_7_599,
input [18:0] Wgt_7_600,
input [18:0] Wgt_7_601,
input [18:0] Wgt_7_602,
input [18:0] Wgt_7_603,
input [18:0] Wgt_7_604,
input [18:0] Wgt_7_605,
input [18:0] Wgt_7_606,
input [18:0] Wgt_7_607,
input [18:0] Wgt_7_608,
input [18:0] Wgt_7_609,
input [18:0] Wgt_7_610,
input [18:0] Wgt_7_611,
input [18:0] Wgt_7_612,
input [18:0] Wgt_7_613,
input [18:0] Wgt_7_614,
input [18:0] Wgt_7_615,
input [18:0] Wgt_7_616,
input [18:0] Wgt_7_617,
input [18:0] Wgt_7_618,
input [18:0] Wgt_7_619,
input [18:0] Wgt_7_620,
input [18:0] Wgt_7_621,
input [18:0] Wgt_7_622,
input [18:0] Wgt_7_623,
input [18:0] Wgt_7_624,
input [18:0] Wgt_7_625,
input [18:0] Wgt_7_626,
input [18:0] Wgt_7_627,
input [18:0] Wgt_7_628,
input [18:0] Wgt_7_629,
input [18:0] Wgt_7_630,
input [18:0] Wgt_7_631,
input [18:0] Wgt_7_632,
input [18:0] Wgt_7_633,
input [18:0] Wgt_7_634,
input [18:0] Wgt_7_635,
input [18:0] Wgt_7_636,
input [18:0] Wgt_7_637,
input [18:0] Wgt_7_638,
input [18:0] Wgt_7_639,
input [18:0] Wgt_7_640,
input [18:0] Wgt_7_641,
input [18:0] Wgt_7_642,
input [18:0] Wgt_7_643,
input [18:0] Wgt_7_644,
input [18:0] Wgt_7_645,
input [18:0] Wgt_7_646,
input [18:0] Wgt_7_647,
input [18:0] Wgt_7_648,
input [18:0] Wgt_7_649,
input [18:0] Wgt_7_650,
input [18:0] Wgt_7_651,
input [18:0] Wgt_7_652,
input [18:0] Wgt_7_653,
input [18:0] Wgt_7_654,
input [18:0] Wgt_7_655,
input [18:0] Wgt_7_656,
input [18:0] Wgt_7_657,
input [18:0] Wgt_7_658,
input [18:0] Wgt_7_659,
input [18:0] Wgt_7_660,
input [18:0] Wgt_7_661,
input [18:0] Wgt_7_662,
input [18:0] Wgt_7_663,
input [18:0] Wgt_7_664,
input [18:0] Wgt_7_665,
input [18:0] Wgt_7_666,
input [18:0] Wgt_7_667,
input [18:0] Wgt_7_668,
input [18:0] Wgt_7_669,
input [18:0] Wgt_7_670,
input [18:0] Wgt_7_671,
input [18:0] Wgt_7_672,
input [18:0] Wgt_7_673,
input [18:0] Wgt_7_674,
input [18:0] Wgt_7_675,
input [18:0] Wgt_7_676,
input [18:0] Wgt_7_677,
input [18:0] Wgt_7_678,
input [18:0] Wgt_7_679,
input [18:0] Wgt_7_680,
input [18:0] Wgt_7_681,
input [18:0] Wgt_7_682,
input [18:0] Wgt_7_683,
input [18:0] Wgt_7_684,
input [18:0] Wgt_7_685,
input [18:0] Wgt_7_686,
input [18:0] Wgt_7_687,
input [18:0] Wgt_7_688,
input [18:0] Wgt_7_689,
input [18:0] Wgt_7_690,
input [18:0] Wgt_7_691,
input [18:0] Wgt_7_692,
input [18:0] Wgt_7_693,
input [18:0] Wgt_7_694,
input [18:0] Wgt_7_695,
input [18:0] Wgt_7_696,
input [18:0] Wgt_7_697,
input [18:0] Wgt_7_698,
input [18:0] Wgt_7_699,
input [18:0] Wgt_7_700,
input [18:0] Wgt_7_701,
input [18:0] Wgt_7_702,
input [18:0] Wgt_7_703,
input [18:0] Wgt_7_704,
input [18:0] Wgt_7_705,
input [18:0] Wgt_7_706,
input [18:0] Wgt_7_707,
input [18:0] Wgt_7_708,
input [18:0] Wgt_7_709,
input [18:0] Wgt_7_710,
input [18:0] Wgt_7_711,
input [18:0] Wgt_7_712,
input [18:0] Wgt_7_713,
input [18:0] Wgt_7_714,
input [18:0] Wgt_7_715,
input [18:0] Wgt_7_716,
input [18:0] Wgt_7_717,
input [18:0] Wgt_7_718,
input [18:0] Wgt_7_719,
input [18:0] Wgt_7_720,
input [18:0] Wgt_7_721,
input [18:0] Wgt_7_722,
input [18:0] Wgt_7_723,
input [18:0] Wgt_7_724,
input [18:0] Wgt_7_725,
input [18:0] Wgt_7_726,
input [18:0] Wgt_7_727,
input [18:0] Wgt_7_728,
input [18:0] Wgt_7_729,
input [18:0] Wgt_7_730,
input [18:0] Wgt_7_731,
input [18:0] Wgt_7_732,
input [18:0] Wgt_7_733,
input [18:0] Wgt_7_734,
input [18:0] Wgt_7_735,
input [18:0] Wgt_7_736,
input [18:0] Wgt_7_737,
input [18:0] Wgt_7_738,
input [18:0] Wgt_7_739,
input [18:0] Wgt_7_740,
input [18:0] Wgt_7_741,
input [18:0] Wgt_7_742,
input [18:0] Wgt_7_743,
input [18:0] Wgt_7_744,
input [18:0] Wgt_7_745,
input [18:0] Wgt_7_746,
input [18:0] Wgt_7_747,
input [18:0] Wgt_7_748,
input [18:0] Wgt_7_749,
input [18:0] Wgt_7_750,
input [18:0] Wgt_7_751,
input [18:0] Wgt_7_752,
input [18:0] Wgt_7_753,
input [18:0] Wgt_7_754,
input [18:0] Wgt_7_755,
input [18:0] Wgt_7_756,
input [18:0] Wgt_7_757,
input [18:0] Wgt_7_758,
input [18:0] Wgt_7_759,
input [18:0] Wgt_7_760,
input [18:0] Wgt_7_761,
input [18:0] Wgt_7_762,
input [18:0] Wgt_7_763,
input [18:0] Wgt_7_764,
input [18:0] Wgt_7_765,
input [18:0] Wgt_7_766,
input [18:0] Wgt_7_767,
input [18:0] Wgt_7_768,
input [18:0] Wgt_7_769,
input [18:0] Wgt_7_770,
input [18:0] Wgt_7_771,
input [18:0] Wgt_7_772,
input [18:0] Wgt_7_773,
input [18:0] Wgt_7_774,
input [18:0] Wgt_7_775,
input [18:0] Wgt_7_776,
input [18:0] Wgt_7_777,
input [18:0] Wgt_7_778,
input [18:0] Wgt_7_779,
input [18:0] Wgt_7_780,
input [18:0] Wgt_7_781,
input [18:0] Wgt_7_782,
input [18:0] Wgt_7_783,
input [18:0] Wgt_7_784,
input [18:0] Wgt_8_0,
input [18:0] Wgt_8_1,
input [18:0] Wgt_8_2,
input [18:0] Wgt_8_3,
input [18:0] Wgt_8_4,
input [18:0] Wgt_8_5,
input [18:0] Wgt_8_6,
input [18:0] Wgt_8_7,
input [18:0] Wgt_8_8,
input [18:0] Wgt_8_9,
input [18:0] Wgt_8_10,
input [18:0] Wgt_8_11,
input [18:0] Wgt_8_12,
input [18:0] Wgt_8_13,
input [18:0] Wgt_8_14,
input [18:0] Wgt_8_15,
input [18:0] Wgt_8_16,
input [18:0] Wgt_8_17,
input [18:0] Wgt_8_18,
input [18:0] Wgt_8_19,
input [18:0] Wgt_8_20,
input [18:0] Wgt_8_21,
input [18:0] Wgt_8_22,
input [18:0] Wgt_8_23,
input [18:0] Wgt_8_24,
input [18:0] Wgt_8_25,
input [18:0] Wgt_8_26,
input [18:0] Wgt_8_27,
input [18:0] Wgt_8_28,
input [18:0] Wgt_8_29,
input [18:0] Wgt_8_30,
input [18:0] Wgt_8_31,
input [18:0] Wgt_8_32,
input [18:0] Wgt_8_33,
input [18:0] Wgt_8_34,
input [18:0] Wgt_8_35,
input [18:0] Wgt_8_36,
input [18:0] Wgt_8_37,
input [18:0] Wgt_8_38,
input [18:0] Wgt_8_39,
input [18:0] Wgt_8_40,
input [18:0] Wgt_8_41,
input [18:0] Wgt_8_42,
input [18:0] Wgt_8_43,
input [18:0] Wgt_8_44,
input [18:0] Wgt_8_45,
input [18:0] Wgt_8_46,
input [18:0] Wgt_8_47,
input [18:0] Wgt_8_48,
input [18:0] Wgt_8_49,
input [18:0] Wgt_8_50,
input [18:0] Wgt_8_51,
input [18:0] Wgt_8_52,
input [18:0] Wgt_8_53,
input [18:0] Wgt_8_54,
input [18:0] Wgt_8_55,
input [18:0] Wgt_8_56,
input [18:0] Wgt_8_57,
input [18:0] Wgt_8_58,
input [18:0] Wgt_8_59,
input [18:0] Wgt_8_60,
input [18:0] Wgt_8_61,
input [18:0] Wgt_8_62,
input [18:0] Wgt_8_63,
input [18:0] Wgt_8_64,
input [18:0] Wgt_8_65,
input [18:0] Wgt_8_66,
input [18:0] Wgt_8_67,
input [18:0] Wgt_8_68,
input [18:0] Wgt_8_69,
input [18:0] Wgt_8_70,
input [18:0] Wgt_8_71,
input [18:0] Wgt_8_72,
input [18:0] Wgt_8_73,
input [18:0] Wgt_8_74,
input [18:0] Wgt_8_75,
input [18:0] Wgt_8_76,
input [18:0] Wgt_8_77,
input [18:0] Wgt_8_78,
input [18:0] Wgt_8_79,
input [18:0] Wgt_8_80,
input [18:0] Wgt_8_81,
input [18:0] Wgt_8_82,
input [18:0] Wgt_8_83,
input [18:0] Wgt_8_84,
input [18:0] Wgt_8_85,
input [18:0] Wgt_8_86,
input [18:0] Wgt_8_87,
input [18:0] Wgt_8_88,
input [18:0] Wgt_8_89,
input [18:0] Wgt_8_90,
input [18:0] Wgt_8_91,
input [18:0] Wgt_8_92,
input [18:0] Wgt_8_93,
input [18:0] Wgt_8_94,
input [18:0] Wgt_8_95,
input [18:0] Wgt_8_96,
input [18:0] Wgt_8_97,
input [18:0] Wgt_8_98,
input [18:0] Wgt_8_99,
input [18:0] Wgt_8_100,
input [18:0] Wgt_8_101,
input [18:0] Wgt_8_102,
input [18:0] Wgt_8_103,
input [18:0] Wgt_8_104,
input [18:0] Wgt_8_105,
input [18:0] Wgt_8_106,
input [18:0] Wgt_8_107,
input [18:0] Wgt_8_108,
input [18:0] Wgt_8_109,
input [18:0] Wgt_8_110,
input [18:0] Wgt_8_111,
input [18:0] Wgt_8_112,
input [18:0] Wgt_8_113,
input [18:0] Wgt_8_114,
input [18:0] Wgt_8_115,
input [18:0] Wgt_8_116,
input [18:0] Wgt_8_117,
input [18:0] Wgt_8_118,
input [18:0] Wgt_8_119,
input [18:0] Wgt_8_120,
input [18:0] Wgt_8_121,
input [18:0] Wgt_8_122,
input [18:0] Wgt_8_123,
input [18:0] Wgt_8_124,
input [18:0] Wgt_8_125,
input [18:0] Wgt_8_126,
input [18:0] Wgt_8_127,
input [18:0] Wgt_8_128,
input [18:0] Wgt_8_129,
input [18:0] Wgt_8_130,
input [18:0] Wgt_8_131,
input [18:0] Wgt_8_132,
input [18:0] Wgt_8_133,
input [18:0] Wgt_8_134,
input [18:0] Wgt_8_135,
input [18:0] Wgt_8_136,
input [18:0] Wgt_8_137,
input [18:0] Wgt_8_138,
input [18:0] Wgt_8_139,
input [18:0] Wgt_8_140,
input [18:0] Wgt_8_141,
input [18:0] Wgt_8_142,
input [18:0] Wgt_8_143,
input [18:0] Wgt_8_144,
input [18:0] Wgt_8_145,
input [18:0] Wgt_8_146,
input [18:0] Wgt_8_147,
input [18:0] Wgt_8_148,
input [18:0] Wgt_8_149,
input [18:0] Wgt_8_150,
input [18:0] Wgt_8_151,
input [18:0] Wgt_8_152,
input [18:0] Wgt_8_153,
input [18:0] Wgt_8_154,
input [18:0] Wgt_8_155,
input [18:0] Wgt_8_156,
input [18:0] Wgt_8_157,
input [18:0] Wgt_8_158,
input [18:0] Wgt_8_159,
input [18:0] Wgt_8_160,
input [18:0] Wgt_8_161,
input [18:0] Wgt_8_162,
input [18:0] Wgt_8_163,
input [18:0] Wgt_8_164,
input [18:0] Wgt_8_165,
input [18:0] Wgt_8_166,
input [18:0] Wgt_8_167,
input [18:0] Wgt_8_168,
input [18:0] Wgt_8_169,
input [18:0] Wgt_8_170,
input [18:0] Wgt_8_171,
input [18:0] Wgt_8_172,
input [18:0] Wgt_8_173,
input [18:0] Wgt_8_174,
input [18:0] Wgt_8_175,
input [18:0] Wgt_8_176,
input [18:0] Wgt_8_177,
input [18:0] Wgt_8_178,
input [18:0] Wgt_8_179,
input [18:0] Wgt_8_180,
input [18:0] Wgt_8_181,
input [18:0] Wgt_8_182,
input [18:0] Wgt_8_183,
input [18:0] Wgt_8_184,
input [18:0] Wgt_8_185,
input [18:0] Wgt_8_186,
input [18:0] Wgt_8_187,
input [18:0] Wgt_8_188,
input [18:0] Wgt_8_189,
input [18:0] Wgt_8_190,
input [18:0] Wgt_8_191,
input [18:0] Wgt_8_192,
input [18:0] Wgt_8_193,
input [18:0] Wgt_8_194,
input [18:0] Wgt_8_195,
input [18:0] Wgt_8_196,
input [18:0] Wgt_8_197,
input [18:0] Wgt_8_198,
input [18:0] Wgt_8_199,
input [18:0] Wgt_8_200,
input [18:0] Wgt_8_201,
input [18:0] Wgt_8_202,
input [18:0] Wgt_8_203,
input [18:0] Wgt_8_204,
input [18:0] Wgt_8_205,
input [18:0] Wgt_8_206,
input [18:0] Wgt_8_207,
input [18:0] Wgt_8_208,
input [18:0] Wgt_8_209,
input [18:0] Wgt_8_210,
input [18:0] Wgt_8_211,
input [18:0] Wgt_8_212,
input [18:0] Wgt_8_213,
input [18:0] Wgt_8_214,
input [18:0] Wgt_8_215,
input [18:0] Wgt_8_216,
input [18:0] Wgt_8_217,
input [18:0] Wgt_8_218,
input [18:0] Wgt_8_219,
input [18:0] Wgt_8_220,
input [18:0] Wgt_8_221,
input [18:0] Wgt_8_222,
input [18:0] Wgt_8_223,
input [18:0] Wgt_8_224,
input [18:0] Wgt_8_225,
input [18:0] Wgt_8_226,
input [18:0] Wgt_8_227,
input [18:0] Wgt_8_228,
input [18:0] Wgt_8_229,
input [18:0] Wgt_8_230,
input [18:0] Wgt_8_231,
input [18:0] Wgt_8_232,
input [18:0] Wgt_8_233,
input [18:0] Wgt_8_234,
input [18:0] Wgt_8_235,
input [18:0] Wgt_8_236,
input [18:0] Wgt_8_237,
input [18:0] Wgt_8_238,
input [18:0] Wgt_8_239,
input [18:0] Wgt_8_240,
input [18:0] Wgt_8_241,
input [18:0] Wgt_8_242,
input [18:0] Wgt_8_243,
input [18:0] Wgt_8_244,
input [18:0] Wgt_8_245,
input [18:0] Wgt_8_246,
input [18:0] Wgt_8_247,
input [18:0] Wgt_8_248,
input [18:0] Wgt_8_249,
input [18:0] Wgt_8_250,
input [18:0] Wgt_8_251,
input [18:0] Wgt_8_252,
input [18:0] Wgt_8_253,
input [18:0] Wgt_8_254,
input [18:0] Wgt_8_255,
input [18:0] Wgt_8_256,
input [18:0] Wgt_8_257,
input [18:0] Wgt_8_258,
input [18:0] Wgt_8_259,
input [18:0] Wgt_8_260,
input [18:0] Wgt_8_261,
input [18:0] Wgt_8_262,
input [18:0] Wgt_8_263,
input [18:0] Wgt_8_264,
input [18:0] Wgt_8_265,
input [18:0] Wgt_8_266,
input [18:0] Wgt_8_267,
input [18:0] Wgt_8_268,
input [18:0] Wgt_8_269,
input [18:0] Wgt_8_270,
input [18:0] Wgt_8_271,
input [18:0] Wgt_8_272,
input [18:0] Wgt_8_273,
input [18:0] Wgt_8_274,
input [18:0] Wgt_8_275,
input [18:0] Wgt_8_276,
input [18:0] Wgt_8_277,
input [18:0] Wgt_8_278,
input [18:0] Wgt_8_279,
input [18:0] Wgt_8_280,
input [18:0] Wgt_8_281,
input [18:0] Wgt_8_282,
input [18:0] Wgt_8_283,
input [18:0] Wgt_8_284,
input [18:0] Wgt_8_285,
input [18:0] Wgt_8_286,
input [18:0] Wgt_8_287,
input [18:0] Wgt_8_288,
input [18:0] Wgt_8_289,
input [18:0] Wgt_8_290,
input [18:0] Wgt_8_291,
input [18:0] Wgt_8_292,
input [18:0] Wgt_8_293,
input [18:0] Wgt_8_294,
input [18:0] Wgt_8_295,
input [18:0] Wgt_8_296,
input [18:0] Wgt_8_297,
input [18:0] Wgt_8_298,
input [18:0] Wgt_8_299,
input [18:0] Wgt_8_300,
input [18:0] Wgt_8_301,
input [18:0] Wgt_8_302,
input [18:0] Wgt_8_303,
input [18:0] Wgt_8_304,
input [18:0] Wgt_8_305,
input [18:0] Wgt_8_306,
input [18:0] Wgt_8_307,
input [18:0] Wgt_8_308,
input [18:0] Wgt_8_309,
input [18:0] Wgt_8_310,
input [18:0] Wgt_8_311,
input [18:0] Wgt_8_312,
input [18:0] Wgt_8_313,
input [18:0] Wgt_8_314,
input [18:0] Wgt_8_315,
input [18:0] Wgt_8_316,
input [18:0] Wgt_8_317,
input [18:0] Wgt_8_318,
input [18:0] Wgt_8_319,
input [18:0] Wgt_8_320,
input [18:0] Wgt_8_321,
input [18:0] Wgt_8_322,
input [18:0] Wgt_8_323,
input [18:0] Wgt_8_324,
input [18:0] Wgt_8_325,
input [18:0] Wgt_8_326,
input [18:0] Wgt_8_327,
input [18:0] Wgt_8_328,
input [18:0] Wgt_8_329,
input [18:0] Wgt_8_330,
input [18:0] Wgt_8_331,
input [18:0] Wgt_8_332,
input [18:0] Wgt_8_333,
input [18:0] Wgt_8_334,
input [18:0] Wgt_8_335,
input [18:0] Wgt_8_336,
input [18:0] Wgt_8_337,
input [18:0] Wgt_8_338,
input [18:0] Wgt_8_339,
input [18:0] Wgt_8_340,
input [18:0] Wgt_8_341,
input [18:0] Wgt_8_342,
input [18:0] Wgt_8_343,
input [18:0] Wgt_8_344,
input [18:0] Wgt_8_345,
input [18:0] Wgt_8_346,
input [18:0] Wgt_8_347,
input [18:0] Wgt_8_348,
input [18:0] Wgt_8_349,
input [18:0] Wgt_8_350,
input [18:0] Wgt_8_351,
input [18:0] Wgt_8_352,
input [18:0] Wgt_8_353,
input [18:0] Wgt_8_354,
input [18:0] Wgt_8_355,
input [18:0] Wgt_8_356,
input [18:0] Wgt_8_357,
input [18:0] Wgt_8_358,
input [18:0] Wgt_8_359,
input [18:0] Wgt_8_360,
input [18:0] Wgt_8_361,
input [18:0] Wgt_8_362,
input [18:0] Wgt_8_363,
input [18:0] Wgt_8_364,
input [18:0] Wgt_8_365,
input [18:0] Wgt_8_366,
input [18:0] Wgt_8_367,
input [18:0] Wgt_8_368,
input [18:0] Wgt_8_369,
input [18:0] Wgt_8_370,
input [18:0] Wgt_8_371,
input [18:0] Wgt_8_372,
input [18:0] Wgt_8_373,
input [18:0] Wgt_8_374,
input [18:0] Wgt_8_375,
input [18:0] Wgt_8_376,
input [18:0] Wgt_8_377,
input [18:0] Wgt_8_378,
input [18:0] Wgt_8_379,
input [18:0] Wgt_8_380,
input [18:0] Wgt_8_381,
input [18:0] Wgt_8_382,
input [18:0] Wgt_8_383,
input [18:0] Wgt_8_384,
input [18:0] Wgt_8_385,
input [18:0] Wgt_8_386,
input [18:0] Wgt_8_387,
input [18:0] Wgt_8_388,
input [18:0] Wgt_8_389,
input [18:0] Wgt_8_390,
input [18:0] Wgt_8_391,
input [18:0] Wgt_8_392,
input [18:0] Wgt_8_393,
input [18:0] Wgt_8_394,
input [18:0] Wgt_8_395,
input [18:0] Wgt_8_396,
input [18:0] Wgt_8_397,
input [18:0] Wgt_8_398,
input [18:0] Wgt_8_399,
input [18:0] Wgt_8_400,
input [18:0] Wgt_8_401,
input [18:0] Wgt_8_402,
input [18:0] Wgt_8_403,
input [18:0] Wgt_8_404,
input [18:0] Wgt_8_405,
input [18:0] Wgt_8_406,
input [18:0] Wgt_8_407,
input [18:0] Wgt_8_408,
input [18:0] Wgt_8_409,
input [18:0] Wgt_8_410,
input [18:0] Wgt_8_411,
input [18:0] Wgt_8_412,
input [18:0] Wgt_8_413,
input [18:0] Wgt_8_414,
input [18:0] Wgt_8_415,
input [18:0] Wgt_8_416,
input [18:0] Wgt_8_417,
input [18:0] Wgt_8_418,
input [18:0] Wgt_8_419,
input [18:0] Wgt_8_420,
input [18:0] Wgt_8_421,
input [18:0] Wgt_8_422,
input [18:0] Wgt_8_423,
input [18:0] Wgt_8_424,
input [18:0] Wgt_8_425,
input [18:0] Wgt_8_426,
input [18:0] Wgt_8_427,
input [18:0] Wgt_8_428,
input [18:0] Wgt_8_429,
input [18:0] Wgt_8_430,
input [18:0] Wgt_8_431,
input [18:0] Wgt_8_432,
input [18:0] Wgt_8_433,
input [18:0] Wgt_8_434,
input [18:0] Wgt_8_435,
input [18:0] Wgt_8_436,
input [18:0] Wgt_8_437,
input [18:0] Wgt_8_438,
input [18:0] Wgt_8_439,
input [18:0] Wgt_8_440,
input [18:0] Wgt_8_441,
input [18:0] Wgt_8_442,
input [18:0] Wgt_8_443,
input [18:0] Wgt_8_444,
input [18:0] Wgt_8_445,
input [18:0] Wgt_8_446,
input [18:0] Wgt_8_447,
input [18:0] Wgt_8_448,
input [18:0] Wgt_8_449,
input [18:0] Wgt_8_450,
input [18:0] Wgt_8_451,
input [18:0] Wgt_8_452,
input [18:0] Wgt_8_453,
input [18:0] Wgt_8_454,
input [18:0] Wgt_8_455,
input [18:0] Wgt_8_456,
input [18:0] Wgt_8_457,
input [18:0] Wgt_8_458,
input [18:0] Wgt_8_459,
input [18:0] Wgt_8_460,
input [18:0] Wgt_8_461,
input [18:0] Wgt_8_462,
input [18:0] Wgt_8_463,
input [18:0] Wgt_8_464,
input [18:0] Wgt_8_465,
input [18:0] Wgt_8_466,
input [18:0] Wgt_8_467,
input [18:0] Wgt_8_468,
input [18:0] Wgt_8_469,
input [18:0] Wgt_8_470,
input [18:0] Wgt_8_471,
input [18:0] Wgt_8_472,
input [18:0] Wgt_8_473,
input [18:0] Wgt_8_474,
input [18:0] Wgt_8_475,
input [18:0] Wgt_8_476,
input [18:0] Wgt_8_477,
input [18:0] Wgt_8_478,
input [18:0] Wgt_8_479,
input [18:0] Wgt_8_480,
input [18:0] Wgt_8_481,
input [18:0] Wgt_8_482,
input [18:0] Wgt_8_483,
input [18:0] Wgt_8_484,
input [18:0] Wgt_8_485,
input [18:0] Wgt_8_486,
input [18:0] Wgt_8_487,
input [18:0] Wgt_8_488,
input [18:0] Wgt_8_489,
input [18:0] Wgt_8_490,
input [18:0] Wgt_8_491,
input [18:0] Wgt_8_492,
input [18:0] Wgt_8_493,
input [18:0] Wgt_8_494,
input [18:0] Wgt_8_495,
input [18:0] Wgt_8_496,
input [18:0] Wgt_8_497,
input [18:0] Wgt_8_498,
input [18:0] Wgt_8_499,
input [18:0] Wgt_8_500,
input [18:0] Wgt_8_501,
input [18:0] Wgt_8_502,
input [18:0] Wgt_8_503,
input [18:0] Wgt_8_504,
input [18:0] Wgt_8_505,
input [18:0] Wgt_8_506,
input [18:0] Wgt_8_507,
input [18:0] Wgt_8_508,
input [18:0] Wgt_8_509,
input [18:0] Wgt_8_510,
input [18:0] Wgt_8_511,
input [18:0] Wgt_8_512,
input [18:0] Wgt_8_513,
input [18:0] Wgt_8_514,
input [18:0] Wgt_8_515,
input [18:0] Wgt_8_516,
input [18:0] Wgt_8_517,
input [18:0] Wgt_8_518,
input [18:0] Wgt_8_519,
input [18:0] Wgt_8_520,
input [18:0] Wgt_8_521,
input [18:0] Wgt_8_522,
input [18:0] Wgt_8_523,
input [18:0] Wgt_8_524,
input [18:0] Wgt_8_525,
input [18:0] Wgt_8_526,
input [18:0] Wgt_8_527,
input [18:0] Wgt_8_528,
input [18:0] Wgt_8_529,
input [18:0] Wgt_8_530,
input [18:0] Wgt_8_531,
input [18:0] Wgt_8_532,
input [18:0] Wgt_8_533,
input [18:0] Wgt_8_534,
input [18:0] Wgt_8_535,
input [18:0] Wgt_8_536,
input [18:0] Wgt_8_537,
input [18:0] Wgt_8_538,
input [18:0] Wgt_8_539,
input [18:0] Wgt_8_540,
input [18:0] Wgt_8_541,
input [18:0] Wgt_8_542,
input [18:0] Wgt_8_543,
input [18:0] Wgt_8_544,
input [18:0] Wgt_8_545,
input [18:0] Wgt_8_546,
input [18:0] Wgt_8_547,
input [18:0] Wgt_8_548,
input [18:0] Wgt_8_549,
input [18:0] Wgt_8_550,
input [18:0] Wgt_8_551,
input [18:0] Wgt_8_552,
input [18:0] Wgt_8_553,
input [18:0] Wgt_8_554,
input [18:0] Wgt_8_555,
input [18:0] Wgt_8_556,
input [18:0] Wgt_8_557,
input [18:0] Wgt_8_558,
input [18:0] Wgt_8_559,
input [18:0] Wgt_8_560,
input [18:0] Wgt_8_561,
input [18:0] Wgt_8_562,
input [18:0] Wgt_8_563,
input [18:0] Wgt_8_564,
input [18:0] Wgt_8_565,
input [18:0] Wgt_8_566,
input [18:0] Wgt_8_567,
input [18:0] Wgt_8_568,
input [18:0] Wgt_8_569,
input [18:0] Wgt_8_570,
input [18:0] Wgt_8_571,
input [18:0] Wgt_8_572,
input [18:0] Wgt_8_573,
input [18:0] Wgt_8_574,
input [18:0] Wgt_8_575,
input [18:0] Wgt_8_576,
input [18:0] Wgt_8_577,
input [18:0] Wgt_8_578,
input [18:0] Wgt_8_579,
input [18:0] Wgt_8_580,
input [18:0] Wgt_8_581,
input [18:0] Wgt_8_582,
input [18:0] Wgt_8_583,
input [18:0] Wgt_8_584,
input [18:0] Wgt_8_585,
input [18:0] Wgt_8_586,
input [18:0] Wgt_8_587,
input [18:0] Wgt_8_588,
input [18:0] Wgt_8_589,
input [18:0] Wgt_8_590,
input [18:0] Wgt_8_591,
input [18:0] Wgt_8_592,
input [18:0] Wgt_8_593,
input [18:0] Wgt_8_594,
input [18:0] Wgt_8_595,
input [18:0] Wgt_8_596,
input [18:0] Wgt_8_597,
input [18:0] Wgt_8_598,
input [18:0] Wgt_8_599,
input [18:0] Wgt_8_600,
input [18:0] Wgt_8_601,
input [18:0] Wgt_8_602,
input [18:0] Wgt_8_603,
input [18:0] Wgt_8_604,
input [18:0] Wgt_8_605,
input [18:0] Wgt_8_606,
input [18:0] Wgt_8_607,
input [18:0] Wgt_8_608,
input [18:0] Wgt_8_609,
input [18:0] Wgt_8_610,
input [18:0] Wgt_8_611,
input [18:0] Wgt_8_612,
input [18:0] Wgt_8_613,
input [18:0] Wgt_8_614,
input [18:0] Wgt_8_615,
input [18:0] Wgt_8_616,
input [18:0] Wgt_8_617,
input [18:0] Wgt_8_618,
input [18:0] Wgt_8_619,
input [18:0] Wgt_8_620,
input [18:0] Wgt_8_621,
input [18:0] Wgt_8_622,
input [18:0] Wgt_8_623,
input [18:0] Wgt_8_624,
input [18:0] Wgt_8_625,
input [18:0] Wgt_8_626,
input [18:0] Wgt_8_627,
input [18:0] Wgt_8_628,
input [18:0] Wgt_8_629,
input [18:0] Wgt_8_630,
input [18:0] Wgt_8_631,
input [18:0] Wgt_8_632,
input [18:0] Wgt_8_633,
input [18:0] Wgt_8_634,
input [18:0] Wgt_8_635,
input [18:0] Wgt_8_636,
input [18:0] Wgt_8_637,
input [18:0] Wgt_8_638,
input [18:0] Wgt_8_639,
input [18:0] Wgt_8_640,
input [18:0] Wgt_8_641,
input [18:0] Wgt_8_642,
input [18:0] Wgt_8_643,
input [18:0] Wgt_8_644,
input [18:0] Wgt_8_645,
input [18:0] Wgt_8_646,
input [18:0] Wgt_8_647,
input [18:0] Wgt_8_648,
input [18:0] Wgt_8_649,
input [18:0] Wgt_8_650,
input [18:0] Wgt_8_651,
input [18:0] Wgt_8_652,
input [18:0] Wgt_8_653,
input [18:0] Wgt_8_654,
input [18:0] Wgt_8_655,
input [18:0] Wgt_8_656,
input [18:0] Wgt_8_657,
input [18:0] Wgt_8_658,
input [18:0] Wgt_8_659,
input [18:0] Wgt_8_660,
input [18:0] Wgt_8_661,
input [18:0] Wgt_8_662,
input [18:0] Wgt_8_663,
input [18:0] Wgt_8_664,
input [18:0] Wgt_8_665,
input [18:0] Wgt_8_666,
input [18:0] Wgt_8_667,
input [18:0] Wgt_8_668,
input [18:0] Wgt_8_669,
input [18:0] Wgt_8_670,
input [18:0] Wgt_8_671,
input [18:0] Wgt_8_672,
input [18:0] Wgt_8_673,
input [18:0] Wgt_8_674,
input [18:0] Wgt_8_675,
input [18:0] Wgt_8_676,
input [18:0] Wgt_8_677,
input [18:0] Wgt_8_678,
input [18:0] Wgt_8_679,
input [18:0] Wgt_8_680,
input [18:0] Wgt_8_681,
input [18:0] Wgt_8_682,
input [18:0] Wgt_8_683,
input [18:0] Wgt_8_684,
input [18:0] Wgt_8_685,
input [18:0] Wgt_8_686,
input [18:0] Wgt_8_687,
input [18:0] Wgt_8_688,
input [18:0] Wgt_8_689,
input [18:0] Wgt_8_690,
input [18:0] Wgt_8_691,
input [18:0] Wgt_8_692,
input [18:0] Wgt_8_693,
input [18:0] Wgt_8_694,
input [18:0] Wgt_8_695,
input [18:0] Wgt_8_696,
input [18:0] Wgt_8_697,
input [18:0] Wgt_8_698,
input [18:0] Wgt_8_699,
input [18:0] Wgt_8_700,
input [18:0] Wgt_8_701,
input [18:0] Wgt_8_702,
input [18:0] Wgt_8_703,
input [18:0] Wgt_8_704,
input [18:0] Wgt_8_705,
input [18:0] Wgt_8_706,
input [18:0] Wgt_8_707,
input [18:0] Wgt_8_708,
input [18:0] Wgt_8_709,
input [18:0] Wgt_8_710,
input [18:0] Wgt_8_711,
input [18:0] Wgt_8_712,
input [18:0] Wgt_8_713,
input [18:0] Wgt_8_714,
input [18:0] Wgt_8_715,
input [18:0] Wgt_8_716,
input [18:0] Wgt_8_717,
input [18:0] Wgt_8_718,
input [18:0] Wgt_8_719,
input [18:0] Wgt_8_720,
input [18:0] Wgt_8_721,
input [18:0] Wgt_8_722,
input [18:0] Wgt_8_723,
input [18:0] Wgt_8_724,
input [18:0] Wgt_8_725,
input [18:0] Wgt_8_726,
input [18:0] Wgt_8_727,
input [18:0] Wgt_8_728,
input [18:0] Wgt_8_729,
input [18:0] Wgt_8_730,
input [18:0] Wgt_8_731,
input [18:0] Wgt_8_732,
input [18:0] Wgt_8_733,
input [18:0] Wgt_8_734,
input [18:0] Wgt_8_735,
input [18:0] Wgt_8_736,
input [18:0] Wgt_8_737,
input [18:0] Wgt_8_738,
input [18:0] Wgt_8_739,
input [18:0] Wgt_8_740,
input [18:0] Wgt_8_741,
input [18:0] Wgt_8_742,
input [18:0] Wgt_8_743,
input [18:0] Wgt_8_744,
input [18:0] Wgt_8_745,
input [18:0] Wgt_8_746,
input [18:0] Wgt_8_747,
input [18:0] Wgt_8_748,
input [18:0] Wgt_8_749,
input [18:0] Wgt_8_750,
input [18:0] Wgt_8_751,
input [18:0] Wgt_8_752,
input [18:0] Wgt_8_753,
input [18:0] Wgt_8_754,
input [18:0] Wgt_8_755,
input [18:0] Wgt_8_756,
input [18:0] Wgt_8_757,
input [18:0] Wgt_8_758,
input [18:0] Wgt_8_759,
input [18:0] Wgt_8_760,
input [18:0] Wgt_8_761,
input [18:0] Wgt_8_762,
input [18:0] Wgt_8_763,
input [18:0] Wgt_8_764,
input [18:0] Wgt_8_765,
input [18:0] Wgt_8_766,
input [18:0] Wgt_8_767,
input [18:0] Wgt_8_768,
input [18:0] Wgt_8_769,
input [18:0] Wgt_8_770,
input [18:0] Wgt_8_771,
input [18:0] Wgt_8_772,
input [18:0] Wgt_8_773,
input [18:0] Wgt_8_774,
input [18:0] Wgt_8_775,
input [18:0] Wgt_8_776,
input [18:0] Wgt_8_777,
input [18:0] Wgt_8_778,
input [18:0] Wgt_8_779,
input [18:0] Wgt_8_780,
input [18:0] Wgt_8_781,
input [18:0] Wgt_8_782,
input [18:0] Wgt_8_783,
input [18:0] Wgt_8_784,
input [18:0] Wgt_9_0,
input [18:0] Wgt_9_1,
input [18:0] Wgt_9_2,
input [18:0] Wgt_9_3,
input [18:0] Wgt_9_4,
input [18:0] Wgt_9_5,
input [18:0] Wgt_9_6,
input [18:0] Wgt_9_7,
input [18:0] Wgt_9_8,
input [18:0] Wgt_9_9,
input [18:0] Wgt_9_10,
input [18:0] Wgt_9_11,
input [18:0] Wgt_9_12,
input [18:0] Wgt_9_13,
input [18:0] Wgt_9_14,
input [18:0] Wgt_9_15,
input [18:0] Wgt_9_16,
input [18:0] Wgt_9_17,
input [18:0] Wgt_9_18,
input [18:0] Wgt_9_19,
input [18:0] Wgt_9_20,
input [18:0] Wgt_9_21,
input [18:0] Wgt_9_22,
input [18:0] Wgt_9_23,
input [18:0] Wgt_9_24,
input [18:0] Wgt_9_25,
input [18:0] Wgt_9_26,
input [18:0] Wgt_9_27,
input [18:0] Wgt_9_28,
input [18:0] Wgt_9_29,
input [18:0] Wgt_9_30,
input [18:0] Wgt_9_31,
input [18:0] Wgt_9_32,
input [18:0] Wgt_9_33,
input [18:0] Wgt_9_34,
input [18:0] Wgt_9_35,
input [18:0] Wgt_9_36,
input [18:0] Wgt_9_37,
input [18:0] Wgt_9_38,
input [18:0] Wgt_9_39,
input [18:0] Wgt_9_40,
input [18:0] Wgt_9_41,
input [18:0] Wgt_9_42,
input [18:0] Wgt_9_43,
input [18:0] Wgt_9_44,
input [18:0] Wgt_9_45,
input [18:0] Wgt_9_46,
input [18:0] Wgt_9_47,
input [18:0] Wgt_9_48,
input [18:0] Wgt_9_49,
input [18:0] Wgt_9_50,
input [18:0] Wgt_9_51,
input [18:0] Wgt_9_52,
input [18:0] Wgt_9_53,
input [18:0] Wgt_9_54,
input [18:0] Wgt_9_55,
input [18:0] Wgt_9_56,
input [18:0] Wgt_9_57,
input [18:0] Wgt_9_58,
input [18:0] Wgt_9_59,
input [18:0] Wgt_9_60,
input [18:0] Wgt_9_61,
input [18:0] Wgt_9_62,
input [18:0] Wgt_9_63,
input [18:0] Wgt_9_64,
input [18:0] Wgt_9_65,
input [18:0] Wgt_9_66,
input [18:0] Wgt_9_67,
input [18:0] Wgt_9_68,
input [18:0] Wgt_9_69,
input [18:0] Wgt_9_70,
input [18:0] Wgt_9_71,
input [18:0] Wgt_9_72,
input [18:0] Wgt_9_73,
input [18:0] Wgt_9_74,
input [18:0] Wgt_9_75,
input [18:0] Wgt_9_76,
input [18:0] Wgt_9_77,
input [18:0] Wgt_9_78,
input [18:0] Wgt_9_79,
input [18:0] Wgt_9_80,
input [18:0] Wgt_9_81,
input [18:0] Wgt_9_82,
input [18:0] Wgt_9_83,
input [18:0] Wgt_9_84,
input [18:0] Wgt_9_85,
input [18:0] Wgt_9_86,
input [18:0] Wgt_9_87,
input [18:0] Wgt_9_88,
input [18:0] Wgt_9_89,
input [18:0] Wgt_9_90,
input [18:0] Wgt_9_91,
input [18:0] Wgt_9_92,
input [18:0] Wgt_9_93,
input [18:0] Wgt_9_94,
input [18:0] Wgt_9_95,
input [18:0] Wgt_9_96,
input [18:0] Wgt_9_97,
input [18:0] Wgt_9_98,
input [18:0] Wgt_9_99,
input [18:0] Wgt_9_100,
input [18:0] Wgt_9_101,
input [18:0] Wgt_9_102,
input [18:0] Wgt_9_103,
input [18:0] Wgt_9_104,
input [18:0] Wgt_9_105,
input [18:0] Wgt_9_106,
input [18:0] Wgt_9_107,
input [18:0] Wgt_9_108,
input [18:0] Wgt_9_109,
input [18:0] Wgt_9_110,
input [18:0] Wgt_9_111,
input [18:0] Wgt_9_112,
input [18:0] Wgt_9_113,
input [18:0] Wgt_9_114,
input [18:0] Wgt_9_115,
input [18:0] Wgt_9_116,
input [18:0] Wgt_9_117,
input [18:0] Wgt_9_118,
input [18:0] Wgt_9_119,
input [18:0] Wgt_9_120,
input [18:0] Wgt_9_121,
input [18:0] Wgt_9_122,
input [18:0] Wgt_9_123,
input [18:0] Wgt_9_124,
input [18:0] Wgt_9_125,
input [18:0] Wgt_9_126,
input [18:0] Wgt_9_127,
input [18:0] Wgt_9_128,
input [18:0] Wgt_9_129,
input [18:0] Wgt_9_130,
input [18:0] Wgt_9_131,
input [18:0] Wgt_9_132,
input [18:0] Wgt_9_133,
input [18:0] Wgt_9_134,
input [18:0] Wgt_9_135,
input [18:0] Wgt_9_136,
input [18:0] Wgt_9_137,
input [18:0] Wgt_9_138,
input [18:0] Wgt_9_139,
input [18:0] Wgt_9_140,
input [18:0] Wgt_9_141,
input [18:0] Wgt_9_142,
input [18:0] Wgt_9_143,
input [18:0] Wgt_9_144,
input [18:0] Wgt_9_145,
input [18:0] Wgt_9_146,
input [18:0] Wgt_9_147,
input [18:0] Wgt_9_148,
input [18:0] Wgt_9_149,
input [18:0] Wgt_9_150,
input [18:0] Wgt_9_151,
input [18:0] Wgt_9_152,
input [18:0] Wgt_9_153,
input [18:0] Wgt_9_154,
input [18:0] Wgt_9_155,
input [18:0] Wgt_9_156,
input [18:0] Wgt_9_157,
input [18:0] Wgt_9_158,
input [18:0] Wgt_9_159,
input [18:0] Wgt_9_160,
input [18:0] Wgt_9_161,
input [18:0] Wgt_9_162,
input [18:0] Wgt_9_163,
input [18:0] Wgt_9_164,
input [18:0] Wgt_9_165,
input [18:0] Wgt_9_166,
input [18:0] Wgt_9_167,
input [18:0] Wgt_9_168,
input [18:0] Wgt_9_169,
input [18:0] Wgt_9_170,
input [18:0] Wgt_9_171,
input [18:0] Wgt_9_172,
input [18:0] Wgt_9_173,
input [18:0] Wgt_9_174,
input [18:0] Wgt_9_175,
input [18:0] Wgt_9_176,
input [18:0] Wgt_9_177,
input [18:0] Wgt_9_178,
input [18:0] Wgt_9_179,
input [18:0] Wgt_9_180,
input [18:0] Wgt_9_181,
input [18:0] Wgt_9_182,
input [18:0] Wgt_9_183,
input [18:0] Wgt_9_184,
input [18:0] Wgt_9_185,
input [18:0] Wgt_9_186,
input [18:0] Wgt_9_187,
input [18:0] Wgt_9_188,
input [18:0] Wgt_9_189,
input [18:0] Wgt_9_190,
input [18:0] Wgt_9_191,
input [18:0] Wgt_9_192,
input [18:0] Wgt_9_193,
input [18:0] Wgt_9_194,
input [18:0] Wgt_9_195,
input [18:0] Wgt_9_196,
input [18:0] Wgt_9_197,
input [18:0] Wgt_9_198,
input [18:0] Wgt_9_199,
input [18:0] Wgt_9_200,
input [18:0] Wgt_9_201,
input [18:0] Wgt_9_202,
input [18:0] Wgt_9_203,
input [18:0] Wgt_9_204,
input [18:0] Wgt_9_205,
input [18:0] Wgt_9_206,
input [18:0] Wgt_9_207,
input [18:0] Wgt_9_208,
input [18:0] Wgt_9_209,
input [18:0] Wgt_9_210,
input [18:0] Wgt_9_211,
input [18:0] Wgt_9_212,
input [18:0] Wgt_9_213,
input [18:0] Wgt_9_214,
input [18:0] Wgt_9_215,
input [18:0] Wgt_9_216,
input [18:0] Wgt_9_217,
input [18:0] Wgt_9_218,
input [18:0] Wgt_9_219,
input [18:0] Wgt_9_220,
input [18:0] Wgt_9_221,
input [18:0] Wgt_9_222,
input [18:0] Wgt_9_223,
input [18:0] Wgt_9_224,
input [18:0] Wgt_9_225,
input [18:0] Wgt_9_226,
input [18:0] Wgt_9_227,
input [18:0] Wgt_9_228,
input [18:0] Wgt_9_229,
input [18:0] Wgt_9_230,
input [18:0] Wgt_9_231,
input [18:0] Wgt_9_232,
input [18:0] Wgt_9_233,
input [18:0] Wgt_9_234,
input [18:0] Wgt_9_235,
input [18:0] Wgt_9_236,
input [18:0] Wgt_9_237,
input [18:0] Wgt_9_238,
input [18:0] Wgt_9_239,
input [18:0] Wgt_9_240,
input [18:0] Wgt_9_241,
input [18:0] Wgt_9_242,
input [18:0] Wgt_9_243,
input [18:0] Wgt_9_244,
input [18:0] Wgt_9_245,
input [18:0] Wgt_9_246,
input [18:0] Wgt_9_247,
input [18:0] Wgt_9_248,
input [18:0] Wgt_9_249,
input [18:0] Wgt_9_250,
input [18:0] Wgt_9_251,
input [18:0] Wgt_9_252,
input [18:0] Wgt_9_253,
input [18:0] Wgt_9_254,
input [18:0] Wgt_9_255,
input [18:0] Wgt_9_256,
input [18:0] Wgt_9_257,
input [18:0] Wgt_9_258,
input [18:0] Wgt_9_259,
input [18:0] Wgt_9_260,
input [18:0] Wgt_9_261,
input [18:0] Wgt_9_262,
input [18:0] Wgt_9_263,
input [18:0] Wgt_9_264,
input [18:0] Wgt_9_265,
input [18:0] Wgt_9_266,
input [18:0] Wgt_9_267,
input [18:0] Wgt_9_268,
input [18:0] Wgt_9_269,
input [18:0] Wgt_9_270,
input [18:0] Wgt_9_271,
input [18:0] Wgt_9_272,
input [18:0] Wgt_9_273,
input [18:0] Wgt_9_274,
input [18:0] Wgt_9_275,
input [18:0] Wgt_9_276,
input [18:0] Wgt_9_277,
input [18:0] Wgt_9_278,
input [18:0] Wgt_9_279,
input [18:0] Wgt_9_280,
input [18:0] Wgt_9_281,
input [18:0] Wgt_9_282,
input [18:0] Wgt_9_283,
input [18:0] Wgt_9_284,
input [18:0] Wgt_9_285,
input [18:0] Wgt_9_286,
input [18:0] Wgt_9_287,
input [18:0] Wgt_9_288,
input [18:0] Wgt_9_289,
input [18:0] Wgt_9_290,
input [18:0] Wgt_9_291,
input [18:0] Wgt_9_292,
input [18:0] Wgt_9_293,
input [18:0] Wgt_9_294,
input [18:0] Wgt_9_295,
input [18:0] Wgt_9_296,
input [18:0] Wgt_9_297,
input [18:0] Wgt_9_298,
input [18:0] Wgt_9_299,
input [18:0] Wgt_9_300,
input [18:0] Wgt_9_301,
input [18:0] Wgt_9_302,
input [18:0] Wgt_9_303,
input [18:0] Wgt_9_304,
input [18:0] Wgt_9_305,
input [18:0] Wgt_9_306,
input [18:0] Wgt_9_307,
input [18:0] Wgt_9_308,
input [18:0] Wgt_9_309,
input [18:0] Wgt_9_310,
input [18:0] Wgt_9_311,
input [18:0] Wgt_9_312,
input [18:0] Wgt_9_313,
input [18:0] Wgt_9_314,
input [18:0] Wgt_9_315,
input [18:0] Wgt_9_316,
input [18:0] Wgt_9_317,
input [18:0] Wgt_9_318,
input [18:0] Wgt_9_319,
input [18:0] Wgt_9_320,
input [18:0] Wgt_9_321,
input [18:0] Wgt_9_322,
input [18:0] Wgt_9_323,
input [18:0] Wgt_9_324,
input [18:0] Wgt_9_325,
input [18:0] Wgt_9_326,
input [18:0] Wgt_9_327,
input [18:0] Wgt_9_328,
input [18:0] Wgt_9_329,
input [18:0] Wgt_9_330,
input [18:0] Wgt_9_331,
input [18:0] Wgt_9_332,
input [18:0] Wgt_9_333,
input [18:0] Wgt_9_334,
input [18:0] Wgt_9_335,
input [18:0] Wgt_9_336,
input [18:0] Wgt_9_337,
input [18:0] Wgt_9_338,
input [18:0] Wgt_9_339,
input [18:0] Wgt_9_340,
input [18:0] Wgt_9_341,
input [18:0] Wgt_9_342,
input [18:0] Wgt_9_343,
input [18:0] Wgt_9_344,
input [18:0] Wgt_9_345,
input [18:0] Wgt_9_346,
input [18:0] Wgt_9_347,
input [18:0] Wgt_9_348,
input [18:0] Wgt_9_349,
input [18:0] Wgt_9_350,
input [18:0] Wgt_9_351,
input [18:0] Wgt_9_352,
input [18:0] Wgt_9_353,
input [18:0] Wgt_9_354,
input [18:0] Wgt_9_355,
input [18:0] Wgt_9_356,
input [18:0] Wgt_9_357,
input [18:0] Wgt_9_358,
input [18:0] Wgt_9_359,
input [18:0] Wgt_9_360,
input [18:0] Wgt_9_361,
input [18:0] Wgt_9_362,
input [18:0] Wgt_9_363,
input [18:0] Wgt_9_364,
input [18:0] Wgt_9_365,
input [18:0] Wgt_9_366,
input [18:0] Wgt_9_367,
input [18:0] Wgt_9_368,
input [18:0] Wgt_9_369,
input [18:0] Wgt_9_370,
input [18:0] Wgt_9_371,
input [18:0] Wgt_9_372,
input [18:0] Wgt_9_373,
input [18:0] Wgt_9_374,
input [18:0] Wgt_9_375,
input [18:0] Wgt_9_376,
input [18:0] Wgt_9_377,
input [18:0] Wgt_9_378,
input [18:0] Wgt_9_379,
input [18:0] Wgt_9_380,
input [18:0] Wgt_9_381,
input [18:0] Wgt_9_382,
input [18:0] Wgt_9_383,
input [18:0] Wgt_9_384,
input [18:0] Wgt_9_385,
input [18:0] Wgt_9_386,
input [18:0] Wgt_9_387,
input [18:0] Wgt_9_388,
input [18:0] Wgt_9_389,
input [18:0] Wgt_9_390,
input [18:0] Wgt_9_391,
input [18:0] Wgt_9_392,
input [18:0] Wgt_9_393,
input [18:0] Wgt_9_394,
input [18:0] Wgt_9_395,
input [18:0] Wgt_9_396,
input [18:0] Wgt_9_397,
input [18:0] Wgt_9_398,
input [18:0] Wgt_9_399,
input [18:0] Wgt_9_400,
input [18:0] Wgt_9_401,
input [18:0] Wgt_9_402,
input [18:0] Wgt_9_403,
input [18:0] Wgt_9_404,
input [18:0] Wgt_9_405,
input [18:0] Wgt_9_406,
input [18:0] Wgt_9_407,
input [18:0] Wgt_9_408,
input [18:0] Wgt_9_409,
input [18:0] Wgt_9_410,
input [18:0] Wgt_9_411,
input [18:0] Wgt_9_412,
input [18:0] Wgt_9_413,
input [18:0] Wgt_9_414,
input [18:0] Wgt_9_415,
input [18:0] Wgt_9_416,
input [18:0] Wgt_9_417,
input [18:0] Wgt_9_418,
input [18:0] Wgt_9_419,
input [18:0] Wgt_9_420,
input [18:0] Wgt_9_421,
input [18:0] Wgt_9_422,
input [18:0] Wgt_9_423,
input [18:0] Wgt_9_424,
input [18:0] Wgt_9_425,
input [18:0] Wgt_9_426,
input [18:0] Wgt_9_427,
input [18:0] Wgt_9_428,
input [18:0] Wgt_9_429,
input [18:0] Wgt_9_430,
input [18:0] Wgt_9_431,
input [18:0] Wgt_9_432,
input [18:0] Wgt_9_433,
input [18:0] Wgt_9_434,
input [18:0] Wgt_9_435,
input [18:0] Wgt_9_436,
input [18:0] Wgt_9_437,
input [18:0] Wgt_9_438,
input [18:0] Wgt_9_439,
input [18:0] Wgt_9_440,
input [18:0] Wgt_9_441,
input [18:0] Wgt_9_442,
input [18:0] Wgt_9_443,
input [18:0] Wgt_9_444,
input [18:0] Wgt_9_445,
input [18:0] Wgt_9_446,
input [18:0] Wgt_9_447,
input [18:0] Wgt_9_448,
input [18:0] Wgt_9_449,
input [18:0] Wgt_9_450,
input [18:0] Wgt_9_451,
input [18:0] Wgt_9_452,
input [18:0] Wgt_9_453,
input [18:0] Wgt_9_454,
input [18:0] Wgt_9_455,
input [18:0] Wgt_9_456,
input [18:0] Wgt_9_457,
input [18:0] Wgt_9_458,
input [18:0] Wgt_9_459,
input [18:0] Wgt_9_460,
input [18:0] Wgt_9_461,
input [18:0] Wgt_9_462,
input [18:0] Wgt_9_463,
input [18:0] Wgt_9_464,
input [18:0] Wgt_9_465,
input [18:0] Wgt_9_466,
input [18:0] Wgt_9_467,
input [18:0] Wgt_9_468,
input [18:0] Wgt_9_469,
input [18:0] Wgt_9_470,
input [18:0] Wgt_9_471,
input [18:0] Wgt_9_472,
input [18:0] Wgt_9_473,
input [18:0] Wgt_9_474,
input [18:0] Wgt_9_475,
input [18:0] Wgt_9_476,
input [18:0] Wgt_9_477,
input [18:0] Wgt_9_478,
input [18:0] Wgt_9_479,
input [18:0] Wgt_9_480,
input [18:0] Wgt_9_481,
input [18:0] Wgt_9_482,
input [18:0] Wgt_9_483,
input [18:0] Wgt_9_484,
input [18:0] Wgt_9_485,
input [18:0] Wgt_9_486,
input [18:0] Wgt_9_487,
input [18:0] Wgt_9_488,
input [18:0] Wgt_9_489,
input [18:0] Wgt_9_490,
input [18:0] Wgt_9_491,
input [18:0] Wgt_9_492,
input [18:0] Wgt_9_493,
input [18:0] Wgt_9_494,
input [18:0] Wgt_9_495,
input [18:0] Wgt_9_496,
input [18:0] Wgt_9_497,
input [18:0] Wgt_9_498,
input [18:0] Wgt_9_499,
input [18:0] Wgt_9_500,
input [18:0] Wgt_9_501,
input [18:0] Wgt_9_502,
input [18:0] Wgt_9_503,
input [18:0] Wgt_9_504,
input [18:0] Wgt_9_505,
input [18:0] Wgt_9_506,
input [18:0] Wgt_9_507,
input [18:0] Wgt_9_508,
input [18:0] Wgt_9_509,
input [18:0] Wgt_9_510,
input [18:0] Wgt_9_511,
input [18:0] Wgt_9_512,
input [18:0] Wgt_9_513,
input [18:0] Wgt_9_514,
input [18:0] Wgt_9_515,
input [18:0] Wgt_9_516,
input [18:0] Wgt_9_517,
input [18:0] Wgt_9_518,
input [18:0] Wgt_9_519,
input [18:0] Wgt_9_520,
input [18:0] Wgt_9_521,
input [18:0] Wgt_9_522,
input [18:0] Wgt_9_523,
input [18:0] Wgt_9_524,
input [18:0] Wgt_9_525,
input [18:0] Wgt_9_526,
input [18:0] Wgt_9_527,
input [18:0] Wgt_9_528,
input [18:0] Wgt_9_529,
input [18:0] Wgt_9_530,
input [18:0] Wgt_9_531,
input [18:0] Wgt_9_532,
input [18:0] Wgt_9_533,
input [18:0] Wgt_9_534,
input [18:0] Wgt_9_535,
input [18:0] Wgt_9_536,
input [18:0] Wgt_9_537,
input [18:0] Wgt_9_538,
input [18:0] Wgt_9_539,
input [18:0] Wgt_9_540,
input [18:0] Wgt_9_541,
input [18:0] Wgt_9_542,
input [18:0] Wgt_9_543,
input [18:0] Wgt_9_544,
input [18:0] Wgt_9_545,
input [18:0] Wgt_9_546,
input [18:0] Wgt_9_547,
input [18:0] Wgt_9_548,
input [18:0] Wgt_9_549,
input [18:0] Wgt_9_550,
input [18:0] Wgt_9_551,
input [18:0] Wgt_9_552,
input [18:0] Wgt_9_553,
input [18:0] Wgt_9_554,
input [18:0] Wgt_9_555,
input [18:0] Wgt_9_556,
input [18:0] Wgt_9_557,
input [18:0] Wgt_9_558,
input [18:0] Wgt_9_559,
input [18:0] Wgt_9_560,
input [18:0] Wgt_9_561,
input [18:0] Wgt_9_562,
input [18:0] Wgt_9_563,
input [18:0] Wgt_9_564,
input [18:0] Wgt_9_565,
input [18:0] Wgt_9_566,
input [18:0] Wgt_9_567,
input [18:0] Wgt_9_568,
input [18:0] Wgt_9_569,
input [18:0] Wgt_9_570,
input [18:0] Wgt_9_571,
input [18:0] Wgt_9_572,
input [18:0] Wgt_9_573,
input [18:0] Wgt_9_574,
input [18:0] Wgt_9_575,
input [18:0] Wgt_9_576,
input [18:0] Wgt_9_577,
input [18:0] Wgt_9_578,
input [18:0] Wgt_9_579,
input [18:0] Wgt_9_580,
input [18:0] Wgt_9_581,
input [18:0] Wgt_9_582,
input [18:0] Wgt_9_583,
input [18:0] Wgt_9_584,
input [18:0] Wgt_9_585,
input [18:0] Wgt_9_586,
input [18:0] Wgt_9_587,
input [18:0] Wgt_9_588,
input [18:0] Wgt_9_589,
input [18:0] Wgt_9_590,
input [18:0] Wgt_9_591,
input [18:0] Wgt_9_592,
input [18:0] Wgt_9_593,
input [18:0] Wgt_9_594,
input [18:0] Wgt_9_595,
input [18:0] Wgt_9_596,
input [18:0] Wgt_9_597,
input [18:0] Wgt_9_598,
input [18:0] Wgt_9_599,
input [18:0] Wgt_9_600,
input [18:0] Wgt_9_601,
input [18:0] Wgt_9_602,
input [18:0] Wgt_9_603,
input [18:0] Wgt_9_604,
input [18:0] Wgt_9_605,
input [18:0] Wgt_9_606,
input [18:0] Wgt_9_607,
input [18:0] Wgt_9_608,
input [18:0] Wgt_9_609,
input [18:0] Wgt_9_610,
input [18:0] Wgt_9_611,
input [18:0] Wgt_9_612,
input [18:0] Wgt_9_613,
input [18:0] Wgt_9_614,
input [18:0] Wgt_9_615,
input [18:0] Wgt_9_616,
input [18:0] Wgt_9_617,
input [18:0] Wgt_9_618,
input [18:0] Wgt_9_619,
input [18:0] Wgt_9_620,
input [18:0] Wgt_9_621,
input [18:0] Wgt_9_622,
input [18:0] Wgt_9_623,
input [18:0] Wgt_9_624,
input [18:0] Wgt_9_625,
input [18:0] Wgt_9_626,
input [18:0] Wgt_9_627,
input [18:0] Wgt_9_628,
input [18:0] Wgt_9_629,
input [18:0] Wgt_9_630,
input [18:0] Wgt_9_631,
input [18:0] Wgt_9_632,
input [18:0] Wgt_9_633,
input [18:0] Wgt_9_634,
input [18:0] Wgt_9_635,
input [18:0] Wgt_9_636,
input [18:0] Wgt_9_637,
input [18:0] Wgt_9_638,
input [18:0] Wgt_9_639,
input [18:0] Wgt_9_640,
input [18:0] Wgt_9_641,
input [18:0] Wgt_9_642,
input [18:0] Wgt_9_643,
input [18:0] Wgt_9_644,
input [18:0] Wgt_9_645,
input [18:0] Wgt_9_646,
input [18:0] Wgt_9_647,
input [18:0] Wgt_9_648,
input [18:0] Wgt_9_649,
input [18:0] Wgt_9_650,
input [18:0] Wgt_9_651,
input [18:0] Wgt_9_652,
input [18:0] Wgt_9_653,
input [18:0] Wgt_9_654,
input [18:0] Wgt_9_655,
input [18:0] Wgt_9_656,
input [18:0] Wgt_9_657,
input [18:0] Wgt_9_658,
input [18:0] Wgt_9_659,
input [18:0] Wgt_9_660,
input [18:0] Wgt_9_661,
input [18:0] Wgt_9_662,
input [18:0] Wgt_9_663,
input [18:0] Wgt_9_664,
input [18:0] Wgt_9_665,
input [18:0] Wgt_9_666,
input [18:0] Wgt_9_667,
input [18:0] Wgt_9_668,
input [18:0] Wgt_9_669,
input [18:0] Wgt_9_670,
input [18:0] Wgt_9_671,
input [18:0] Wgt_9_672,
input [18:0] Wgt_9_673,
input [18:0] Wgt_9_674,
input [18:0] Wgt_9_675,
input [18:0] Wgt_9_676,
input [18:0] Wgt_9_677,
input [18:0] Wgt_9_678,
input [18:0] Wgt_9_679,
input [18:0] Wgt_9_680,
input [18:0] Wgt_9_681,
input [18:0] Wgt_9_682,
input [18:0] Wgt_9_683,
input [18:0] Wgt_9_684,
input [18:0] Wgt_9_685,
input [18:0] Wgt_9_686,
input [18:0] Wgt_9_687,
input [18:0] Wgt_9_688,
input [18:0] Wgt_9_689,
input [18:0] Wgt_9_690,
input [18:0] Wgt_9_691,
input [18:0] Wgt_9_692,
input [18:0] Wgt_9_693,
input [18:0] Wgt_9_694,
input [18:0] Wgt_9_695,
input [18:0] Wgt_9_696,
input [18:0] Wgt_9_697,
input [18:0] Wgt_9_698,
input [18:0] Wgt_9_699,
input [18:0] Wgt_9_700,
input [18:0] Wgt_9_701,
input [18:0] Wgt_9_702,
input [18:0] Wgt_9_703,
input [18:0] Wgt_9_704,
input [18:0] Wgt_9_705,
input [18:0] Wgt_9_706,
input [18:0] Wgt_9_707,
input [18:0] Wgt_9_708,
input [18:0] Wgt_9_709,
input [18:0] Wgt_9_710,
input [18:0] Wgt_9_711,
input [18:0] Wgt_9_712,
input [18:0] Wgt_9_713,
input [18:0] Wgt_9_714,
input [18:0] Wgt_9_715,
input [18:0] Wgt_9_716,
input [18:0] Wgt_9_717,
input [18:0] Wgt_9_718,
input [18:0] Wgt_9_719,
input [18:0] Wgt_9_720,
input [18:0] Wgt_9_721,
input [18:0] Wgt_9_722,
input [18:0] Wgt_9_723,
input [18:0] Wgt_9_724,
input [18:0] Wgt_9_725,
input [18:0] Wgt_9_726,
input [18:0] Wgt_9_727,
input [18:0] Wgt_9_728,
input [18:0] Wgt_9_729,
input [18:0] Wgt_9_730,
input [18:0] Wgt_9_731,
input [18:0] Wgt_9_732,
input [18:0] Wgt_9_733,
input [18:0] Wgt_9_734,
input [18:0] Wgt_9_735,
input [18:0] Wgt_9_736,
input [18:0] Wgt_9_737,
input [18:0] Wgt_9_738,
input [18:0] Wgt_9_739,
input [18:0] Wgt_9_740,
input [18:0] Wgt_9_741,
input [18:0] Wgt_9_742,
input [18:0] Wgt_9_743,
input [18:0] Wgt_9_744,
input [18:0] Wgt_9_745,
input [18:0] Wgt_9_746,
input [18:0] Wgt_9_747,
input [18:0] Wgt_9_748,
input [18:0] Wgt_9_749,
input [18:0] Wgt_9_750,
input [18:0] Wgt_9_751,
input [18:0] Wgt_9_752,
input [18:0] Wgt_9_753,
input [18:0] Wgt_9_754,
input [18:0] Wgt_9_755,
input [18:0] Wgt_9_756,
input [18:0] Wgt_9_757,
input [18:0] Wgt_9_758,
input [18:0] Wgt_9_759,
input [18:0] Wgt_9_760,
input [18:0] Wgt_9_761,
input [18:0] Wgt_9_762,
input [18:0] Wgt_9_763,
input [18:0] Wgt_9_764,
input [18:0] Wgt_9_765,
input [18:0] Wgt_9_766,
input [18:0] Wgt_9_767,
input [18:0] Wgt_9_768,
input [18:0] Wgt_9_769,
input [18:0] Wgt_9_770,
input [18:0] Wgt_9_771,
input [18:0] Wgt_9_772,
input [18:0] Wgt_9_773,
input [18:0] Wgt_9_774,
input [18:0] Wgt_9_775,
input [18:0] Wgt_9_776,
input [18:0] Wgt_9_777,
input [18:0] Wgt_9_778,
input [18:0] Wgt_9_779,
input [18:0] Wgt_9_780,
input [18:0] Wgt_9_781,
input [18:0] Wgt_9_782,
input [18:0] Wgt_9_783,
input [18:0] Wgt_9_784,
input [9:0] Pix_0,
input [9:0] Pix_1,
input [9:0] Pix_2,
input [9:0] Pix_3,
input [9:0] Pix_4,
input [9:0] Pix_5,
input [9:0] Pix_6,
input [9:0] Pix_7,
input [9:0] Pix_8,
input [9:0] Pix_9,
input [9:0] Pix_10,
input [9:0] Pix_11,
input [9:0] Pix_12,
input [9:0] Pix_13,
input [9:0] Pix_14,
input [9:0] Pix_15,
input [9:0] Pix_16,
input [9:0] Pix_17,
input [9:0] Pix_18,
input [9:0] Pix_19,
input [9:0] Pix_20,
input [9:0] Pix_21,
input [9:0] Pix_22,
input [9:0] Pix_23,
input [9:0] Pix_24,
input [9:0] Pix_25,
input [9:0] Pix_26,
input [9:0] Pix_27,
input [9:0] Pix_28,
input [9:0] Pix_29,
input [9:0] Pix_30,
input [9:0] Pix_31,
input [9:0] Pix_32,
input [9:0] Pix_33,
input [9:0] Pix_34,
input [9:0] Pix_35,
input [9:0] Pix_36,
input [9:0] Pix_37,
input [9:0] Pix_38,
input [9:0] Pix_39,
input [9:0] Pix_40,
input [9:0] Pix_41,
input [9:0] Pix_42,
input [9:0] Pix_43,
input [9:0] Pix_44,
input [9:0] Pix_45,
input [9:0] Pix_46,
input [9:0] Pix_47,
input [9:0] Pix_48,
input [9:0] Pix_49,
input [9:0] Pix_50,
input [9:0] Pix_51,
input [9:0] Pix_52,
input [9:0] Pix_53,
input [9:0] Pix_54,
input [9:0] Pix_55,
input [9:0] Pix_56,
input [9:0] Pix_57,
input [9:0] Pix_58,
input [9:0] Pix_59,
input [9:0] Pix_60,
input [9:0] Pix_61,
input [9:0] Pix_62,
input [9:0] Pix_63,
input [9:0] Pix_64,
input [9:0] Pix_65,
input [9:0] Pix_66,
input [9:0] Pix_67,
input [9:0] Pix_68,
input [9:0] Pix_69,
input [9:0] Pix_70,
input [9:0] Pix_71,
input [9:0] Pix_72,
input [9:0] Pix_73,
input [9:0] Pix_74,
input [9:0] Pix_75,
input [9:0] Pix_76,
input [9:0] Pix_77,
input [9:0] Pix_78,
input [9:0] Pix_79,
input [9:0] Pix_80,
input [9:0] Pix_81,
input [9:0] Pix_82,
input [9:0] Pix_83,
input [9:0] Pix_84,
input [9:0] Pix_85,
input [9:0] Pix_86,
input [9:0] Pix_87,
input [9:0] Pix_88,
input [9:0] Pix_89,
input [9:0] Pix_90,
input [9:0] Pix_91,
input [9:0] Pix_92,
input [9:0] Pix_93,
input [9:0] Pix_94,
input [9:0] Pix_95,
input [9:0] Pix_96,
input [9:0] Pix_97,
input [9:0] Pix_98,
input [9:0] Pix_99,
input [9:0] Pix_100,
input [9:0] Pix_101,
input [9:0] Pix_102,
input [9:0] Pix_103,
input [9:0] Pix_104,
input [9:0] Pix_105,
input [9:0] Pix_106,
input [9:0] Pix_107,
input [9:0] Pix_108,
input [9:0] Pix_109,
input [9:0] Pix_110,
input [9:0] Pix_111,
input [9:0] Pix_112,
input [9:0] Pix_113,
input [9:0] Pix_114,
input [9:0] Pix_115,
input [9:0] Pix_116,
input [9:0] Pix_117,
input [9:0] Pix_118,
input [9:0] Pix_119,
input [9:0] Pix_120,
input [9:0] Pix_121,
input [9:0] Pix_122,
input [9:0] Pix_123,
input [9:0] Pix_124,
input [9:0] Pix_125,
input [9:0] Pix_126,
input [9:0] Pix_127,
input [9:0] Pix_128,
input [9:0] Pix_129,
input [9:0] Pix_130,
input [9:0] Pix_131,
input [9:0] Pix_132,
input [9:0] Pix_133,
input [9:0] Pix_134,
input [9:0] Pix_135,
input [9:0] Pix_136,
input [9:0] Pix_137,
input [9:0] Pix_138,
input [9:0] Pix_139,
input [9:0] Pix_140,
input [9:0] Pix_141,
input [9:0] Pix_142,
input [9:0] Pix_143,
input [9:0] Pix_144,
input [9:0] Pix_145,
input [9:0] Pix_146,
input [9:0] Pix_147,
input [9:0] Pix_148,
input [9:0] Pix_149,
input [9:0] Pix_150,
input [9:0] Pix_151,
input [9:0] Pix_152,
input [9:0] Pix_153,
input [9:0] Pix_154,
input [9:0] Pix_155,
input [9:0] Pix_156,
input [9:0] Pix_157,
input [9:0] Pix_158,
input [9:0] Pix_159,
input [9:0] Pix_160,
input [9:0] Pix_161,
input [9:0] Pix_162,
input [9:0] Pix_163,
input [9:0] Pix_164,
input [9:0] Pix_165,
input [9:0] Pix_166,
input [9:0] Pix_167,
input [9:0] Pix_168,
input [9:0] Pix_169,
input [9:0] Pix_170,
input [9:0] Pix_171,
input [9:0] Pix_172,
input [9:0] Pix_173,
input [9:0] Pix_174,
input [9:0] Pix_175,
input [9:0] Pix_176,
input [9:0] Pix_177,
input [9:0] Pix_178,
input [9:0] Pix_179,
input [9:0] Pix_180,
input [9:0] Pix_181,
input [9:0] Pix_182,
input [9:0] Pix_183,
input [9:0] Pix_184,
input [9:0] Pix_185,
input [9:0] Pix_186,
input [9:0] Pix_187,
input [9:0] Pix_188,
input [9:0] Pix_189,
input [9:0] Pix_190,
input [9:0] Pix_191,
input [9:0] Pix_192,
input [9:0] Pix_193,
input [9:0] Pix_194,
input [9:0] Pix_195,
input [9:0] Pix_196,
input [9:0] Pix_197,
input [9:0] Pix_198,
input [9:0] Pix_199,
input [9:0] Pix_200,
input [9:0] Pix_201,
input [9:0] Pix_202,
input [9:0] Pix_203,
input [9:0] Pix_204,
input [9:0] Pix_205,
input [9:0] Pix_206,
input [9:0] Pix_207,
input [9:0] Pix_208,
input [9:0] Pix_209,
input [9:0] Pix_210,
input [9:0] Pix_211,
input [9:0] Pix_212,
input [9:0] Pix_213,
input [9:0] Pix_214,
input [9:0] Pix_215,
input [9:0] Pix_216,
input [9:0] Pix_217,
input [9:0] Pix_218,
input [9:0] Pix_219,
input [9:0] Pix_220,
input [9:0] Pix_221,
input [9:0] Pix_222,
input [9:0] Pix_223,
input [9:0] Pix_224,
input [9:0] Pix_225,
input [9:0] Pix_226,
input [9:0] Pix_227,
input [9:0] Pix_228,
input [9:0] Pix_229,
input [9:0] Pix_230,
input [9:0] Pix_231,
input [9:0] Pix_232,
input [9:0] Pix_233,
input [9:0] Pix_234,
input [9:0] Pix_235,
input [9:0] Pix_236,
input [9:0] Pix_237,
input [9:0] Pix_238,
input [9:0] Pix_239,
input [9:0] Pix_240,
input [9:0] Pix_241,
input [9:0] Pix_242,
input [9:0] Pix_243,
input [9:0] Pix_244,
input [9:0] Pix_245,
input [9:0] Pix_246,
input [9:0] Pix_247,
input [9:0] Pix_248,
input [9:0] Pix_249,
input [9:0] Pix_250,
input [9:0] Pix_251,
input [9:0] Pix_252,
input [9:0] Pix_253,
input [9:0] Pix_254,
input [9:0] Pix_255,
input [9:0] Pix_256,
input [9:0] Pix_257,
input [9:0] Pix_258,
input [9:0] Pix_259,
input [9:0] Pix_260,
input [9:0] Pix_261,
input [9:0] Pix_262,
input [9:0] Pix_263,
input [9:0] Pix_264,
input [9:0] Pix_265,
input [9:0] Pix_266,
input [9:0] Pix_267,
input [9:0] Pix_268,
input [9:0] Pix_269,
input [9:0] Pix_270,
input [9:0] Pix_271,
input [9:0] Pix_272,
input [9:0] Pix_273,
input [9:0] Pix_274,
input [9:0] Pix_275,
input [9:0] Pix_276,
input [9:0] Pix_277,
input [9:0] Pix_278,
input [9:0] Pix_279,
input [9:0] Pix_280,
input [9:0] Pix_281,
input [9:0] Pix_282,
input [9:0] Pix_283,
input [9:0] Pix_284,
input [9:0] Pix_285,
input [9:0] Pix_286,
input [9:0] Pix_287,
input [9:0] Pix_288,
input [9:0] Pix_289,
input [9:0] Pix_290,
input [9:0] Pix_291,
input [9:0] Pix_292,
input [9:0] Pix_293,
input [9:0] Pix_294,
input [9:0] Pix_295,
input [9:0] Pix_296,
input [9:0] Pix_297,
input [9:0] Pix_298,
input [9:0] Pix_299,
input [9:0] Pix_300,
input [9:0] Pix_301,
input [9:0] Pix_302,
input [9:0] Pix_303,
input [9:0] Pix_304,
input [9:0] Pix_305,
input [9:0] Pix_306,
input [9:0] Pix_307,
input [9:0] Pix_308,
input [9:0] Pix_309,
input [9:0] Pix_310,
input [9:0] Pix_311,
input [9:0] Pix_312,
input [9:0] Pix_313,
input [9:0] Pix_314,
input [9:0] Pix_315,
input [9:0] Pix_316,
input [9:0] Pix_317,
input [9:0] Pix_318,
input [9:0] Pix_319,
input [9:0] Pix_320,
input [9:0] Pix_321,
input [9:0] Pix_322,
input [9:0] Pix_323,
input [9:0] Pix_324,
input [9:0] Pix_325,
input [9:0] Pix_326,
input [9:0] Pix_327,
input [9:0] Pix_328,
input [9:0] Pix_329,
input [9:0] Pix_330,
input [9:0] Pix_331,
input [9:0] Pix_332,
input [9:0] Pix_333,
input [9:0] Pix_334,
input [9:0] Pix_335,
input [9:0] Pix_336,
input [9:0] Pix_337,
input [9:0] Pix_338,
input [9:0] Pix_339,
input [9:0] Pix_340,
input [9:0] Pix_341,
input [9:0] Pix_342,
input [9:0] Pix_343,
input [9:0] Pix_344,
input [9:0] Pix_345,
input [9:0] Pix_346,
input [9:0] Pix_347,
input [9:0] Pix_348,
input [9:0] Pix_349,
input [9:0] Pix_350,
input [9:0] Pix_351,
input [9:0] Pix_352,
input [9:0] Pix_353,
input [9:0] Pix_354,
input [9:0] Pix_355,
input [9:0] Pix_356,
input [9:0] Pix_357,
input [9:0] Pix_358,
input [9:0] Pix_359,
input [9:0] Pix_360,
input [9:0] Pix_361,
input [9:0] Pix_362,
input [9:0] Pix_363,
input [9:0] Pix_364,
input [9:0] Pix_365,
input [9:0] Pix_366,
input [9:0] Pix_367,
input [9:0] Pix_368,
input [9:0] Pix_369,
input [9:0] Pix_370,
input [9:0] Pix_371,
input [9:0] Pix_372,
input [9:0] Pix_373,
input [9:0] Pix_374,
input [9:0] Pix_375,
input [9:0] Pix_376,
input [9:0] Pix_377,
input [9:0] Pix_378,
input [9:0] Pix_379,
input [9:0] Pix_380,
input [9:0] Pix_381,
input [9:0] Pix_382,
input [9:0] Pix_383,
input [9:0] Pix_384,
input [9:0] Pix_385,
input [9:0] Pix_386,
input [9:0] Pix_387,
input [9:0] Pix_388,
input [9:0] Pix_389,
input [9:0] Pix_390,
input [9:0] Pix_391,
input [9:0] Pix_392,
input [9:0] Pix_393,
input [9:0] Pix_394,
input [9:0] Pix_395,
input [9:0] Pix_396,
input [9:0] Pix_397,
input [9:0] Pix_398,
input [9:0] Pix_399,
input [9:0] Pix_400,
input [9:0] Pix_401,
input [9:0] Pix_402,
input [9:0] Pix_403,
input [9:0] Pix_404,
input [9:0] Pix_405,
input [9:0] Pix_406,
input [9:0] Pix_407,
input [9:0] Pix_408,
input [9:0] Pix_409,
input [9:0] Pix_410,
input [9:0] Pix_411,
input [9:0] Pix_412,
input [9:0] Pix_413,
input [9:0] Pix_414,
input [9:0] Pix_415,
input [9:0] Pix_416,
input [9:0] Pix_417,
input [9:0] Pix_418,
input [9:0] Pix_419,
input [9:0] Pix_420,
input [9:0] Pix_421,
input [9:0] Pix_422,
input [9:0] Pix_423,
input [9:0] Pix_424,
input [9:0] Pix_425,
input [9:0] Pix_426,
input [9:0] Pix_427,
input [9:0] Pix_428,
input [9:0] Pix_429,
input [9:0] Pix_430,
input [9:0] Pix_431,
input [9:0] Pix_432,
input [9:0] Pix_433,
input [9:0] Pix_434,
input [9:0] Pix_435,
input [9:0] Pix_436,
input [9:0] Pix_437,
input [9:0] Pix_438,
input [9:0] Pix_439,
input [9:0] Pix_440,
input [9:0] Pix_441,
input [9:0] Pix_442,
input [9:0] Pix_443,
input [9:0] Pix_444,
input [9:0] Pix_445,
input [9:0] Pix_446,
input [9:0] Pix_447,
input [9:0] Pix_448,
input [9:0] Pix_449,
input [9:0] Pix_450,
input [9:0] Pix_451,
input [9:0] Pix_452,
input [9:0] Pix_453,
input [9:0] Pix_454,
input [9:0] Pix_455,
input [9:0] Pix_456,
input [9:0] Pix_457,
input [9:0] Pix_458,
input [9:0] Pix_459,
input [9:0] Pix_460,
input [9:0] Pix_461,
input [9:0] Pix_462,
input [9:0] Pix_463,
input [9:0] Pix_464,
input [9:0] Pix_465,
input [9:0] Pix_466,
input [9:0] Pix_467,
input [9:0] Pix_468,
input [9:0] Pix_469,
input [9:0] Pix_470,
input [9:0] Pix_471,
input [9:0] Pix_472,
input [9:0] Pix_473,
input [9:0] Pix_474,
input [9:0] Pix_475,
input [9:0] Pix_476,
input [9:0] Pix_477,
input [9:0] Pix_478,
input [9:0] Pix_479,
input [9:0] Pix_480,
input [9:0] Pix_481,
input [9:0] Pix_482,
input [9:0] Pix_483,
input [9:0] Pix_484,
input [9:0] Pix_485,
input [9:0] Pix_486,
input [9:0] Pix_487,
input [9:0] Pix_488,
input [9:0] Pix_489,
input [9:0] Pix_490,
input [9:0] Pix_491,
input [9:0] Pix_492,
input [9:0] Pix_493,
input [9:0] Pix_494,
input [9:0] Pix_495,
input [9:0] Pix_496,
input [9:0] Pix_497,
input [9:0] Pix_498,
input [9:0] Pix_499,
input [9:0] Pix_500,
input [9:0] Pix_501,
input [9:0] Pix_502,
input [9:0] Pix_503,
input [9:0] Pix_504,
input [9:0] Pix_505,
input [9:0] Pix_506,
input [9:0] Pix_507,
input [9:0] Pix_508,
input [9:0] Pix_509,
input [9:0] Pix_510,
input [9:0] Pix_511,
input [9:0] Pix_512,
input [9:0] Pix_513,
input [9:0] Pix_514,
input [9:0] Pix_515,
input [9:0] Pix_516,
input [9:0] Pix_517,
input [9:0] Pix_518,
input [9:0] Pix_519,
input [9:0] Pix_520,
input [9:0] Pix_521,
input [9:0] Pix_522,
input [9:0] Pix_523,
input [9:0] Pix_524,
input [9:0] Pix_525,
input [9:0] Pix_526,
input [9:0] Pix_527,
input [9:0] Pix_528,
input [9:0] Pix_529,
input [9:0] Pix_530,
input [9:0] Pix_531,
input [9:0] Pix_532,
input [9:0] Pix_533,
input [9:0] Pix_534,
input [9:0] Pix_535,
input [9:0] Pix_536,
input [9:0] Pix_537,
input [9:0] Pix_538,
input [9:0] Pix_539,
input [9:0] Pix_540,
input [9:0] Pix_541,
input [9:0] Pix_542,
input [9:0] Pix_543,
input [9:0] Pix_544,
input [9:0] Pix_545,
input [9:0] Pix_546,
input [9:0] Pix_547,
input [9:0] Pix_548,
input [9:0] Pix_549,
input [9:0] Pix_550,
input [9:0] Pix_551,
input [9:0] Pix_552,
input [9:0] Pix_553,
input [9:0] Pix_554,
input [9:0] Pix_555,
input [9:0] Pix_556,
input [9:0] Pix_557,
input [9:0] Pix_558,
input [9:0] Pix_559,
input [9:0] Pix_560,
input [9:0] Pix_561,
input [9:0] Pix_562,
input [9:0] Pix_563,
input [9:0] Pix_564,
input [9:0] Pix_565,
input [9:0] Pix_566,
input [9:0] Pix_567,
input [9:0] Pix_568,
input [9:0] Pix_569,
input [9:0] Pix_570,
input [9:0] Pix_571,
input [9:0] Pix_572,
input [9:0] Pix_573,
input [9:0] Pix_574,
input [9:0] Pix_575,
input [9:0] Pix_576,
input [9:0] Pix_577,
input [9:0] Pix_578,
input [9:0] Pix_579,
input [9:0] Pix_580,
input [9:0] Pix_581,
input [9:0] Pix_582,
input [9:0] Pix_583,
input [9:0] Pix_584,
input [9:0] Pix_585,
input [9:0] Pix_586,
input [9:0] Pix_587,
input [9:0] Pix_588,
input [9:0] Pix_589,
input [9:0] Pix_590,
input [9:0] Pix_591,
input [9:0] Pix_592,
input [9:0] Pix_593,
input [9:0] Pix_594,
input [9:0] Pix_595,
input [9:0] Pix_596,
input [9:0] Pix_597,
input [9:0] Pix_598,
input [9:0] Pix_599,
input [9:0] Pix_600,
input [9:0] Pix_601,
input [9:0] Pix_602,
input [9:0] Pix_603,
input [9:0] Pix_604,
input [9:0] Pix_605,
input [9:0] Pix_606,
input [9:0] Pix_607,
input [9:0] Pix_608,
input [9:0] Pix_609,
input [9:0] Pix_610,
input [9:0] Pix_611,
input [9:0] Pix_612,
input [9:0] Pix_613,
input [9:0] Pix_614,
input [9:0] Pix_615,
input [9:0] Pix_616,
input [9:0] Pix_617,
input [9:0] Pix_618,
input [9:0] Pix_619,
input [9:0] Pix_620,
input [9:0] Pix_621,
input [9:0] Pix_622,
input [9:0] Pix_623,
input [9:0] Pix_624,
input [9:0] Pix_625,
input [9:0] Pix_626,
input [9:0] Pix_627,
input [9:0] Pix_628,
input [9:0] Pix_629,
input [9:0] Pix_630,
input [9:0] Pix_631,
input [9:0] Pix_632,
input [9:0] Pix_633,
input [9:0] Pix_634,
input [9:0] Pix_635,
input [9:0] Pix_636,
input [9:0] Pix_637,
input [9:0] Pix_638,
input [9:0] Pix_639,
input [9:0] Pix_640,
input [9:0] Pix_641,
input [9:0] Pix_642,
input [9:0] Pix_643,
input [9:0] Pix_644,
input [9:0] Pix_645,
input [9:0] Pix_646,
input [9:0] Pix_647,
input [9:0] Pix_648,
input [9:0] Pix_649,
input [9:0] Pix_650,
input [9:0] Pix_651,
input [9:0] Pix_652,
input [9:0] Pix_653,
input [9:0] Pix_654,
input [9:0] Pix_655,
input [9:0] Pix_656,
input [9:0] Pix_657,
input [9:0] Pix_658,
input [9:0] Pix_659,
input [9:0] Pix_660,
input [9:0] Pix_661,
input [9:0] Pix_662,
input [9:0] Pix_663,
input [9:0] Pix_664,
input [9:0] Pix_665,
input [9:0] Pix_666,
input [9:0] Pix_667,
input [9:0] Pix_668,
input [9:0] Pix_669,
input [9:0] Pix_670,
input [9:0] Pix_671,
input [9:0] Pix_672,
input [9:0] Pix_673,
input [9:0] Pix_674,
input [9:0] Pix_675,
input [9:0] Pix_676,
input [9:0] Pix_677,
input [9:0] Pix_678,
input [9:0] Pix_679,
input [9:0] Pix_680,
input [9:0] Pix_681,
input [9:0] Pix_682,
input [9:0] Pix_683,
input [9:0] Pix_684,
input [9:0] Pix_685,
input [9:0] Pix_686,
input [9:0] Pix_687,
input [9:0] Pix_688,
input [9:0] Pix_689,
input [9:0] Pix_690,
input [9:0] Pix_691,
input [9:0] Pix_692,
input [9:0] Pix_693,
input [9:0] Pix_694,
input [9:0] Pix_695,
input [9:0] Pix_696,
input [9:0] Pix_697,
input [9:0] Pix_698,
input [9:0] Pix_699,
input [9:0] Pix_700,
input [9:0] Pix_701,
input [9:0] Pix_702,
input [9:0] Pix_703,
input [9:0] Pix_704,
input [9:0] Pix_705,
input [9:0] Pix_706,
input [9:0] Pix_707,
input [9:0] Pix_708,
input [9:0] Pix_709,
input [9:0] Pix_710,
input [9:0] Pix_711,
input [9:0] Pix_712,
input [9:0] Pix_713,
input [9:0] Pix_714,
input [9:0] Pix_715,
input [9:0] Pix_716,
input [9:0] Pix_717,
input [9:0] Pix_718,
input [9:0] Pix_719,
input [9:0] Pix_720,
input [9:0] Pix_721,
input [9:0] Pix_722,
input [9:0] Pix_723,
input [9:0] Pix_724,
input [9:0] Pix_725,
input [9:0] Pix_726,
input [9:0] Pix_727,
input [9:0] Pix_728,
input [9:0] Pix_729,
input [9:0] Pix_730,
input [9:0] Pix_731,
input [9:0] Pix_732,
input [9:0] Pix_733,
input [9:0] Pix_734,
input [9:0] Pix_735,
input [9:0] Pix_736,
input [9:0] Pix_737,
input [9:0] Pix_738,
input [9:0] Pix_739,
input [9:0] Pix_740,
input [9:0] Pix_741,
input [9:0] Pix_742,
input [9:0] Pix_743,
input [9:0] Pix_744,
input [9:0] Pix_745,
input [9:0] Pix_746,
input [9:0] Pix_747,
input [9:0] Pix_748,
input [9:0] Pix_749,
input [9:0] Pix_750,
input [9:0] Pix_751,
input [9:0] Pix_752,
input [9:0] Pix_753,
input [9:0] Pix_754,
input [9:0] Pix_755,
input [9:0] Pix_756,
input [9:0] Pix_757,
input [9:0] Pix_758,
input [9:0] Pix_759,
input [9:0] Pix_760,
input [9:0] Pix_761,
input [9:0] Pix_762,
input [9:0] Pix_763,
input [9:0] Pix_764,
input [9:0] Pix_765,
input [9:0] Pix_766,
input [9:0] Pix_767,
input [9:0] Pix_768,
input [9:0] Pix_769,
input [9:0] Pix_770,
input [9:0] Pix_771,
input [9:0] Pix_772,
input [9:0] Pix_773,
input [9:0] Pix_774,
input [9:0] Pix_775,
input [9:0] Pix_776,
input [9:0] Pix_777,
input [9:0] Pix_778,
input [9:0] Pix_779,
input [9:0] Pix_780,
input [9:0] Pix_781,
input [9:0] Pix_782,
input [9:0] Pix_783,
input [9:0] Pix_784,
output [3:0] Image_Number,
output Output_Valid
);

reg[9:0] PixelsStore[0:784];
reg[18:0] WeightsStore0[0:784];
reg[18:0] WeightsStore1[0:784];
reg[18:0] WeightsStore2[0:784];
reg[18:0] WeightsStore3[0:784];
reg[18:0] WeightsStore4[0:784];
reg[18:0] WeightsStore5[0:784];
reg[18:0] WeightsStore6[0:784];
reg[18:0] WeightsStore7[0:784];
reg[18:0] WeightsStore8[0:784];
reg[18:0] WeightsStore9[0:784];
reg[31:0] switchCounter;
reg ready;
reg internalReset;
wire[259:0] value;

assign Output_Valid = ready;

DotProduct784 DP0(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore0[0]),
	.Weight1(WeightsStore0[1]),
	.Weight2(WeightsStore0[2]),
	.Weight3(WeightsStore0[3]),
	.Weight4(WeightsStore0[4]),
	.Weight5(WeightsStore0[5]),
	.Weight6(WeightsStore0[6]),
	.Weight7(WeightsStore0[7]),
	.Weight8(WeightsStore0[8]),
	.Weight9(WeightsStore0[9]),
	.Weight10(WeightsStore0[10]),
	.Weight11(WeightsStore0[11]),
	.Weight12(WeightsStore0[12]),
	.Weight13(WeightsStore0[13]),
	.Weight14(WeightsStore0[14]),
	.Weight15(WeightsStore0[15]),
	.Weight16(WeightsStore0[16]),
	.Weight17(WeightsStore0[17]),
	.Weight18(WeightsStore0[18]),
	.Weight19(WeightsStore0[19]),
	.Weight20(WeightsStore0[20]),
	.Weight21(WeightsStore0[21]),
	.Weight22(WeightsStore0[22]),
	.Weight23(WeightsStore0[23]),
	.Weight24(WeightsStore0[24]),
	.Weight25(WeightsStore0[25]),
	.Weight26(WeightsStore0[26]),
	.Weight27(WeightsStore0[27]),
	.WeightBias(WeightsStore0[784]),
	.value(value[25:0])
	);
DotProduct784 DP1(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore1[0]),
	.Weight1(WeightsStore1[1]),
	.Weight2(WeightsStore1[2]),
	.Weight3(WeightsStore1[3]),
	.Weight4(WeightsStore1[4]),
	.Weight5(WeightsStore1[5]),
	.Weight6(WeightsStore1[6]),
	.Weight7(WeightsStore1[7]),
	.Weight8(WeightsStore1[8]),
	.Weight9(WeightsStore1[9]),
	.Weight10(WeightsStore1[10]),
	.Weight11(WeightsStore1[11]),
	.Weight12(WeightsStore1[12]),
	.Weight13(WeightsStore1[13]),
	.Weight14(WeightsStore1[14]),
	.Weight15(WeightsStore1[15]),
	.Weight16(WeightsStore1[16]),
	.Weight17(WeightsStore1[17]),
	.Weight18(WeightsStore1[18]),
	.Weight19(WeightsStore1[19]),
	.Weight20(WeightsStore1[20]),
	.Weight21(WeightsStore1[21]),
	.Weight22(WeightsStore1[22]),
	.Weight23(WeightsStore1[23]),
	.Weight24(WeightsStore1[24]),
	.Weight25(WeightsStore1[25]),
	.Weight26(WeightsStore1[26]),
	.Weight27(WeightsStore1[27]),
	.WeightBias(WeightsStore1[784]),
	.value(value[51:26])
	);
DotProduct784 DP2(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore2[0]),
	.Weight1(WeightsStore2[1]),
	.Weight2(WeightsStore2[2]),
	.Weight3(WeightsStore2[3]),
	.Weight4(WeightsStore2[4]),
	.Weight5(WeightsStore2[5]),
	.Weight6(WeightsStore2[6]),
	.Weight7(WeightsStore2[7]),
	.Weight8(WeightsStore2[8]),
	.Weight9(WeightsStore2[9]),
	.Weight10(WeightsStore2[10]),
	.Weight11(WeightsStore2[11]),
	.Weight12(WeightsStore2[12]),
	.Weight13(WeightsStore2[13]),
	.Weight14(WeightsStore2[14]),
	.Weight15(WeightsStore2[15]),
	.Weight16(WeightsStore2[16]),
	.Weight17(WeightsStore2[17]),
	.Weight18(WeightsStore2[18]),
	.Weight19(WeightsStore2[19]),
	.Weight20(WeightsStore2[20]),
	.Weight21(WeightsStore2[21]),
	.Weight22(WeightsStore2[22]),
	.Weight23(WeightsStore2[23]),
	.Weight24(WeightsStore2[24]),
	.Weight25(WeightsStore2[25]),
	.Weight26(WeightsStore2[26]),
	.Weight27(WeightsStore2[27]),
	.WeightBias(WeightsStore2[784]),
	.value(value[77:52])
	);
DotProduct784 DP3(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore3[0]),
	.Weight1(WeightsStore3[1]),
	.Weight2(WeightsStore3[2]),
	.Weight3(WeightsStore3[3]),
	.Weight4(WeightsStore3[4]),
	.Weight5(WeightsStore3[5]),
	.Weight6(WeightsStore3[6]),
	.Weight7(WeightsStore3[7]),
	.Weight8(WeightsStore3[8]),
	.Weight9(WeightsStore3[9]),
	.Weight10(WeightsStore3[10]),
	.Weight11(WeightsStore3[11]),
	.Weight12(WeightsStore3[12]),
	.Weight13(WeightsStore3[13]),
	.Weight14(WeightsStore3[14]),
	.Weight15(WeightsStore3[15]),
	.Weight16(WeightsStore3[16]),
	.Weight17(WeightsStore3[17]),
	.Weight18(WeightsStore3[18]),
	.Weight19(WeightsStore3[19]),
	.Weight20(WeightsStore3[20]),
	.Weight21(WeightsStore3[21]),
	.Weight22(WeightsStore3[22]),
	.Weight23(WeightsStore3[23]),
	.Weight24(WeightsStore3[24]),
	.Weight25(WeightsStore3[25]),
	.Weight26(WeightsStore3[26]),
	.Weight27(WeightsStore3[27]),
	.WeightBias(WeightsStore3[784]),
	.value(value[103:78])
	);
DotProduct784 DP4(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore4[0]),
	.Weight1(WeightsStore4[1]),
	.Weight2(WeightsStore4[2]),
	.Weight3(WeightsStore4[3]),
	.Weight4(WeightsStore4[4]),
	.Weight5(WeightsStore4[5]),
	.Weight6(WeightsStore4[6]),
	.Weight7(WeightsStore4[7]),
	.Weight8(WeightsStore4[8]),
	.Weight9(WeightsStore4[9]),
	.Weight10(WeightsStore4[10]),
	.Weight11(WeightsStore4[11]),
	.Weight12(WeightsStore4[12]),
	.Weight13(WeightsStore4[13]),
	.Weight14(WeightsStore4[14]),
	.Weight15(WeightsStore4[15]),
	.Weight16(WeightsStore4[16]),
	.Weight17(WeightsStore4[17]),
	.Weight18(WeightsStore4[18]),
	.Weight19(WeightsStore4[19]),
	.Weight20(WeightsStore4[20]),
	.Weight21(WeightsStore4[21]),
	.Weight22(WeightsStore4[22]),
	.Weight23(WeightsStore4[23]),
	.Weight24(WeightsStore4[24]),
	.Weight25(WeightsStore4[25]),
	.Weight26(WeightsStore4[26]),
	.Weight27(WeightsStore4[27]),
	.WeightBias(WeightsStore4[784]),
	.value(value[129:104])
	);
DotProduct784 DP5(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore5[0]),
	.Weight1(WeightsStore5[1]),
	.Weight2(WeightsStore5[2]),
	.Weight3(WeightsStore5[3]),
	.Weight4(WeightsStore5[4]),
	.Weight5(WeightsStore5[5]),
	.Weight6(WeightsStore5[6]),
	.Weight7(WeightsStore5[7]),
	.Weight8(WeightsStore5[8]),
	.Weight9(WeightsStore5[9]),
	.Weight10(WeightsStore5[10]),
	.Weight11(WeightsStore5[11]),
	.Weight12(WeightsStore5[12]),
	.Weight13(WeightsStore5[13]),
	.Weight14(WeightsStore5[14]),
	.Weight15(WeightsStore5[15]),
	.Weight16(WeightsStore5[16]),
	.Weight17(WeightsStore5[17]),
	.Weight18(WeightsStore5[18]),
	.Weight19(WeightsStore5[19]),
	.Weight20(WeightsStore5[20]),
	.Weight21(WeightsStore5[21]),
	.Weight22(WeightsStore5[22]),
	.Weight23(WeightsStore5[23]),
	.Weight24(WeightsStore5[24]),
	.Weight25(WeightsStore5[25]),
	.Weight26(WeightsStore5[26]),
	.Weight27(WeightsStore5[27]),
	.WeightBias(WeightsStore5[784]),
	.value(value[155:130])
	);
DotProduct784 DP6(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore6[0]),
	.Weight1(WeightsStore6[1]),
	.Weight2(WeightsStore6[2]),
	.Weight3(WeightsStore6[3]),
	.Weight4(WeightsStore6[4]),
	.Weight5(WeightsStore6[5]),
	.Weight6(WeightsStore6[6]),
	.Weight7(WeightsStore6[7]),
	.Weight8(WeightsStore6[8]),
	.Weight9(WeightsStore6[9]),
	.Weight10(WeightsStore6[10]),
	.Weight11(WeightsStore6[11]),
	.Weight12(WeightsStore6[12]),
	.Weight13(WeightsStore6[13]),
	.Weight14(WeightsStore6[14]),
	.Weight15(WeightsStore6[15]),
	.Weight16(WeightsStore6[16]),
	.Weight17(WeightsStore6[17]),
	.Weight18(WeightsStore6[18]),
	.Weight19(WeightsStore6[19]),
	.Weight20(WeightsStore6[20]),
	.Weight21(WeightsStore6[21]),
	.Weight22(WeightsStore6[22]),
	.Weight23(WeightsStore6[23]),
	.Weight24(WeightsStore6[24]),
	.Weight25(WeightsStore6[25]),
	.Weight26(WeightsStore6[26]),
	.Weight27(WeightsStore6[27]),
	.WeightBias(WeightsStore6[784]),
	.value(value[181:156])
	);
DotProduct784 DP7(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore7[0]),
	.Weight1(WeightsStore7[1]),
	.Weight2(WeightsStore7[2]),
	.Weight3(WeightsStore7[3]),
	.Weight4(WeightsStore7[4]),
	.Weight5(WeightsStore7[5]),
	.Weight6(WeightsStore7[6]),
	.Weight7(WeightsStore7[7]),
	.Weight8(WeightsStore7[8]),
	.Weight9(WeightsStore7[9]),
	.Weight10(WeightsStore7[10]),
	.Weight11(WeightsStore7[11]),
	.Weight12(WeightsStore7[12]),
	.Weight13(WeightsStore7[13]),
	.Weight14(WeightsStore7[14]),
	.Weight15(WeightsStore7[15]),
	.Weight16(WeightsStore7[16]),
	.Weight17(WeightsStore7[17]),
	.Weight18(WeightsStore7[18]),
	.Weight19(WeightsStore7[19]),
	.Weight20(WeightsStore7[20]),
	.Weight21(WeightsStore7[21]),
	.Weight22(WeightsStore7[22]),
	.Weight23(WeightsStore7[23]),
	.Weight24(WeightsStore7[24]),
	.Weight25(WeightsStore7[25]),
	.Weight26(WeightsStore7[26]),
	.Weight27(WeightsStore7[27]),
	.WeightBias(WeightsStore7[784]),
	.value(value[207:182])
	);
DotProduct784 DP8(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore8[0]),
	.Weight1(WeightsStore8[1]),
	.Weight2(WeightsStore8[2]),
	.Weight3(WeightsStore8[3]),
	.Weight4(WeightsStore8[4]),
	.Weight5(WeightsStore8[5]),
	.Weight6(WeightsStore8[6]),
	.Weight7(WeightsStore8[7]),
	.Weight8(WeightsStore8[8]),
	.Weight9(WeightsStore8[9]),
	.Weight10(WeightsStore8[10]),
	.Weight11(WeightsStore8[11]),
	.Weight12(WeightsStore8[12]),
	.Weight13(WeightsStore8[13]),
	.Weight14(WeightsStore8[14]),
	.Weight15(WeightsStore8[15]),
	.Weight16(WeightsStore8[16]),
	.Weight17(WeightsStore8[17]),
	.Weight18(WeightsStore8[18]),
	.Weight19(WeightsStore8[19]),
	.Weight20(WeightsStore8[20]),
	.Weight21(WeightsStore8[21]),
	.Weight22(WeightsStore8[22]),
	.Weight23(WeightsStore8[23]),
	.Weight24(WeightsStore8[24]),
	.Weight25(WeightsStore8[25]),
	.Weight26(WeightsStore8[26]),
	.Weight27(WeightsStore8[27]),
	.WeightBias(WeightsStore8[784]),
	.value(value[233:208])
	);
DotProduct784 DP9(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore9[0]),
	.Weight1(WeightsStore9[1]),
	.Weight2(WeightsStore9[2]),
	.Weight3(WeightsStore9[3]),
	.Weight4(WeightsStore9[4]),
	.Weight5(WeightsStore9[5]),
	.Weight6(WeightsStore9[6]),
	.Weight7(WeightsStore9[7]),
	.Weight8(WeightsStore9[8]),
	.Weight9(WeightsStore9[9]),
	.Weight10(WeightsStore9[10]),
	.Weight11(WeightsStore9[11]),
	.Weight12(WeightsStore9[12]),
	.Weight13(WeightsStore9[13]),
	.Weight14(WeightsStore9[14]),
	.Weight15(WeightsStore9[15]),
	.Weight16(WeightsStore9[16]),
	.Weight17(WeightsStore9[17]),
	.Weight18(WeightsStore9[18]),
	.Weight19(WeightsStore9[19]),
	.Weight20(WeightsStore9[20]),
	.Weight21(WeightsStore9[21]),
	.Weight22(WeightsStore9[22]),
	.Weight23(WeightsStore9[23]),
	.Weight24(WeightsStore9[24]),
	.Weight25(WeightsStore9[25]),
	.Weight26(WeightsStore9[26]),
	.Weight27(WeightsStore9[27]),
	.WeightBias(WeightsStore9[784]),
	.value(value[259:234])
	);
Max max(.GlobalReset(internalReset),
	.Num(value),
	.Index(Image_Number)
	);

always@(posedge clk)begin
	if(GlobalReset == 1'b0)begin
		switchCounter <= 32'd0;
		ready <= 1'b0;
		internalReset = 1'b0;
		PixelsStore[0] <= 10'd0;
		PixelsStore[1] <= 10'd0;
		PixelsStore[2] <= 10'd0;
		PixelsStore[3] <= 10'd0;
		PixelsStore[4] <= 10'd0;
		PixelsStore[5] <= 10'd0;
		PixelsStore[6] <= 10'd0;
		PixelsStore[7] <= 10'd0;
		PixelsStore[8] <= 10'd0;
		PixelsStore[9] <= 10'd0;
		PixelsStore[10] <= 10'd0;
		PixelsStore[11] <= 10'd0;
		PixelsStore[12] <= 10'd0;
		PixelsStore[13] <= 10'd0;
		PixelsStore[14] <= 10'd0;
		PixelsStore[15] <= 10'd0;
		PixelsStore[16] <= 10'd0;
		PixelsStore[17] <= 10'd0;
		PixelsStore[18] <= 10'd0;
		PixelsStore[19] <= 10'd0;
		PixelsStore[20] <= 10'd0;
		PixelsStore[21] <= 10'd0;
		PixelsStore[22] <= 10'd0;
		PixelsStore[23] <= 10'd0;
		PixelsStore[24] <= 10'd0;
		PixelsStore[25] <= 10'd0;
		PixelsStore[26] <= 10'd0;
		PixelsStore[27] <= 10'd0;
		PixelsStore[28] <= 10'd0;
		PixelsStore[29] <= 10'd0;
		PixelsStore[30] <= 10'd0;
		PixelsStore[31] <= 10'd0;
		PixelsStore[32] <= 10'd0;
		PixelsStore[33] <= 10'd0;
		PixelsStore[34] <= 10'd0;
		PixelsStore[35] <= 10'd0;
		PixelsStore[36] <= 10'd0;
		PixelsStore[37] <= 10'd0;
		PixelsStore[38] <= 10'd0;
		PixelsStore[39] <= 10'd0;
		PixelsStore[40] <= 10'd0;
		PixelsStore[41] <= 10'd0;
		PixelsStore[42] <= 10'd0;
		PixelsStore[43] <= 10'd0;
		PixelsStore[44] <= 10'd0;
		PixelsStore[45] <= 10'd0;
		PixelsStore[46] <= 10'd0;
		PixelsStore[47] <= 10'd0;
		PixelsStore[48] <= 10'd0;
		PixelsStore[49] <= 10'd0;
		PixelsStore[50] <= 10'd0;
		PixelsStore[51] <= 10'd0;
		PixelsStore[52] <= 10'd0;
		PixelsStore[53] <= 10'd0;
		PixelsStore[54] <= 10'd0;
		PixelsStore[55] <= 10'd0;
		PixelsStore[56] <= 10'd0;
		PixelsStore[57] <= 10'd0;
		PixelsStore[58] <= 10'd0;
		PixelsStore[59] <= 10'd0;
		PixelsStore[60] <= 10'd0;
		PixelsStore[61] <= 10'd0;
		PixelsStore[62] <= 10'd0;
		PixelsStore[63] <= 10'd0;
		PixelsStore[64] <= 10'd0;
		PixelsStore[65] <= 10'd0;
		PixelsStore[66] <= 10'd0;
		PixelsStore[67] <= 10'd0;
		PixelsStore[68] <= 10'd0;
		PixelsStore[69] <= 10'd0;
		PixelsStore[70] <= 10'd0;
		PixelsStore[71] <= 10'd0;
		PixelsStore[72] <= 10'd0;
		PixelsStore[73] <= 10'd0;
		PixelsStore[74] <= 10'd0;
		PixelsStore[75] <= 10'd0;
		PixelsStore[76] <= 10'd0;
		PixelsStore[77] <= 10'd0;
		PixelsStore[78] <= 10'd0;
		PixelsStore[79] <= 10'd0;
		PixelsStore[80] <= 10'd0;
		PixelsStore[81] <= 10'd0;
		PixelsStore[82] <= 10'd0;
		PixelsStore[83] <= 10'd0;
		PixelsStore[84] <= 10'd0;
		PixelsStore[85] <= 10'd0;
		PixelsStore[86] <= 10'd0;
		PixelsStore[87] <= 10'd0;
		PixelsStore[88] <= 10'd0;
		PixelsStore[89] <= 10'd0;
		PixelsStore[90] <= 10'd0;
		PixelsStore[91] <= 10'd0;
		PixelsStore[92] <= 10'd0;
		PixelsStore[93] <= 10'd0;
		PixelsStore[94] <= 10'd0;
		PixelsStore[95] <= 10'd0;
		PixelsStore[96] <= 10'd0;
		PixelsStore[97] <= 10'd0;
		PixelsStore[98] <= 10'd0;
		PixelsStore[99] <= 10'd0;
		PixelsStore[100] <= 10'd0;
		PixelsStore[101] <= 10'd0;
		PixelsStore[102] <= 10'd0;
		PixelsStore[103] <= 10'd0;
		PixelsStore[104] <= 10'd0;
		PixelsStore[105] <= 10'd0;
		PixelsStore[106] <= 10'd0;
		PixelsStore[107] <= 10'd0;
		PixelsStore[108] <= 10'd0;
		PixelsStore[109] <= 10'd0;
		PixelsStore[110] <= 10'd0;
		PixelsStore[111] <= 10'd0;
		PixelsStore[112] <= 10'd0;
		PixelsStore[113] <= 10'd0;
		PixelsStore[114] <= 10'd0;
		PixelsStore[115] <= 10'd0;
		PixelsStore[116] <= 10'd0;
		PixelsStore[117] <= 10'd0;
		PixelsStore[118] <= 10'd0;
		PixelsStore[119] <= 10'd0;
		PixelsStore[120] <= 10'd0;
		PixelsStore[121] <= 10'd0;
		PixelsStore[122] <= 10'd0;
		PixelsStore[123] <= 10'd0;
		PixelsStore[124] <= 10'd0;
		PixelsStore[125] <= 10'd0;
		PixelsStore[126] <= 10'd0;
		PixelsStore[127] <= 10'd0;
		PixelsStore[128] <= 10'd0;
		PixelsStore[129] <= 10'd0;
		PixelsStore[130] <= 10'd0;
		PixelsStore[131] <= 10'd0;
		PixelsStore[132] <= 10'd0;
		PixelsStore[133] <= 10'd0;
		PixelsStore[134] <= 10'd0;
		PixelsStore[135] <= 10'd0;
		PixelsStore[136] <= 10'd0;
		PixelsStore[137] <= 10'd0;
		PixelsStore[138] <= 10'd0;
		PixelsStore[139] <= 10'd0;
		PixelsStore[140] <= 10'd0;
		PixelsStore[141] <= 10'd0;
		PixelsStore[142] <= 10'd0;
		PixelsStore[143] <= 10'd0;
		PixelsStore[144] <= 10'd0;
		PixelsStore[145] <= 10'd0;
		PixelsStore[146] <= 10'd0;
		PixelsStore[147] <= 10'd0;
		PixelsStore[148] <= 10'd0;
		PixelsStore[149] <= 10'd0;
		PixelsStore[150] <= 10'd0;
		PixelsStore[151] <= 10'd0;
		PixelsStore[152] <= 10'd0;
		PixelsStore[153] <= 10'd0;
		PixelsStore[154] <= 10'd0;
		PixelsStore[155] <= 10'd0;
		PixelsStore[156] <= 10'd0;
		PixelsStore[157] <= 10'd0;
		PixelsStore[158] <= 10'd0;
		PixelsStore[159] <= 10'd0;
		PixelsStore[160] <= 10'd0;
		PixelsStore[161] <= 10'd0;
		PixelsStore[162] <= 10'd0;
		PixelsStore[163] <= 10'd0;
		PixelsStore[164] <= 10'd0;
		PixelsStore[165] <= 10'd0;
		PixelsStore[166] <= 10'd0;
		PixelsStore[167] <= 10'd0;
		PixelsStore[168] <= 10'd0;
		PixelsStore[169] <= 10'd0;
		PixelsStore[170] <= 10'd0;
		PixelsStore[171] <= 10'd0;
		PixelsStore[172] <= 10'd0;
		PixelsStore[173] <= 10'd0;
		PixelsStore[174] <= 10'd0;
		PixelsStore[175] <= 10'd0;
		PixelsStore[176] <= 10'd0;
		PixelsStore[177] <= 10'd0;
		PixelsStore[178] <= 10'd0;
		PixelsStore[179] <= 10'd0;
		PixelsStore[180] <= 10'd0;
		PixelsStore[181] <= 10'd0;
		PixelsStore[182] <= 10'd0;
		PixelsStore[183] <= 10'd0;
		PixelsStore[184] <= 10'd0;
		PixelsStore[185] <= 10'd0;
		PixelsStore[186] <= 10'd0;
		PixelsStore[187] <= 10'd0;
		PixelsStore[188] <= 10'd0;
		PixelsStore[189] <= 10'd0;
		PixelsStore[190] <= 10'd0;
		PixelsStore[191] <= 10'd0;
		PixelsStore[192] <= 10'd0;
		PixelsStore[193] <= 10'd0;
		PixelsStore[194] <= 10'd0;
		PixelsStore[195] <= 10'd0;
		PixelsStore[196] <= 10'd0;
		PixelsStore[197] <= 10'd0;
		PixelsStore[198] <= 10'd0;
		PixelsStore[199] <= 10'd0;
		PixelsStore[200] <= 10'd0;
		PixelsStore[201] <= 10'd0;
		PixelsStore[202] <= 10'd0;
		PixelsStore[203] <= 10'd0;
		PixelsStore[204] <= 10'd0;
		PixelsStore[205] <= 10'd0;
		PixelsStore[206] <= 10'd0;
		PixelsStore[207] <= 10'd0;
		PixelsStore[208] <= 10'd0;
		PixelsStore[209] <= 10'd0;
		PixelsStore[210] <= 10'd0;
		PixelsStore[211] <= 10'd0;
		PixelsStore[212] <= 10'd0;
		PixelsStore[213] <= 10'd0;
		PixelsStore[214] <= 10'd0;
		PixelsStore[215] <= 10'd0;
		PixelsStore[216] <= 10'd0;
		PixelsStore[217] <= 10'd0;
		PixelsStore[218] <= 10'd0;
		PixelsStore[219] <= 10'd0;
		PixelsStore[220] <= 10'd0;
		PixelsStore[221] <= 10'd0;
		PixelsStore[222] <= 10'd0;
		PixelsStore[223] <= 10'd0;
		PixelsStore[224] <= 10'd0;
		PixelsStore[225] <= 10'd0;
		PixelsStore[226] <= 10'd0;
		PixelsStore[227] <= 10'd0;
		PixelsStore[228] <= 10'd0;
		PixelsStore[229] <= 10'd0;
		PixelsStore[230] <= 10'd0;
		PixelsStore[231] <= 10'd0;
		PixelsStore[232] <= 10'd0;
		PixelsStore[233] <= 10'd0;
		PixelsStore[234] <= 10'd0;
		PixelsStore[235] <= 10'd0;
		PixelsStore[236] <= 10'd0;
		PixelsStore[237] <= 10'd0;
		PixelsStore[238] <= 10'd0;
		PixelsStore[239] <= 10'd0;
		PixelsStore[240] <= 10'd0;
		PixelsStore[241] <= 10'd0;
		PixelsStore[242] <= 10'd0;
		PixelsStore[243] <= 10'd0;
		PixelsStore[244] <= 10'd0;
		PixelsStore[245] <= 10'd0;
		PixelsStore[246] <= 10'd0;
		PixelsStore[247] <= 10'd0;
		PixelsStore[248] <= 10'd0;
		PixelsStore[249] <= 10'd0;
		PixelsStore[250] <= 10'd0;
		PixelsStore[251] <= 10'd0;
		PixelsStore[252] <= 10'd0;
		PixelsStore[253] <= 10'd0;
		PixelsStore[254] <= 10'd0;
		PixelsStore[255] <= 10'd0;
		PixelsStore[256] <= 10'd0;
		PixelsStore[257] <= 10'd0;
		PixelsStore[258] <= 10'd0;
		PixelsStore[259] <= 10'd0;
		PixelsStore[260] <= 10'd0;
		PixelsStore[261] <= 10'd0;
		PixelsStore[262] <= 10'd0;
		PixelsStore[263] <= 10'd0;
		PixelsStore[264] <= 10'd0;
		PixelsStore[265] <= 10'd0;
		PixelsStore[266] <= 10'd0;
		PixelsStore[267] <= 10'd0;
		PixelsStore[268] <= 10'd0;
		PixelsStore[269] <= 10'd0;
		PixelsStore[270] <= 10'd0;
		PixelsStore[271] <= 10'd0;
		PixelsStore[272] <= 10'd0;
		PixelsStore[273] <= 10'd0;
		PixelsStore[274] <= 10'd0;
		PixelsStore[275] <= 10'd0;
		PixelsStore[276] <= 10'd0;
		PixelsStore[277] <= 10'd0;
		PixelsStore[278] <= 10'd0;
		PixelsStore[279] <= 10'd0;
		PixelsStore[280] <= 10'd0;
		PixelsStore[281] <= 10'd0;
		PixelsStore[282] <= 10'd0;
		PixelsStore[283] <= 10'd0;
		PixelsStore[284] <= 10'd0;
		PixelsStore[285] <= 10'd0;
		PixelsStore[286] <= 10'd0;
		PixelsStore[287] <= 10'd0;
		PixelsStore[288] <= 10'd0;
		PixelsStore[289] <= 10'd0;
		PixelsStore[290] <= 10'd0;
		PixelsStore[291] <= 10'd0;
		PixelsStore[292] <= 10'd0;
		PixelsStore[293] <= 10'd0;
		PixelsStore[294] <= 10'd0;
		PixelsStore[295] <= 10'd0;
		PixelsStore[296] <= 10'd0;
		PixelsStore[297] <= 10'd0;
		PixelsStore[298] <= 10'd0;
		PixelsStore[299] <= 10'd0;
		PixelsStore[300] <= 10'd0;
		PixelsStore[301] <= 10'd0;
		PixelsStore[302] <= 10'd0;
		PixelsStore[303] <= 10'd0;
		PixelsStore[304] <= 10'd0;
		PixelsStore[305] <= 10'd0;
		PixelsStore[306] <= 10'd0;
		PixelsStore[307] <= 10'd0;
		PixelsStore[308] <= 10'd0;
		PixelsStore[309] <= 10'd0;
		PixelsStore[310] <= 10'd0;
		PixelsStore[311] <= 10'd0;
		PixelsStore[312] <= 10'd0;
		PixelsStore[313] <= 10'd0;
		PixelsStore[314] <= 10'd0;
		PixelsStore[315] <= 10'd0;
		PixelsStore[316] <= 10'd0;
		PixelsStore[317] <= 10'd0;
		PixelsStore[318] <= 10'd0;
		PixelsStore[319] <= 10'd0;
		PixelsStore[320] <= 10'd0;
		PixelsStore[321] <= 10'd0;
		PixelsStore[322] <= 10'd0;
		PixelsStore[323] <= 10'd0;
		PixelsStore[324] <= 10'd0;
		PixelsStore[325] <= 10'd0;
		PixelsStore[326] <= 10'd0;
		PixelsStore[327] <= 10'd0;
		PixelsStore[328] <= 10'd0;
		PixelsStore[329] <= 10'd0;
		PixelsStore[330] <= 10'd0;
		PixelsStore[331] <= 10'd0;
		PixelsStore[332] <= 10'd0;
		PixelsStore[333] <= 10'd0;
		PixelsStore[334] <= 10'd0;
		PixelsStore[335] <= 10'd0;
		PixelsStore[336] <= 10'd0;
		PixelsStore[337] <= 10'd0;
		PixelsStore[338] <= 10'd0;
		PixelsStore[339] <= 10'd0;
		PixelsStore[340] <= 10'd0;
		PixelsStore[341] <= 10'd0;
		PixelsStore[342] <= 10'd0;
		PixelsStore[343] <= 10'd0;
		PixelsStore[344] <= 10'd0;
		PixelsStore[345] <= 10'd0;
		PixelsStore[346] <= 10'd0;
		PixelsStore[347] <= 10'd0;
		PixelsStore[348] <= 10'd0;
		PixelsStore[349] <= 10'd0;
		PixelsStore[350] <= 10'd0;
		PixelsStore[351] <= 10'd0;
		PixelsStore[352] <= 10'd0;
		PixelsStore[353] <= 10'd0;
		PixelsStore[354] <= 10'd0;
		PixelsStore[355] <= 10'd0;
		PixelsStore[356] <= 10'd0;
		PixelsStore[357] <= 10'd0;
		PixelsStore[358] <= 10'd0;
		PixelsStore[359] <= 10'd0;
		PixelsStore[360] <= 10'd0;
		PixelsStore[361] <= 10'd0;
		PixelsStore[362] <= 10'd0;
		PixelsStore[363] <= 10'd0;
		PixelsStore[364] <= 10'd0;
		PixelsStore[365] <= 10'd0;
		PixelsStore[366] <= 10'd0;
		PixelsStore[367] <= 10'd0;
		PixelsStore[368] <= 10'd0;
		PixelsStore[369] <= 10'd0;
		PixelsStore[370] <= 10'd0;
		PixelsStore[371] <= 10'd0;
		PixelsStore[372] <= 10'd0;
		PixelsStore[373] <= 10'd0;
		PixelsStore[374] <= 10'd0;
		PixelsStore[375] <= 10'd0;
		PixelsStore[376] <= 10'd0;
		PixelsStore[377] <= 10'd0;
		PixelsStore[378] <= 10'd0;
		PixelsStore[379] <= 10'd0;
		PixelsStore[380] <= 10'd0;
		PixelsStore[381] <= 10'd0;
		PixelsStore[382] <= 10'd0;
		PixelsStore[383] <= 10'd0;
		PixelsStore[384] <= 10'd0;
		PixelsStore[385] <= 10'd0;
		PixelsStore[386] <= 10'd0;
		PixelsStore[387] <= 10'd0;
		PixelsStore[388] <= 10'd0;
		PixelsStore[389] <= 10'd0;
		PixelsStore[390] <= 10'd0;
		PixelsStore[391] <= 10'd0;
		PixelsStore[392] <= 10'd0;
		PixelsStore[393] <= 10'd0;
		PixelsStore[394] <= 10'd0;
		PixelsStore[395] <= 10'd0;
		PixelsStore[396] <= 10'd0;
		PixelsStore[397] <= 10'd0;
		PixelsStore[398] <= 10'd0;
		PixelsStore[399] <= 10'd0;
		PixelsStore[400] <= 10'd0;
		PixelsStore[401] <= 10'd0;
		PixelsStore[402] <= 10'd0;
		PixelsStore[403] <= 10'd0;
		PixelsStore[404] <= 10'd0;
		PixelsStore[405] <= 10'd0;
		PixelsStore[406] <= 10'd0;
		PixelsStore[407] <= 10'd0;
		PixelsStore[408] <= 10'd0;
		PixelsStore[409] <= 10'd0;
		PixelsStore[410] <= 10'd0;
		PixelsStore[411] <= 10'd0;
		PixelsStore[412] <= 10'd0;
		PixelsStore[413] <= 10'd0;
		PixelsStore[414] <= 10'd0;
		PixelsStore[415] <= 10'd0;
		PixelsStore[416] <= 10'd0;
		PixelsStore[417] <= 10'd0;
		PixelsStore[418] <= 10'd0;
		PixelsStore[419] <= 10'd0;
		PixelsStore[420] <= 10'd0;
		PixelsStore[421] <= 10'd0;
		PixelsStore[422] <= 10'd0;
		PixelsStore[423] <= 10'd0;
		PixelsStore[424] <= 10'd0;
		PixelsStore[425] <= 10'd0;
		PixelsStore[426] <= 10'd0;
		PixelsStore[427] <= 10'd0;
		PixelsStore[428] <= 10'd0;
		PixelsStore[429] <= 10'd0;
		PixelsStore[430] <= 10'd0;
		PixelsStore[431] <= 10'd0;
		PixelsStore[432] <= 10'd0;
		PixelsStore[433] <= 10'd0;
		PixelsStore[434] <= 10'd0;
		PixelsStore[435] <= 10'd0;
		PixelsStore[436] <= 10'd0;
		PixelsStore[437] <= 10'd0;
		PixelsStore[438] <= 10'd0;
		PixelsStore[439] <= 10'd0;
		PixelsStore[440] <= 10'd0;
		PixelsStore[441] <= 10'd0;
		PixelsStore[442] <= 10'd0;
		PixelsStore[443] <= 10'd0;
		PixelsStore[444] <= 10'd0;
		PixelsStore[445] <= 10'd0;
		PixelsStore[446] <= 10'd0;
		PixelsStore[447] <= 10'd0;
		PixelsStore[448] <= 10'd0;
		PixelsStore[449] <= 10'd0;
		PixelsStore[450] <= 10'd0;
		PixelsStore[451] <= 10'd0;
		PixelsStore[452] <= 10'd0;
		PixelsStore[453] <= 10'd0;
		PixelsStore[454] <= 10'd0;
		PixelsStore[455] <= 10'd0;
		PixelsStore[456] <= 10'd0;
		PixelsStore[457] <= 10'd0;
		PixelsStore[458] <= 10'd0;
		PixelsStore[459] <= 10'd0;
		PixelsStore[460] <= 10'd0;
		PixelsStore[461] <= 10'd0;
		PixelsStore[462] <= 10'd0;
		PixelsStore[463] <= 10'd0;
		PixelsStore[464] <= 10'd0;
		PixelsStore[465] <= 10'd0;
		PixelsStore[466] <= 10'd0;
		PixelsStore[467] <= 10'd0;
		PixelsStore[468] <= 10'd0;
		PixelsStore[469] <= 10'd0;
		PixelsStore[470] <= 10'd0;
		PixelsStore[471] <= 10'd0;
		PixelsStore[472] <= 10'd0;
		PixelsStore[473] <= 10'd0;
		PixelsStore[474] <= 10'd0;
		PixelsStore[475] <= 10'd0;
		PixelsStore[476] <= 10'd0;
		PixelsStore[477] <= 10'd0;
		PixelsStore[478] <= 10'd0;
		PixelsStore[479] <= 10'd0;
		PixelsStore[480] <= 10'd0;
		PixelsStore[481] <= 10'd0;
		PixelsStore[482] <= 10'd0;
		PixelsStore[483] <= 10'd0;
		PixelsStore[484] <= 10'd0;
		PixelsStore[485] <= 10'd0;
		PixelsStore[486] <= 10'd0;
		PixelsStore[487] <= 10'd0;
		PixelsStore[488] <= 10'd0;
		PixelsStore[489] <= 10'd0;
		PixelsStore[490] <= 10'd0;
		PixelsStore[491] <= 10'd0;
		PixelsStore[492] <= 10'd0;
		PixelsStore[493] <= 10'd0;
		PixelsStore[494] <= 10'd0;
		PixelsStore[495] <= 10'd0;
		PixelsStore[496] <= 10'd0;
		PixelsStore[497] <= 10'd0;
		PixelsStore[498] <= 10'd0;
		PixelsStore[499] <= 10'd0;
		PixelsStore[500] <= 10'd0;
		PixelsStore[501] <= 10'd0;
		PixelsStore[502] <= 10'd0;
		PixelsStore[503] <= 10'd0;
		PixelsStore[504] <= 10'd0;
		PixelsStore[505] <= 10'd0;
		PixelsStore[506] <= 10'd0;
		PixelsStore[507] <= 10'd0;
		PixelsStore[508] <= 10'd0;
		PixelsStore[509] <= 10'd0;
		PixelsStore[510] <= 10'd0;
		PixelsStore[511] <= 10'd0;
		PixelsStore[512] <= 10'd0;
		PixelsStore[513] <= 10'd0;
		PixelsStore[514] <= 10'd0;
		PixelsStore[515] <= 10'd0;
		PixelsStore[516] <= 10'd0;
		PixelsStore[517] <= 10'd0;
		PixelsStore[518] <= 10'd0;
		PixelsStore[519] <= 10'd0;
		PixelsStore[520] <= 10'd0;
		PixelsStore[521] <= 10'd0;
		PixelsStore[522] <= 10'd0;
		PixelsStore[523] <= 10'd0;
		PixelsStore[524] <= 10'd0;
		PixelsStore[525] <= 10'd0;
		PixelsStore[526] <= 10'd0;
		PixelsStore[527] <= 10'd0;
		PixelsStore[528] <= 10'd0;
		PixelsStore[529] <= 10'd0;
		PixelsStore[530] <= 10'd0;
		PixelsStore[531] <= 10'd0;
		PixelsStore[532] <= 10'd0;
		PixelsStore[533] <= 10'd0;
		PixelsStore[534] <= 10'd0;
		PixelsStore[535] <= 10'd0;
		PixelsStore[536] <= 10'd0;
		PixelsStore[537] <= 10'd0;
		PixelsStore[538] <= 10'd0;
		PixelsStore[539] <= 10'd0;
		PixelsStore[540] <= 10'd0;
		PixelsStore[541] <= 10'd0;
		PixelsStore[542] <= 10'd0;
		PixelsStore[543] <= 10'd0;
		PixelsStore[544] <= 10'd0;
		PixelsStore[545] <= 10'd0;
		PixelsStore[546] <= 10'd0;
		PixelsStore[547] <= 10'd0;
		PixelsStore[548] <= 10'd0;
		PixelsStore[549] <= 10'd0;
		PixelsStore[550] <= 10'd0;
		PixelsStore[551] <= 10'd0;
		PixelsStore[552] <= 10'd0;
		PixelsStore[553] <= 10'd0;
		PixelsStore[554] <= 10'd0;
		PixelsStore[555] <= 10'd0;
		PixelsStore[556] <= 10'd0;
		PixelsStore[557] <= 10'd0;
		PixelsStore[558] <= 10'd0;
		PixelsStore[559] <= 10'd0;
		PixelsStore[560] <= 10'd0;
		PixelsStore[561] <= 10'd0;
		PixelsStore[562] <= 10'd0;
		PixelsStore[563] <= 10'd0;
		PixelsStore[564] <= 10'd0;
		PixelsStore[565] <= 10'd0;
		PixelsStore[566] <= 10'd0;
		PixelsStore[567] <= 10'd0;
		PixelsStore[568] <= 10'd0;
		PixelsStore[569] <= 10'd0;
		PixelsStore[570] <= 10'd0;
		PixelsStore[571] <= 10'd0;
		PixelsStore[572] <= 10'd0;
		PixelsStore[573] <= 10'd0;
		PixelsStore[574] <= 10'd0;
		PixelsStore[575] <= 10'd0;
		PixelsStore[576] <= 10'd0;
		PixelsStore[577] <= 10'd0;
		PixelsStore[578] <= 10'd0;
		PixelsStore[579] <= 10'd0;
		PixelsStore[580] <= 10'd0;
		PixelsStore[581] <= 10'd0;
		PixelsStore[582] <= 10'd0;
		PixelsStore[583] <= 10'd0;
		PixelsStore[584] <= 10'd0;
		PixelsStore[585] <= 10'd0;
		PixelsStore[586] <= 10'd0;
		PixelsStore[587] <= 10'd0;
		PixelsStore[588] <= 10'd0;
		PixelsStore[589] <= 10'd0;
		PixelsStore[590] <= 10'd0;
		PixelsStore[591] <= 10'd0;
		PixelsStore[592] <= 10'd0;
		PixelsStore[593] <= 10'd0;
		PixelsStore[594] <= 10'd0;
		PixelsStore[595] <= 10'd0;
		PixelsStore[596] <= 10'd0;
		PixelsStore[597] <= 10'd0;
		PixelsStore[598] <= 10'd0;
		PixelsStore[599] <= 10'd0;
		PixelsStore[600] <= 10'd0;
		PixelsStore[601] <= 10'd0;
		PixelsStore[602] <= 10'd0;
		PixelsStore[603] <= 10'd0;
		PixelsStore[604] <= 10'd0;
		PixelsStore[605] <= 10'd0;
		PixelsStore[606] <= 10'd0;
		PixelsStore[607] <= 10'd0;
		PixelsStore[608] <= 10'd0;
		PixelsStore[609] <= 10'd0;
		PixelsStore[610] <= 10'd0;
		PixelsStore[611] <= 10'd0;
		PixelsStore[612] <= 10'd0;
		PixelsStore[613] <= 10'd0;
		PixelsStore[614] <= 10'd0;
		PixelsStore[615] <= 10'd0;
		PixelsStore[616] <= 10'd0;
		PixelsStore[617] <= 10'd0;
		PixelsStore[618] <= 10'd0;
		PixelsStore[619] <= 10'd0;
		PixelsStore[620] <= 10'd0;
		PixelsStore[621] <= 10'd0;
		PixelsStore[622] <= 10'd0;
		PixelsStore[623] <= 10'd0;
		PixelsStore[624] <= 10'd0;
		PixelsStore[625] <= 10'd0;
		PixelsStore[626] <= 10'd0;
		PixelsStore[627] <= 10'd0;
		PixelsStore[628] <= 10'd0;
		PixelsStore[629] <= 10'd0;
		PixelsStore[630] <= 10'd0;
		PixelsStore[631] <= 10'd0;
		PixelsStore[632] <= 10'd0;
		PixelsStore[633] <= 10'd0;
		PixelsStore[634] <= 10'd0;
		PixelsStore[635] <= 10'd0;
		PixelsStore[636] <= 10'd0;
		PixelsStore[637] <= 10'd0;
		PixelsStore[638] <= 10'd0;
		PixelsStore[639] <= 10'd0;
		PixelsStore[640] <= 10'd0;
		PixelsStore[641] <= 10'd0;
		PixelsStore[642] <= 10'd0;
		PixelsStore[643] <= 10'd0;
		PixelsStore[644] <= 10'd0;
		PixelsStore[645] <= 10'd0;
		PixelsStore[646] <= 10'd0;
		PixelsStore[647] <= 10'd0;
		PixelsStore[648] <= 10'd0;
		PixelsStore[649] <= 10'd0;
		PixelsStore[650] <= 10'd0;
		PixelsStore[651] <= 10'd0;
		PixelsStore[652] <= 10'd0;
		PixelsStore[653] <= 10'd0;
		PixelsStore[654] <= 10'd0;
		PixelsStore[655] <= 10'd0;
		PixelsStore[656] <= 10'd0;
		PixelsStore[657] <= 10'd0;
		PixelsStore[658] <= 10'd0;
		PixelsStore[659] <= 10'd0;
		PixelsStore[660] <= 10'd0;
		PixelsStore[661] <= 10'd0;
		PixelsStore[662] <= 10'd0;
		PixelsStore[663] <= 10'd0;
		PixelsStore[664] <= 10'd0;
		PixelsStore[665] <= 10'd0;
		PixelsStore[666] <= 10'd0;
		PixelsStore[667] <= 10'd0;
		PixelsStore[668] <= 10'd0;
		PixelsStore[669] <= 10'd0;
		PixelsStore[670] <= 10'd0;
		PixelsStore[671] <= 10'd0;
		PixelsStore[672] <= 10'd0;
		PixelsStore[673] <= 10'd0;
		PixelsStore[674] <= 10'd0;
		PixelsStore[675] <= 10'd0;
		PixelsStore[676] <= 10'd0;
		PixelsStore[677] <= 10'd0;
		PixelsStore[678] <= 10'd0;
		PixelsStore[679] <= 10'd0;
		PixelsStore[680] <= 10'd0;
		PixelsStore[681] <= 10'd0;
		PixelsStore[682] <= 10'd0;
		PixelsStore[683] <= 10'd0;
		PixelsStore[684] <= 10'd0;
		PixelsStore[685] <= 10'd0;
		PixelsStore[686] <= 10'd0;
		PixelsStore[687] <= 10'd0;
		PixelsStore[688] <= 10'd0;
		PixelsStore[689] <= 10'd0;
		PixelsStore[690] <= 10'd0;
		PixelsStore[691] <= 10'd0;
		PixelsStore[692] <= 10'd0;
		PixelsStore[693] <= 10'd0;
		PixelsStore[694] <= 10'd0;
		PixelsStore[695] <= 10'd0;
		PixelsStore[696] <= 10'd0;
		PixelsStore[697] <= 10'd0;
		PixelsStore[698] <= 10'd0;
		PixelsStore[699] <= 10'd0;
		PixelsStore[700] <= 10'd0;
		PixelsStore[701] <= 10'd0;
		PixelsStore[702] <= 10'd0;
		PixelsStore[703] <= 10'd0;
		PixelsStore[704] <= 10'd0;
		PixelsStore[705] <= 10'd0;
		PixelsStore[706] <= 10'd0;
		PixelsStore[707] <= 10'd0;
		PixelsStore[708] <= 10'd0;
		PixelsStore[709] <= 10'd0;
		PixelsStore[710] <= 10'd0;
		PixelsStore[711] <= 10'd0;
		PixelsStore[712] <= 10'd0;
		PixelsStore[713] <= 10'd0;
		PixelsStore[714] <= 10'd0;
		PixelsStore[715] <= 10'd0;
		PixelsStore[716] <= 10'd0;
		PixelsStore[717] <= 10'd0;
		PixelsStore[718] <= 10'd0;
		PixelsStore[719] <= 10'd0;
		PixelsStore[720] <= 10'd0;
		PixelsStore[721] <= 10'd0;
		PixelsStore[722] <= 10'd0;
		PixelsStore[723] <= 10'd0;
		PixelsStore[724] <= 10'd0;
		PixelsStore[725] <= 10'd0;
		PixelsStore[726] <= 10'd0;
		PixelsStore[727] <= 10'd0;
		PixelsStore[728] <= 10'd0;
		PixelsStore[729] <= 10'd0;
		PixelsStore[730] <= 10'd0;
		PixelsStore[731] <= 10'd0;
		PixelsStore[732] <= 10'd0;
		PixelsStore[733] <= 10'd0;
		PixelsStore[734] <= 10'd0;
		PixelsStore[735] <= 10'd0;
		PixelsStore[736] <= 10'd0;
		PixelsStore[737] <= 10'd0;
		PixelsStore[738] <= 10'd0;
		PixelsStore[739] <= 10'd0;
		PixelsStore[740] <= 10'd0;
		PixelsStore[741] <= 10'd0;
		PixelsStore[742] <= 10'd0;
		PixelsStore[743] <= 10'd0;
		PixelsStore[744] <= 10'd0;
		PixelsStore[745] <= 10'd0;
		PixelsStore[746] <= 10'd0;
		PixelsStore[747] <= 10'd0;
		PixelsStore[748] <= 10'd0;
		PixelsStore[749] <= 10'd0;
		PixelsStore[750] <= 10'd0;
		PixelsStore[751] <= 10'd0;
		PixelsStore[752] <= 10'd0;
		PixelsStore[753] <= 10'd0;
		PixelsStore[754] <= 10'd0;
		PixelsStore[755] <= 10'd0;
		PixelsStore[756] <= 10'd0;
		PixelsStore[757] <= 10'd0;
		PixelsStore[758] <= 10'd0;
		PixelsStore[759] <= 10'd0;
		PixelsStore[760] <= 10'd0;
		PixelsStore[761] <= 10'd0;
		PixelsStore[762] <= 10'd0;
		PixelsStore[763] <= 10'd0;
		PixelsStore[764] <= 10'd0;
		PixelsStore[765] <= 10'd0;
		PixelsStore[766] <= 10'd0;
		PixelsStore[767] <= 10'd0;
		PixelsStore[768] <= 10'd0;
		PixelsStore[769] <= 10'd0;
		PixelsStore[770] <= 10'd0;
		PixelsStore[771] <= 10'd0;
		PixelsStore[772] <= 10'd0;
		PixelsStore[773] <= 10'd0;
		PixelsStore[774] <= 10'd0;
		PixelsStore[775] <= 10'd0;
		PixelsStore[776] <= 10'd0;
		PixelsStore[777] <= 10'd0;
		PixelsStore[778] <= 10'd0;
		PixelsStore[779] <= 10'd0;
		PixelsStore[780] <= 10'd0;
		PixelsStore[781] <= 10'd0;
		PixelsStore[782] <= 10'd0;
		PixelsStore[783] <= 10'd0;
		PixelsStore[784] <= 10'd0;
		WeightsStore0[0] <= 19'd0;
		WeightsStore0[1] <= 19'd0;
		WeightsStore0[2] <= 19'd0;
		WeightsStore0[3] <= 19'd0;
		WeightsStore0[4] <= 19'd0;
		WeightsStore0[5] <= 19'd0;
		WeightsStore0[6] <= 19'd0;
		WeightsStore0[7] <= 19'd0;
		WeightsStore0[8] <= 19'd0;
		WeightsStore0[9] <= 19'd0;
		WeightsStore0[10] <= 19'd0;
		WeightsStore0[11] <= 19'd0;
		WeightsStore0[12] <= 19'd0;
		WeightsStore0[13] <= 19'd0;
		WeightsStore0[14] <= 19'd0;
		WeightsStore0[15] <= 19'd0;
		WeightsStore0[16] <= 19'd0;
		WeightsStore0[17] <= 19'd0;
		WeightsStore0[18] <= 19'd0;
		WeightsStore0[19] <= 19'd0;
		WeightsStore0[20] <= 19'd0;
		WeightsStore0[21] <= 19'd0;
		WeightsStore0[22] <= 19'd0;
		WeightsStore0[23] <= 19'd0;
		WeightsStore0[24] <= 19'd0;
		WeightsStore0[25] <= 19'd0;
		WeightsStore0[26] <= 19'd0;
		WeightsStore0[27] <= 19'd0;
		WeightsStore0[28] <= 19'd0;
		WeightsStore0[29] <= 19'd0;
		WeightsStore0[30] <= 19'd0;
		WeightsStore0[31] <= 19'd0;
		WeightsStore0[32] <= 19'd0;
		WeightsStore0[33] <= 19'd0;
		WeightsStore0[34] <= 19'd0;
		WeightsStore0[35] <= 19'd0;
		WeightsStore0[36] <= 19'd0;
		WeightsStore0[37] <= 19'd0;
		WeightsStore0[38] <= 19'd0;
		WeightsStore0[39] <= 19'd0;
		WeightsStore0[40] <= 19'd0;
		WeightsStore0[41] <= 19'd0;
		WeightsStore0[42] <= 19'd0;
		WeightsStore0[43] <= 19'd0;
		WeightsStore0[44] <= 19'd0;
		WeightsStore0[45] <= 19'd0;
		WeightsStore0[46] <= 19'd0;
		WeightsStore0[47] <= 19'd0;
		WeightsStore0[48] <= 19'd0;
		WeightsStore0[49] <= 19'd0;
		WeightsStore0[50] <= 19'd0;
		WeightsStore0[51] <= 19'd0;
		WeightsStore0[52] <= 19'd0;
		WeightsStore0[53] <= 19'd0;
		WeightsStore0[54] <= 19'd0;
		WeightsStore0[55] <= 19'd0;
		WeightsStore0[56] <= 19'd0;
		WeightsStore0[57] <= 19'd0;
		WeightsStore0[58] <= 19'd0;
		WeightsStore0[59] <= 19'd0;
		WeightsStore0[60] <= 19'd0;
		WeightsStore0[61] <= 19'd0;
		WeightsStore0[62] <= 19'd0;
		WeightsStore0[63] <= 19'd0;
		WeightsStore0[64] <= 19'd0;
		WeightsStore0[65] <= 19'd0;
		WeightsStore0[66] <= 19'd0;
		WeightsStore0[67] <= 19'd0;
		WeightsStore0[68] <= 19'd0;
		WeightsStore0[69] <= 19'd0;
		WeightsStore0[70] <= 19'd0;
		WeightsStore0[71] <= 19'd0;
		WeightsStore0[72] <= 19'd0;
		WeightsStore0[73] <= 19'd0;
		WeightsStore0[74] <= 19'd0;
		WeightsStore0[75] <= 19'd0;
		WeightsStore0[76] <= 19'd0;
		WeightsStore0[77] <= 19'd0;
		WeightsStore0[78] <= 19'd0;
		WeightsStore0[79] <= 19'd0;
		WeightsStore0[80] <= 19'd0;
		WeightsStore0[81] <= 19'd0;
		WeightsStore0[82] <= 19'd0;
		WeightsStore0[83] <= 19'd0;
		WeightsStore0[84] <= 19'd0;
		WeightsStore0[85] <= 19'd0;
		WeightsStore0[86] <= 19'd0;
		WeightsStore0[87] <= 19'd0;
		WeightsStore0[88] <= 19'd0;
		WeightsStore0[89] <= 19'd0;
		WeightsStore0[90] <= 19'd0;
		WeightsStore0[91] <= 19'd0;
		WeightsStore0[92] <= 19'd0;
		WeightsStore0[93] <= 19'd0;
		WeightsStore0[94] <= 19'd0;
		WeightsStore0[95] <= 19'd0;
		WeightsStore0[96] <= 19'd0;
		WeightsStore0[97] <= 19'd0;
		WeightsStore0[98] <= 19'd0;
		WeightsStore0[99] <= 19'd0;
		WeightsStore0[100] <= 19'd0;
		WeightsStore0[101] <= 19'd0;
		WeightsStore0[102] <= 19'd0;
		WeightsStore0[103] <= 19'd0;
		WeightsStore0[104] <= 19'd0;
		WeightsStore0[105] <= 19'd0;
		WeightsStore0[106] <= 19'd0;
		WeightsStore0[107] <= 19'd0;
		WeightsStore0[108] <= 19'd0;
		WeightsStore0[109] <= 19'd0;
		WeightsStore0[110] <= 19'd0;
		WeightsStore0[111] <= 19'd0;
		WeightsStore0[112] <= 19'd0;
		WeightsStore0[113] <= 19'd0;
		WeightsStore0[114] <= 19'd0;
		WeightsStore0[115] <= 19'd0;
		WeightsStore0[116] <= 19'd0;
		WeightsStore0[117] <= 19'd0;
		WeightsStore0[118] <= 19'd0;
		WeightsStore0[119] <= 19'd0;
		WeightsStore0[120] <= 19'd0;
		WeightsStore0[121] <= 19'd0;
		WeightsStore0[122] <= 19'd0;
		WeightsStore0[123] <= 19'd0;
		WeightsStore0[124] <= 19'd0;
		WeightsStore0[125] <= 19'd0;
		WeightsStore0[126] <= 19'd0;
		WeightsStore0[127] <= 19'd0;
		WeightsStore0[128] <= 19'd0;
		WeightsStore0[129] <= 19'd0;
		WeightsStore0[130] <= 19'd0;
		WeightsStore0[131] <= 19'd0;
		WeightsStore0[132] <= 19'd0;
		WeightsStore0[133] <= 19'd0;
		WeightsStore0[134] <= 19'd0;
		WeightsStore0[135] <= 19'd0;
		WeightsStore0[136] <= 19'd0;
		WeightsStore0[137] <= 19'd0;
		WeightsStore0[138] <= 19'd0;
		WeightsStore0[139] <= 19'd0;
		WeightsStore0[140] <= 19'd0;
		WeightsStore0[141] <= 19'd0;
		WeightsStore0[142] <= 19'd0;
		WeightsStore0[143] <= 19'd0;
		WeightsStore0[144] <= 19'd0;
		WeightsStore0[145] <= 19'd0;
		WeightsStore0[146] <= 19'd0;
		WeightsStore0[147] <= 19'd0;
		WeightsStore0[148] <= 19'd0;
		WeightsStore0[149] <= 19'd0;
		WeightsStore0[150] <= 19'd0;
		WeightsStore0[151] <= 19'd0;
		WeightsStore0[152] <= 19'd0;
		WeightsStore0[153] <= 19'd0;
		WeightsStore0[154] <= 19'd0;
		WeightsStore0[155] <= 19'd0;
		WeightsStore0[156] <= 19'd0;
		WeightsStore0[157] <= 19'd0;
		WeightsStore0[158] <= 19'd0;
		WeightsStore0[159] <= 19'd0;
		WeightsStore0[160] <= 19'd0;
		WeightsStore0[161] <= 19'd0;
		WeightsStore0[162] <= 19'd0;
		WeightsStore0[163] <= 19'd0;
		WeightsStore0[164] <= 19'd0;
		WeightsStore0[165] <= 19'd0;
		WeightsStore0[166] <= 19'd0;
		WeightsStore0[167] <= 19'd0;
		WeightsStore0[168] <= 19'd0;
		WeightsStore0[169] <= 19'd0;
		WeightsStore0[170] <= 19'd0;
		WeightsStore0[171] <= 19'd0;
		WeightsStore0[172] <= 19'd0;
		WeightsStore0[173] <= 19'd0;
		WeightsStore0[174] <= 19'd0;
		WeightsStore0[175] <= 19'd0;
		WeightsStore0[176] <= 19'd0;
		WeightsStore0[177] <= 19'd0;
		WeightsStore0[178] <= 19'd0;
		WeightsStore0[179] <= 19'd0;
		WeightsStore0[180] <= 19'd0;
		WeightsStore0[181] <= 19'd0;
		WeightsStore0[182] <= 19'd0;
		WeightsStore0[183] <= 19'd0;
		WeightsStore0[184] <= 19'd0;
		WeightsStore0[185] <= 19'd0;
		WeightsStore0[186] <= 19'd0;
		WeightsStore0[187] <= 19'd0;
		WeightsStore0[188] <= 19'd0;
		WeightsStore0[189] <= 19'd0;
		WeightsStore0[190] <= 19'd0;
		WeightsStore0[191] <= 19'd0;
		WeightsStore0[192] <= 19'd0;
		WeightsStore0[193] <= 19'd0;
		WeightsStore0[194] <= 19'd0;
		WeightsStore0[195] <= 19'd0;
		WeightsStore0[196] <= 19'd0;
		WeightsStore0[197] <= 19'd0;
		WeightsStore0[198] <= 19'd0;
		WeightsStore0[199] <= 19'd0;
		WeightsStore0[200] <= 19'd0;
		WeightsStore0[201] <= 19'd0;
		WeightsStore0[202] <= 19'd0;
		WeightsStore0[203] <= 19'd0;
		WeightsStore0[204] <= 19'd0;
		WeightsStore0[205] <= 19'd0;
		WeightsStore0[206] <= 19'd0;
		WeightsStore0[207] <= 19'd0;
		WeightsStore0[208] <= 19'd0;
		WeightsStore0[209] <= 19'd0;
		WeightsStore0[210] <= 19'd0;
		WeightsStore0[211] <= 19'd0;
		WeightsStore0[212] <= 19'd0;
		WeightsStore0[213] <= 19'd0;
		WeightsStore0[214] <= 19'd0;
		WeightsStore0[215] <= 19'd0;
		WeightsStore0[216] <= 19'd0;
		WeightsStore0[217] <= 19'd0;
		WeightsStore0[218] <= 19'd0;
		WeightsStore0[219] <= 19'd0;
		WeightsStore0[220] <= 19'd0;
		WeightsStore0[221] <= 19'd0;
		WeightsStore0[222] <= 19'd0;
		WeightsStore0[223] <= 19'd0;
		WeightsStore0[224] <= 19'd0;
		WeightsStore0[225] <= 19'd0;
		WeightsStore0[226] <= 19'd0;
		WeightsStore0[227] <= 19'd0;
		WeightsStore0[228] <= 19'd0;
		WeightsStore0[229] <= 19'd0;
		WeightsStore0[230] <= 19'd0;
		WeightsStore0[231] <= 19'd0;
		WeightsStore0[232] <= 19'd0;
		WeightsStore0[233] <= 19'd0;
		WeightsStore0[234] <= 19'd0;
		WeightsStore0[235] <= 19'd0;
		WeightsStore0[236] <= 19'd0;
		WeightsStore0[237] <= 19'd0;
		WeightsStore0[238] <= 19'd0;
		WeightsStore0[239] <= 19'd0;
		WeightsStore0[240] <= 19'd0;
		WeightsStore0[241] <= 19'd0;
		WeightsStore0[242] <= 19'd0;
		WeightsStore0[243] <= 19'd0;
		WeightsStore0[244] <= 19'd0;
		WeightsStore0[245] <= 19'd0;
		WeightsStore0[246] <= 19'd0;
		WeightsStore0[247] <= 19'd0;
		WeightsStore0[248] <= 19'd0;
		WeightsStore0[249] <= 19'd0;
		WeightsStore0[250] <= 19'd0;
		WeightsStore0[251] <= 19'd0;
		WeightsStore0[252] <= 19'd0;
		WeightsStore0[253] <= 19'd0;
		WeightsStore0[254] <= 19'd0;
		WeightsStore0[255] <= 19'd0;
		WeightsStore0[256] <= 19'd0;
		WeightsStore0[257] <= 19'd0;
		WeightsStore0[258] <= 19'd0;
		WeightsStore0[259] <= 19'd0;
		WeightsStore0[260] <= 19'd0;
		WeightsStore0[261] <= 19'd0;
		WeightsStore0[262] <= 19'd0;
		WeightsStore0[263] <= 19'd0;
		WeightsStore0[264] <= 19'd0;
		WeightsStore0[265] <= 19'd0;
		WeightsStore0[266] <= 19'd0;
		WeightsStore0[267] <= 19'd0;
		WeightsStore0[268] <= 19'd0;
		WeightsStore0[269] <= 19'd0;
		WeightsStore0[270] <= 19'd0;
		WeightsStore0[271] <= 19'd0;
		WeightsStore0[272] <= 19'd0;
		WeightsStore0[273] <= 19'd0;
		WeightsStore0[274] <= 19'd0;
		WeightsStore0[275] <= 19'd0;
		WeightsStore0[276] <= 19'd0;
		WeightsStore0[277] <= 19'd0;
		WeightsStore0[278] <= 19'd0;
		WeightsStore0[279] <= 19'd0;
		WeightsStore0[280] <= 19'd0;
		WeightsStore0[281] <= 19'd0;
		WeightsStore0[282] <= 19'd0;
		WeightsStore0[283] <= 19'd0;
		WeightsStore0[284] <= 19'd0;
		WeightsStore0[285] <= 19'd0;
		WeightsStore0[286] <= 19'd0;
		WeightsStore0[287] <= 19'd0;
		WeightsStore0[288] <= 19'd0;
		WeightsStore0[289] <= 19'd0;
		WeightsStore0[290] <= 19'd0;
		WeightsStore0[291] <= 19'd0;
		WeightsStore0[292] <= 19'd0;
		WeightsStore0[293] <= 19'd0;
		WeightsStore0[294] <= 19'd0;
		WeightsStore0[295] <= 19'd0;
		WeightsStore0[296] <= 19'd0;
		WeightsStore0[297] <= 19'd0;
		WeightsStore0[298] <= 19'd0;
		WeightsStore0[299] <= 19'd0;
		WeightsStore0[300] <= 19'd0;
		WeightsStore0[301] <= 19'd0;
		WeightsStore0[302] <= 19'd0;
		WeightsStore0[303] <= 19'd0;
		WeightsStore0[304] <= 19'd0;
		WeightsStore0[305] <= 19'd0;
		WeightsStore0[306] <= 19'd0;
		WeightsStore0[307] <= 19'd0;
		WeightsStore0[308] <= 19'd0;
		WeightsStore0[309] <= 19'd0;
		WeightsStore0[310] <= 19'd0;
		WeightsStore0[311] <= 19'd0;
		WeightsStore0[312] <= 19'd0;
		WeightsStore0[313] <= 19'd0;
		WeightsStore0[314] <= 19'd0;
		WeightsStore0[315] <= 19'd0;
		WeightsStore0[316] <= 19'd0;
		WeightsStore0[317] <= 19'd0;
		WeightsStore0[318] <= 19'd0;
		WeightsStore0[319] <= 19'd0;
		WeightsStore0[320] <= 19'd0;
		WeightsStore0[321] <= 19'd0;
		WeightsStore0[322] <= 19'd0;
		WeightsStore0[323] <= 19'd0;
		WeightsStore0[324] <= 19'd0;
		WeightsStore0[325] <= 19'd0;
		WeightsStore0[326] <= 19'd0;
		WeightsStore0[327] <= 19'd0;
		WeightsStore0[328] <= 19'd0;
		WeightsStore0[329] <= 19'd0;
		WeightsStore0[330] <= 19'd0;
		WeightsStore0[331] <= 19'd0;
		WeightsStore0[332] <= 19'd0;
		WeightsStore0[333] <= 19'd0;
		WeightsStore0[334] <= 19'd0;
		WeightsStore0[335] <= 19'd0;
		WeightsStore0[336] <= 19'd0;
		WeightsStore0[337] <= 19'd0;
		WeightsStore0[338] <= 19'd0;
		WeightsStore0[339] <= 19'd0;
		WeightsStore0[340] <= 19'd0;
		WeightsStore0[341] <= 19'd0;
		WeightsStore0[342] <= 19'd0;
		WeightsStore0[343] <= 19'd0;
		WeightsStore0[344] <= 19'd0;
		WeightsStore0[345] <= 19'd0;
		WeightsStore0[346] <= 19'd0;
		WeightsStore0[347] <= 19'd0;
		WeightsStore0[348] <= 19'd0;
		WeightsStore0[349] <= 19'd0;
		WeightsStore0[350] <= 19'd0;
		WeightsStore0[351] <= 19'd0;
		WeightsStore0[352] <= 19'd0;
		WeightsStore0[353] <= 19'd0;
		WeightsStore0[354] <= 19'd0;
		WeightsStore0[355] <= 19'd0;
		WeightsStore0[356] <= 19'd0;
		WeightsStore0[357] <= 19'd0;
		WeightsStore0[358] <= 19'd0;
		WeightsStore0[359] <= 19'd0;
		WeightsStore0[360] <= 19'd0;
		WeightsStore0[361] <= 19'd0;
		WeightsStore0[362] <= 19'd0;
		WeightsStore0[363] <= 19'd0;
		WeightsStore0[364] <= 19'd0;
		WeightsStore0[365] <= 19'd0;
		WeightsStore0[366] <= 19'd0;
		WeightsStore0[367] <= 19'd0;
		WeightsStore0[368] <= 19'd0;
		WeightsStore0[369] <= 19'd0;
		WeightsStore0[370] <= 19'd0;
		WeightsStore0[371] <= 19'd0;
		WeightsStore0[372] <= 19'd0;
		WeightsStore0[373] <= 19'd0;
		WeightsStore0[374] <= 19'd0;
		WeightsStore0[375] <= 19'd0;
		WeightsStore0[376] <= 19'd0;
		WeightsStore0[377] <= 19'd0;
		WeightsStore0[378] <= 19'd0;
		WeightsStore0[379] <= 19'd0;
		WeightsStore0[380] <= 19'd0;
		WeightsStore0[381] <= 19'd0;
		WeightsStore0[382] <= 19'd0;
		WeightsStore0[383] <= 19'd0;
		WeightsStore0[384] <= 19'd0;
		WeightsStore0[385] <= 19'd0;
		WeightsStore0[386] <= 19'd0;
		WeightsStore0[387] <= 19'd0;
		WeightsStore0[388] <= 19'd0;
		WeightsStore0[389] <= 19'd0;
		WeightsStore0[390] <= 19'd0;
		WeightsStore0[391] <= 19'd0;
		WeightsStore0[392] <= 19'd0;
		WeightsStore0[393] <= 19'd0;
		WeightsStore0[394] <= 19'd0;
		WeightsStore0[395] <= 19'd0;
		WeightsStore0[396] <= 19'd0;
		WeightsStore0[397] <= 19'd0;
		WeightsStore0[398] <= 19'd0;
		WeightsStore0[399] <= 19'd0;
		WeightsStore0[400] <= 19'd0;
		WeightsStore0[401] <= 19'd0;
		WeightsStore0[402] <= 19'd0;
		WeightsStore0[403] <= 19'd0;
		WeightsStore0[404] <= 19'd0;
		WeightsStore0[405] <= 19'd0;
		WeightsStore0[406] <= 19'd0;
		WeightsStore0[407] <= 19'd0;
		WeightsStore0[408] <= 19'd0;
		WeightsStore0[409] <= 19'd0;
		WeightsStore0[410] <= 19'd0;
		WeightsStore0[411] <= 19'd0;
		WeightsStore0[412] <= 19'd0;
		WeightsStore0[413] <= 19'd0;
		WeightsStore0[414] <= 19'd0;
		WeightsStore0[415] <= 19'd0;
		WeightsStore0[416] <= 19'd0;
		WeightsStore0[417] <= 19'd0;
		WeightsStore0[418] <= 19'd0;
		WeightsStore0[419] <= 19'd0;
		WeightsStore0[420] <= 19'd0;
		WeightsStore0[421] <= 19'd0;
		WeightsStore0[422] <= 19'd0;
		WeightsStore0[423] <= 19'd0;
		WeightsStore0[424] <= 19'd0;
		WeightsStore0[425] <= 19'd0;
		WeightsStore0[426] <= 19'd0;
		WeightsStore0[427] <= 19'd0;
		WeightsStore0[428] <= 19'd0;
		WeightsStore0[429] <= 19'd0;
		WeightsStore0[430] <= 19'd0;
		WeightsStore0[431] <= 19'd0;
		WeightsStore0[432] <= 19'd0;
		WeightsStore0[433] <= 19'd0;
		WeightsStore0[434] <= 19'd0;
		WeightsStore0[435] <= 19'd0;
		WeightsStore0[436] <= 19'd0;
		WeightsStore0[437] <= 19'd0;
		WeightsStore0[438] <= 19'd0;
		WeightsStore0[439] <= 19'd0;
		WeightsStore0[440] <= 19'd0;
		WeightsStore0[441] <= 19'd0;
		WeightsStore0[442] <= 19'd0;
		WeightsStore0[443] <= 19'd0;
		WeightsStore0[444] <= 19'd0;
		WeightsStore0[445] <= 19'd0;
		WeightsStore0[446] <= 19'd0;
		WeightsStore0[447] <= 19'd0;
		WeightsStore0[448] <= 19'd0;
		WeightsStore0[449] <= 19'd0;
		WeightsStore0[450] <= 19'd0;
		WeightsStore0[451] <= 19'd0;
		WeightsStore0[452] <= 19'd0;
		WeightsStore0[453] <= 19'd0;
		WeightsStore0[454] <= 19'd0;
		WeightsStore0[455] <= 19'd0;
		WeightsStore0[456] <= 19'd0;
		WeightsStore0[457] <= 19'd0;
		WeightsStore0[458] <= 19'd0;
		WeightsStore0[459] <= 19'd0;
		WeightsStore0[460] <= 19'd0;
		WeightsStore0[461] <= 19'd0;
		WeightsStore0[462] <= 19'd0;
		WeightsStore0[463] <= 19'd0;
		WeightsStore0[464] <= 19'd0;
		WeightsStore0[465] <= 19'd0;
		WeightsStore0[466] <= 19'd0;
		WeightsStore0[467] <= 19'd0;
		WeightsStore0[468] <= 19'd0;
		WeightsStore0[469] <= 19'd0;
		WeightsStore0[470] <= 19'd0;
		WeightsStore0[471] <= 19'd0;
		WeightsStore0[472] <= 19'd0;
		WeightsStore0[473] <= 19'd0;
		WeightsStore0[474] <= 19'd0;
		WeightsStore0[475] <= 19'd0;
		WeightsStore0[476] <= 19'd0;
		WeightsStore0[477] <= 19'd0;
		WeightsStore0[478] <= 19'd0;
		WeightsStore0[479] <= 19'd0;
		WeightsStore0[480] <= 19'd0;
		WeightsStore0[481] <= 19'd0;
		WeightsStore0[482] <= 19'd0;
		WeightsStore0[483] <= 19'd0;
		WeightsStore0[484] <= 19'd0;
		WeightsStore0[485] <= 19'd0;
		WeightsStore0[486] <= 19'd0;
		WeightsStore0[487] <= 19'd0;
		WeightsStore0[488] <= 19'd0;
		WeightsStore0[489] <= 19'd0;
		WeightsStore0[490] <= 19'd0;
		WeightsStore0[491] <= 19'd0;
		WeightsStore0[492] <= 19'd0;
		WeightsStore0[493] <= 19'd0;
		WeightsStore0[494] <= 19'd0;
		WeightsStore0[495] <= 19'd0;
		WeightsStore0[496] <= 19'd0;
		WeightsStore0[497] <= 19'd0;
		WeightsStore0[498] <= 19'd0;
		WeightsStore0[499] <= 19'd0;
		WeightsStore0[500] <= 19'd0;
		WeightsStore0[501] <= 19'd0;
		WeightsStore0[502] <= 19'd0;
		WeightsStore0[503] <= 19'd0;
		WeightsStore0[504] <= 19'd0;
		WeightsStore0[505] <= 19'd0;
		WeightsStore0[506] <= 19'd0;
		WeightsStore0[507] <= 19'd0;
		WeightsStore0[508] <= 19'd0;
		WeightsStore0[509] <= 19'd0;
		WeightsStore0[510] <= 19'd0;
		WeightsStore0[511] <= 19'd0;
		WeightsStore0[512] <= 19'd0;
		WeightsStore0[513] <= 19'd0;
		WeightsStore0[514] <= 19'd0;
		WeightsStore0[515] <= 19'd0;
		WeightsStore0[516] <= 19'd0;
		WeightsStore0[517] <= 19'd0;
		WeightsStore0[518] <= 19'd0;
		WeightsStore0[519] <= 19'd0;
		WeightsStore0[520] <= 19'd0;
		WeightsStore0[521] <= 19'd0;
		WeightsStore0[522] <= 19'd0;
		WeightsStore0[523] <= 19'd0;
		WeightsStore0[524] <= 19'd0;
		WeightsStore0[525] <= 19'd0;
		WeightsStore0[526] <= 19'd0;
		WeightsStore0[527] <= 19'd0;
		WeightsStore0[528] <= 19'd0;
		WeightsStore0[529] <= 19'd0;
		WeightsStore0[530] <= 19'd0;
		WeightsStore0[531] <= 19'd0;
		WeightsStore0[532] <= 19'd0;
		WeightsStore0[533] <= 19'd0;
		WeightsStore0[534] <= 19'd0;
		WeightsStore0[535] <= 19'd0;
		WeightsStore0[536] <= 19'd0;
		WeightsStore0[537] <= 19'd0;
		WeightsStore0[538] <= 19'd0;
		WeightsStore0[539] <= 19'd0;
		WeightsStore0[540] <= 19'd0;
		WeightsStore0[541] <= 19'd0;
		WeightsStore0[542] <= 19'd0;
		WeightsStore0[543] <= 19'd0;
		WeightsStore0[544] <= 19'd0;
		WeightsStore0[545] <= 19'd0;
		WeightsStore0[546] <= 19'd0;
		WeightsStore0[547] <= 19'd0;
		WeightsStore0[548] <= 19'd0;
		WeightsStore0[549] <= 19'd0;
		WeightsStore0[550] <= 19'd0;
		WeightsStore0[551] <= 19'd0;
		WeightsStore0[552] <= 19'd0;
		WeightsStore0[553] <= 19'd0;
		WeightsStore0[554] <= 19'd0;
		WeightsStore0[555] <= 19'd0;
		WeightsStore0[556] <= 19'd0;
		WeightsStore0[557] <= 19'd0;
		WeightsStore0[558] <= 19'd0;
		WeightsStore0[559] <= 19'd0;
		WeightsStore0[560] <= 19'd0;
		WeightsStore0[561] <= 19'd0;
		WeightsStore0[562] <= 19'd0;
		WeightsStore0[563] <= 19'd0;
		WeightsStore0[564] <= 19'd0;
		WeightsStore0[565] <= 19'd0;
		WeightsStore0[566] <= 19'd0;
		WeightsStore0[567] <= 19'd0;
		WeightsStore0[568] <= 19'd0;
		WeightsStore0[569] <= 19'd0;
		WeightsStore0[570] <= 19'd0;
		WeightsStore0[571] <= 19'd0;
		WeightsStore0[572] <= 19'd0;
		WeightsStore0[573] <= 19'd0;
		WeightsStore0[574] <= 19'd0;
		WeightsStore0[575] <= 19'd0;
		WeightsStore0[576] <= 19'd0;
		WeightsStore0[577] <= 19'd0;
		WeightsStore0[578] <= 19'd0;
		WeightsStore0[579] <= 19'd0;
		WeightsStore0[580] <= 19'd0;
		WeightsStore0[581] <= 19'd0;
		WeightsStore0[582] <= 19'd0;
		WeightsStore0[583] <= 19'd0;
		WeightsStore0[584] <= 19'd0;
		WeightsStore0[585] <= 19'd0;
		WeightsStore0[586] <= 19'd0;
		WeightsStore0[587] <= 19'd0;
		WeightsStore0[588] <= 19'd0;
		WeightsStore0[589] <= 19'd0;
		WeightsStore0[590] <= 19'd0;
		WeightsStore0[591] <= 19'd0;
		WeightsStore0[592] <= 19'd0;
		WeightsStore0[593] <= 19'd0;
		WeightsStore0[594] <= 19'd0;
		WeightsStore0[595] <= 19'd0;
		WeightsStore0[596] <= 19'd0;
		WeightsStore0[597] <= 19'd0;
		WeightsStore0[598] <= 19'd0;
		WeightsStore0[599] <= 19'd0;
		WeightsStore0[600] <= 19'd0;
		WeightsStore0[601] <= 19'd0;
		WeightsStore0[602] <= 19'd0;
		WeightsStore0[603] <= 19'd0;
		WeightsStore0[604] <= 19'd0;
		WeightsStore0[605] <= 19'd0;
		WeightsStore0[606] <= 19'd0;
		WeightsStore0[607] <= 19'd0;
		WeightsStore0[608] <= 19'd0;
		WeightsStore0[609] <= 19'd0;
		WeightsStore0[610] <= 19'd0;
		WeightsStore0[611] <= 19'd0;
		WeightsStore0[612] <= 19'd0;
		WeightsStore0[613] <= 19'd0;
		WeightsStore0[614] <= 19'd0;
		WeightsStore0[615] <= 19'd0;
		WeightsStore0[616] <= 19'd0;
		WeightsStore0[617] <= 19'd0;
		WeightsStore0[618] <= 19'd0;
		WeightsStore0[619] <= 19'd0;
		WeightsStore0[620] <= 19'd0;
		WeightsStore0[621] <= 19'd0;
		WeightsStore0[622] <= 19'd0;
		WeightsStore0[623] <= 19'd0;
		WeightsStore0[624] <= 19'd0;
		WeightsStore0[625] <= 19'd0;
		WeightsStore0[626] <= 19'd0;
		WeightsStore0[627] <= 19'd0;
		WeightsStore0[628] <= 19'd0;
		WeightsStore0[629] <= 19'd0;
		WeightsStore0[630] <= 19'd0;
		WeightsStore0[631] <= 19'd0;
		WeightsStore0[632] <= 19'd0;
		WeightsStore0[633] <= 19'd0;
		WeightsStore0[634] <= 19'd0;
		WeightsStore0[635] <= 19'd0;
		WeightsStore0[636] <= 19'd0;
		WeightsStore0[637] <= 19'd0;
		WeightsStore0[638] <= 19'd0;
		WeightsStore0[639] <= 19'd0;
		WeightsStore0[640] <= 19'd0;
		WeightsStore0[641] <= 19'd0;
		WeightsStore0[642] <= 19'd0;
		WeightsStore0[643] <= 19'd0;
		WeightsStore0[644] <= 19'd0;
		WeightsStore0[645] <= 19'd0;
		WeightsStore0[646] <= 19'd0;
		WeightsStore0[647] <= 19'd0;
		WeightsStore0[648] <= 19'd0;
		WeightsStore0[649] <= 19'd0;
		WeightsStore0[650] <= 19'd0;
		WeightsStore0[651] <= 19'd0;
		WeightsStore0[652] <= 19'd0;
		WeightsStore0[653] <= 19'd0;
		WeightsStore0[654] <= 19'd0;
		WeightsStore0[655] <= 19'd0;
		WeightsStore0[656] <= 19'd0;
		WeightsStore0[657] <= 19'd0;
		WeightsStore0[658] <= 19'd0;
		WeightsStore0[659] <= 19'd0;
		WeightsStore0[660] <= 19'd0;
		WeightsStore0[661] <= 19'd0;
		WeightsStore0[662] <= 19'd0;
		WeightsStore0[663] <= 19'd0;
		WeightsStore0[664] <= 19'd0;
		WeightsStore0[665] <= 19'd0;
		WeightsStore0[666] <= 19'd0;
		WeightsStore0[667] <= 19'd0;
		WeightsStore0[668] <= 19'd0;
		WeightsStore0[669] <= 19'd0;
		WeightsStore0[670] <= 19'd0;
		WeightsStore0[671] <= 19'd0;
		WeightsStore0[672] <= 19'd0;
		WeightsStore0[673] <= 19'd0;
		WeightsStore0[674] <= 19'd0;
		WeightsStore0[675] <= 19'd0;
		WeightsStore0[676] <= 19'd0;
		WeightsStore0[677] <= 19'd0;
		WeightsStore0[678] <= 19'd0;
		WeightsStore0[679] <= 19'd0;
		WeightsStore0[680] <= 19'd0;
		WeightsStore0[681] <= 19'd0;
		WeightsStore0[682] <= 19'd0;
		WeightsStore0[683] <= 19'd0;
		WeightsStore0[684] <= 19'd0;
		WeightsStore0[685] <= 19'd0;
		WeightsStore0[686] <= 19'd0;
		WeightsStore0[687] <= 19'd0;
		WeightsStore0[688] <= 19'd0;
		WeightsStore0[689] <= 19'd0;
		WeightsStore0[690] <= 19'd0;
		WeightsStore0[691] <= 19'd0;
		WeightsStore0[692] <= 19'd0;
		WeightsStore0[693] <= 19'd0;
		WeightsStore0[694] <= 19'd0;
		WeightsStore0[695] <= 19'd0;
		WeightsStore0[696] <= 19'd0;
		WeightsStore0[697] <= 19'd0;
		WeightsStore0[698] <= 19'd0;
		WeightsStore0[699] <= 19'd0;
		WeightsStore0[700] <= 19'd0;
		WeightsStore0[701] <= 19'd0;
		WeightsStore0[702] <= 19'd0;
		WeightsStore0[703] <= 19'd0;
		WeightsStore0[704] <= 19'd0;
		WeightsStore0[705] <= 19'd0;
		WeightsStore0[706] <= 19'd0;
		WeightsStore0[707] <= 19'd0;
		WeightsStore0[708] <= 19'd0;
		WeightsStore0[709] <= 19'd0;
		WeightsStore0[710] <= 19'd0;
		WeightsStore0[711] <= 19'd0;
		WeightsStore0[712] <= 19'd0;
		WeightsStore0[713] <= 19'd0;
		WeightsStore0[714] <= 19'd0;
		WeightsStore0[715] <= 19'd0;
		WeightsStore0[716] <= 19'd0;
		WeightsStore0[717] <= 19'd0;
		WeightsStore0[718] <= 19'd0;
		WeightsStore0[719] <= 19'd0;
		WeightsStore0[720] <= 19'd0;
		WeightsStore0[721] <= 19'd0;
		WeightsStore0[722] <= 19'd0;
		WeightsStore0[723] <= 19'd0;
		WeightsStore0[724] <= 19'd0;
		WeightsStore0[725] <= 19'd0;
		WeightsStore0[726] <= 19'd0;
		WeightsStore0[727] <= 19'd0;
		WeightsStore0[728] <= 19'd0;
		WeightsStore0[729] <= 19'd0;
		WeightsStore0[730] <= 19'd0;
		WeightsStore0[731] <= 19'd0;
		WeightsStore0[732] <= 19'd0;
		WeightsStore0[733] <= 19'd0;
		WeightsStore0[734] <= 19'd0;
		WeightsStore0[735] <= 19'd0;
		WeightsStore0[736] <= 19'd0;
		WeightsStore0[737] <= 19'd0;
		WeightsStore0[738] <= 19'd0;
		WeightsStore0[739] <= 19'd0;
		WeightsStore0[740] <= 19'd0;
		WeightsStore0[741] <= 19'd0;
		WeightsStore0[742] <= 19'd0;
		WeightsStore0[743] <= 19'd0;
		WeightsStore0[744] <= 19'd0;
		WeightsStore0[745] <= 19'd0;
		WeightsStore0[746] <= 19'd0;
		WeightsStore0[747] <= 19'd0;
		WeightsStore0[748] <= 19'd0;
		WeightsStore0[749] <= 19'd0;
		WeightsStore0[750] <= 19'd0;
		WeightsStore0[751] <= 19'd0;
		WeightsStore0[752] <= 19'd0;
		WeightsStore0[753] <= 19'd0;
		WeightsStore0[754] <= 19'd0;
		WeightsStore0[755] <= 19'd0;
		WeightsStore0[756] <= 19'd0;
		WeightsStore0[757] <= 19'd0;
		WeightsStore0[758] <= 19'd0;
		WeightsStore0[759] <= 19'd0;
		WeightsStore0[760] <= 19'd0;
		WeightsStore0[761] <= 19'd0;
		WeightsStore0[762] <= 19'd0;
		WeightsStore0[763] <= 19'd0;
		WeightsStore0[764] <= 19'd0;
		WeightsStore0[765] <= 19'd0;
		WeightsStore0[766] <= 19'd0;
		WeightsStore0[767] <= 19'd0;
		WeightsStore0[768] <= 19'd0;
		WeightsStore0[769] <= 19'd0;
		WeightsStore0[770] <= 19'd0;
		WeightsStore0[771] <= 19'd0;
		WeightsStore0[772] <= 19'd0;
		WeightsStore0[773] <= 19'd0;
		WeightsStore0[774] <= 19'd0;
		WeightsStore0[775] <= 19'd0;
		WeightsStore0[776] <= 19'd0;
		WeightsStore0[777] <= 19'd0;
		WeightsStore0[778] <= 19'd0;
		WeightsStore0[779] <= 19'd0;
		WeightsStore0[780] <= 19'd0;
		WeightsStore0[781] <= 19'd0;
		WeightsStore0[782] <= 19'd0;
		WeightsStore0[783] <= 19'd0;
		WeightsStore0[784] <= 19'd0;
		WeightsStore1[0] <= 19'd0;
		WeightsStore1[1] <= 19'd0;
		WeightsStore1[2] <= 19'd0;
		WeightsStore1[3] <= 19'd0;
		WeightsStore1[4] <= 19'd0;
		WeightsStore1[5] <= 19'd0;
		WeightsStore1[6] <= 19'd0;
		WeightsStore1[7] <= 19'd0;
		WeightsStore1[8] <= 19'd0;
		WeightsStore1[9] <= 19'd0;
		WeightsStore1[10] <= 19'd0;
		WeightsStore1[11] <= 19'd0;
		WeightsStore1[12] <= 19'd0;
		WeightsStore1[13] <= 19'd0;
		WeightsStore1[14] <= 19'd0;
		WeightsStore1[15] <= 19'd0;
		WeightsStore1[16] <= 19'd0;
		WeightsStore1[17] <= 19'd0;
		WeightsStore1[18] <= 19'd0;
		WeightsStore1[19] <= 19'd0;
		WeightsStore1[20] <= 19'd0;
		WeightsStore1[21] <= 19'd0;
		WeightsStore1[22] <= 19'd0;
		WeightsStore1[23] <= 19'd0;
		WeightsStore1[24] <= 19'd0;
		WeightsStore1[25] <= 19'd0;
		WeightsStore1[26] <= 19'd0;
		WeightsStore1[27] <= 19'd0;
		WeightsStore1[28] <= 19'd0;
		WeightsStore1[29] <= 19'd0;
		WeightsStore1[30] <= 19'd0;
		WeightsStore1[31] <= 19'd0;
		WeightsStore1[32] <= 19'd0;
		WeightsStore1[33] <= 19'd0;
		WeightsStore1[34] <= 19'd0;
		WeightsStore1[35] <= 19'd0;
		WeightsStore1[36] <= 19'd0;
		WeightsStore1[37] <= 19'd0;
		WeightsStore1[38] <= 19'd0;
		WeightsStore1[39] <= 19'd0;
		WeightsStore1[40] <= 19'd0;
		WeightsStore1[41] <= 19'd0;
		WeightsStore1[42] <= 19'd0;
		WeightsStore1[43] <= 19'd0;
		WeightsStore1[44] <= 19'd0;
		WeightsStore1[45] <= 19'd0;
		WeightsStore1[46] <= 19'd0;
		WeightsStore1[47] <= 19'd0;
		WeightsStore1[48] <= 19'd0;
		WeightsStore1[49] <= 19'd0;
		WeightsStore1[50] <= 19'd0;
		WeightsStore1[51] <= 19'd0;
		WeightsStore1[52] <= 19'd0;
		WeightsStore1[53] <= 19'd0;
		WeightsStore1[54] <= 19'd0;
		WeightsStore1[55] <= 19'd0;
		WeightsStore1[56] <= 19'd0;
		WeightsStore1[57] <= 19'd0;
		WeightsStore1[58] <= 19'd0;
		WeightsStore1[59] <= 19'd0;
		WeightsStore1[60] <= 19'd0;
		WeightsStore1[61] <= 19'd0;
		WeightsStore1[62] <= 19'd0;
		WeightsStore1[63] <= 19'd0;
		WeightsStore1[64] <= 19'd0;
		WeightsStore1[65] <= 19'd0;
		WeightsStore1[66] <= 19'd0;
		WeightsStore1[67] <= 19'd0;
		WeightsStore1[68] <= 19'd0;
		WeightsStore1[69] <= 19'd0;
		WeightsStore1[70] <= 19'd0;
		WeightsStore1[71] <= 19'd0;
		WeightsStore1[72] <= 19'd0;
		WeightsStore1[73] <= 19'd0;
		WeightsStore1[74] <= 19'd0;
		WeightsStore1[75] <= 19'd0;
		WeightsStore1[76] <= 19'd0;
		WeightsStore1[77] <= 19'd0;
		WeightsStore1[78] <= 19'd0;
		WeightsStore1[79] <= 19'd0;
		WeightsStore1[80] <= 19'd0;
		WeightsStore1[81] <= 19'd0;
		WeightsStore1[82] <= 19'd0;
		WeightsStore1[83] <= 19'd0;
		WeightsStore1[84] <= 19'd0;
		WeightsStore1[85] <= 19'd0;
		WeightsStore1[86] <= 19'd0;
		WeightsStore1[87] <= 19'd0;
		WeightsStore1[88] <= 19'd0;
		WeightsStore1[89] <= 19'd0;
		WeightsStore1[90] <= 19'd0;
		WeightsStore1[91] <= 19'd0;
		WeightsStore1[92] <= 19'd0;
		WeightsStore1[93] <= 19'd0;
		WeightsStore1[94] <= 19'd0;
		WeightsStore1[95] <= 19'd0;
		WeightsStore1[96] <= 19'd0;
		WeightsStore1[97] <= 19'd0;
		WeightsStore1[98] <= 19'd0;
		WeightsStore1[99] <= 19'd0;
		WeightsStore1[100] <= 19'd0;
		WeightsStore1[101] <= 19'd0;
		WeightsStore1[102] <= 19'd0;
		WeightsStore1[103] <= 19'd0;
		WeightsStore1[104] <= 19'd0;
		WeightsStore1[105] <= 19'd0;
		WeightsStore1[106] <= 19'd0;
		WeightsStore1[107] <= 19'd0;
		WeightsStore1[108] <= 19'd0;
		WeightsStore1[109] <= 19'd0;
		WeightsStore1[110] <= 19'd0;
		WeightsStore1[111] <= 19'd0;
		WeightsStore1[112] <= 19'd0;
		WeightsStore1[113] <= 19'd0;
		WeightsStore1[114] <= 19'd0;
		WeightsStore1[115] <= 19'd0;
		WeightsStore1[116] <= 19'd0;
		WeightsStore1[117] <= 19'd0;
		WeightsStore1[118] <= 19'd0;
		WeightsStore1[119] <= 19'd0;
		WeightsStore1[120] <= 19'd0;
		WeightsStore1[121] <= 19'd0;
		WeightsStore1[122] <= 19'd0;
		WeightsStore1[123] <= 19'd0;
		WeightsStore1[124] <= 19'd0;
		WeightsStore1[125] <= 19'd0;
		WeightsStore1[126] <= 19'd0;
		WeightsStore1[127] <= 19'd0;
		WeightsStore1[128] <= 19'd0;
		WeightsStore1[129] <= 19'd0;
		WeightsStore1[130] <= 19'd0;
		WeightsStore1[131] <= 19'd0;
		WeightsStore1[132] <= 19'd0;
		WeightsStore1[133] <= 19'd0;
		WeightsStore1[134] <= 19'd0;
		WeightsStore1[135] <= 19'd0;
		WeightsStore1[136] <= 19'd0;
		WeightsStore1[137] <= 19'd0;
		WeightsStore1[138] <= 19'd0;
		WeightsStore1[139] <= 19'd0;
		WeightsStore1[140] <= 19'd0;
		WeightsStore1[141] <= 19'd0;
		WeightsStore1[142] <= 19'd0;
		WeightsStore1[143] <= 19'd0;
		WeightsStore1[144] <= 19'd0;
		WeightsStore1[145] <= 19'd0;
		WeightsStore1[146] <= 19'd0;
		WeightsStore1[147] <= 19'd0;
		WeightsStore1[148] <= 19'd0;
		WeightsStore1[149] <= 19'd0;
		WeightsStore1[150] <= 19'd0;
		WeightsStore1[151] <= 19'd0;
		WeightsStore1[152] <= 19'd0;
		WeightsStore1[153] <= 19'd0;
		WeightsStore1[154] <= 19'd0;
		WeightsStore1[155] <= 19'd0;
		WeightsStore1[156] <= 19'd0;
		WeightsStore1[157] <= 19'd0;
		WeightsStore1[158] <= 19'd0;
		WeightsStore1[159] <= 19'd0;
		WeightsStore1[160] <= 19'd0;
		WeightsStore1[161] <= 19'd0;
		WeightsStore1[162] <= 19'd0;
		WeightsStore1[163] <= 19'd0;
		WeightsStore1[164] <= 19'd0;
		WeightsStore1[165] <= 19'd0;
		WeightsStore1[166] <= 19'd0;
		WeightsStore1[167] <= 19'd0;
		WeightsStore1[168] <= 19'd0;
		WeightsStore1[169] <= 19'd0;
		WeightsStore1[170] <= 19'd0;
		WeightsStore1[171] <= 19'd0;
		WeightsStore1[172] <= 19'd0;
		WeightsStore1[173] <= 19'd0;
		WeightsStore1[174] <= 19'd0;
		WeightsStore1[175] <= 19'd0;
		WeightsStore1[176] <= 19'd0;
		WeightsStore1[177] <= 19'd0;
		WeightsStore1[178] <= 19'd0;
		WeightsStore1[179] <= 19'd0;
		WeightsStore1[180] <= 19'd0;
		WeightsStore1[181] <= 19'd0;
		WeightsStore1[182] <= 19'd0;
		WeightsStore1[183] <= 19'd0;
		WeightsStore1[184] <= 19'd0;
		WeightsStore1[185] <= 19'd0;
		WeightsStore1[186] <= 19'd0;
		WeightsStore1[187] <= 19'd0;
		WeightsStore1[188] <= 19'd0;
		WeightsStore1[189] <= 19'd0;
		WeightsStore1[190] <= 19'd0;
		WeightsStore1[191] <= 19'd0;
		WeightsStore1[192] <= 19'd0;
		WeightsStore1[193] <= 19'd0;
		WeightsStore1[194] <= 19'd0;
		WeightsStore1[195] <= 19'd0;
		WeightsStore1[196] <= 19'd0;
		WeightsStore1[197] <= 19'd0;
		WeightsStore1[198] <= 19'd0;
		WeightsStore1[199] <= 19'd0;
		WeightsStore1[200] <= 19'd0;
		WeightsStore1[201] <= 19'd0;
		WeightsStore1[202] <= 19'd0;
		WeightsStore1[203] <= 19'd0;
		WeightsStore1[204] <= 19'd0;
		WeightsStore1[205] <= 19'd0;
		WeightsStore1[206] <= 19'd0;
		WeightsStore1[207] <= 19'd0;
		WeightsStore1[208] <= 19'd0;
		WeightsStore1[209] <= 19'd0;
		WeightsStore1[210] <= 19'd0;
		WeightsStore1[211] <= 19'd0;
		WeightsStore1[212] <= 19'd0;
		WeightsStore1[213] <= 19'd0;
		WeightsStore1[214] <= 19'd0;
		WeightsStore1[215] <= 19'd0;
		WeightsStore1[216] <= 19'd0;
		WeightsStore1[217] <= 19'd0;
		WeightsStore1[218] <= 19'd0;
		WeightsStore1[219] <= 19'd0;
		WeightsStore1[220] <= 19'd0;
		WeightsStore1[221] <= 19'd0;
		WeightsStore1[222] <= 19'd0;
		WeightsStore1[223] <= 19'd0;
		WeightsStore1[224] <= 19'd0;
		WeightsStore1[225] <= 19'd0;
		WeightsStore1[226] <= 19'd0;
		WeightsStore1[227] <= 19'd0;
		WeightsStore1[228] <= 19'd0;
		WeightsStore1[229] <= 19'd0;
		WeightsStore1[230] <= 19'd0;
		WeightsStore1[231] <= 19'd0;
		WeightsStore1[232] <= 19'd0;
		WeightsStore1[233] <= 19'd0;
		WeightsStore1[234] <= 19'd0;
		WeightsStore1[235] <= 19'd0;
		WeightsStore1[236] <= 19'd0;
		WeightsStore1[237] <= 19'd0;
		WeightsStore1[238] <= 19'd0;
		WeightsStore1[239] <= 19'd0;
		WeightsStore1[240] <= 19'd0;
		WeightsStore1[241] <= 19'd0;
		WeightsStore1[242] <= 19'd0;
		WeightsStore1[243] <= 19'd0;
		WeightsStore1[244] <= 19'd0;
		WeightsStore1[245] <= 19'd0;
		WeightsStore1[246] <= 19'd0;
		WeightsStore1[247] <= 19'd0;
		WeightsStore1[248] <= 19'd0;
		WeightsStore1[249] <= 19'd0;
		WeightsStore1[250] <= 19'd0;
		WeightsStore1[251] <= 19'd0;
		WeightsStore1[252] <= 19'd0;
		WeightsStore1[253] <= 19'd0;
		WeightsStore1[254] <= 19'd0;
		WeightsStore1[255] <= 19'd0;
		WeightsStore1[256] <= 19'd0;
		WeightsStore1[257] <= 19'd0;
		WeightsStore1[258] <= 19'd0;
		WeightsStore1[259] <= 19'd0;
		WeightsStore1[260] <= 19'd0;
		WeightsStore1[261] <= 19'd0;
		WeightsStore1[262] <= 19'd0;
		WeightsStore1[263] <= 19'd0;
		WeightsStore1[264] <= 19'd0;
		WeightsStore1[265] <= 19'd0;
		WeightsStore1[266] <= 19'd0;
		WeightsStore1[267] <= 19'd0;
		WeightsStore1[268] <= 19'd0;
		WeightsStore1[269] <= 19'd0;
		WeightsStore1[270] <= 19'd0;
		WeightsStore1[271] <= 19'd0;
		WeightsStore1[272] <= 19'd0;
		WeightsStore1[273] <= 19'd0;
		WeightsStore1[274] <= 19'd0;
		WeightsStore1[275] <= 19'd0;
		WeightsStore1[276] <= 19'd0;
		WeightsStore1[277] <= 19'd0;
		WeightsStore1[278] <= 19'd0;
		WeightsStore1[279] <= 19'd0;
		WeightsStore1[280] <= 19'd0;
		WeightsStore1[281] <= 19'd0;
		WeightsStore1[282] <= 19'd0;
		WeightsStore1[283] <= 19'd0;
		WeightsStore1[284] <= 19'd0;
		WeightsStore1[285] <= 19'd0;
		WeightsStore1[286] <= 19'd0;
		WeightsStore1[287] <= 19'd0;
		WeightsStore1[288] <= 19'd0;
		WeightsStore1[289] <= 19'd0;
		WeightsStore1[290] <= 19'd0;
		WeightsStore1[291] <= 19'd0;
		WeightsStore1[292] <= 19'd0;
		WeightsStore1[293] <= 19'd0;
		WeightsStore1[294] <= 19'd0;
		WeightsStore1[295] <= 19'd0;
		WeightsStore1[296] <= 19'd0;
		WeightsStore1[297] <= 19'd0;
		WeightsStore1[298] <= 19'd0;
		WeightsStore1[299] <= 19'd0;
		WeightsStore1[300] <= 19'd0;
		WeightsStore1[301] <= 19'd0;
		WeightsStore1[302] <= 19'd0;
		WeightsStore1[303] <= 19'd0;
		WeightsStore1[304] <= 19'd0;
		WeightsStore1[305] <= 19'd0;
		WeightsStore1[306] <= 19'd0;
		WeightsStore1[307] <= 19'd0;
		WeightsStore1[308] <= 19'd0;
		WeightsStore1[309] <= 19'd0;
		WeightsStore1[310] <= 19'd0;
		WeightsStore1[311] <= 19'd0;
		WeightsStore1[312] <= 19'd0;
		WeightsStore1[313] <= 19'd0;
		WeightsStore1[314] <= 19'd0;
		WeightsStore1[315] <= 19'd0;
		WeightsStore1[316] <= 19'd0;
		WeightsStore1[317] <= 19'd0;
		WeightsStore1[318] <= 19'd0;
		WeightsStore1[319] <= 19'd0;
		WeightsStore1[320] <= 19'd0;
		WeightsStore1[321] <= 19'd0;
		WeightsStore1[322] <= 19'd0;
		WeightsStore1[323] <= 19'd0;
		WeightsStore1[324] <= 19'd0;
		WeightsStore1[325] <= 19'd0;
		WeightsStore1[326] <= 19'd0;
		WeightsStore1[327] <= 19'd0;
		WeightsStore1[328] <= 19'd0;
		WeightsStore1[329] <= 19'd0;
		WeightsStore1[330] <= 19'd0;
		WeightsStore1[331] <= 19'd0;
		WeightsStore1[332] <= 19'd0;
		WeightsStore1[333] <= 19'd0;
		WeightsStore1[334] <= 19'd0;
		WeightsStore1[335] <= 19'd0;
		WeightsStore1[336] <= 19'd0;
		WeightsStore1[337] <= 19'd0;
		WeightsStore1[338] <= 19'd0;
		WeightsStore1[339] <= 19'd0;
		WeightsStore1[340] <= 19'd0;
		WeightsStore1[341] <= 19'd0;
		WeightsStore1[342] <= 19'd0;
		WeightsStore1[343] <= 19'd0;
		WeightsStore1[344] <= 19'd0;
		WeightsStore1[345] <= 19'd0;
		WeightsStore1[346] <= 19'd0;
		WeightsStore1[347] <= 19'd0;
		WeightsStore1[348] <= 19'd0;
		WeightsStore1[349] <= 19'd0;
		WeightsStore1[350] <= 19'd0;
		WeightsStore1[351] <= 19'd0;
		WeightsStore1[352] <= 19'd0;
		WeightsStore1[353] <= 19'd0;
		WeightsStore1[354] <= 19'd0;
		WeightsStore1[355] <= 19'd0;
		WeightsStore1[356] <= 19'd0;
		WeightsStore1[357] <= 19'd0;
		WeightsStore1[358] <= 19'd0;
		WeightsStore1[359] <= 19'd0;
		WeightsStore1[360] <= 19'd0;
		WeightsStore1[361] <= 19'd0;
		WeightsStore1[362] <= 19'd0;
		WeightsStore1[363] <= 19'd0;
		WeightsStore1[364] <= 19'd0;
		WeightsStore1[365] <= 19'd0;
		WeightsStore1[366] <= 19'd0;
		WeightsStore1[367] <= 19'd0;
		WeightsStore1[368] <= 19'd0;
		WeightsStore1[369] <= 19'd0;
		WeightsStore1[370] <= 19'd0;
		WeightsStore1[371] <= 19'd0;
		WeightsStore1[372] <= 19'd0;
		WeightsStore1[373] <= 19'd0;
		WeightsStore1[374] <= 19'd0;
		WeightsStore1[375] <= 19'd0;
		WeightsStore1[376] <= 19'd0;
		WeightsStore1[377] <= 19'd0;
		WeightsStore1[378] <= 19'd0;
		WeightsStore1[379] <= 19'd0;
		WeightsStore1[380] <= 19'd0;
		WeightsStore1[381] <= 19'd0;
		WeightsStore1[382] <= 19'd0;
		WeightsStore1[383] <= 19'd0;
		WeightsStore1[384] <= 19'd0;
		WeightsStore1[385] <= 19'd0;
		WeightsStore1[386] <= 19'd0;
		WeightsStore1[387] <= 19'd0;
		WeightsStore1[388] <= 19'd0;
		WeightsStore1[389] <= 19'd0;
		WeightsStore1[390] <= 19'd0;
		WeightsStore1[391] <= 19'd0;
		WeightsStore1[392] <= 19'd0;
		WeightsStore1[393] <= 19'd0;
		WeightsStore1[394] <= 19'd0;
		WeightsStore1[395] <= 19'd0;
		WeightsStore1[396] <= 19'd0;
		WeightsStore1[397] <= 19'd0;
		WeightsStore1[398] <= 19'd0;
		WeightsStore1[399] <= 19'd0;
		WeightsStore1[400] <= 19'd0;
		WeightsStore1[401] <= 19'd0;
		WeightsStore1[402] <= 19'd0;
		WeightsStore1[403] <= 19'd0;
		WeightsStore1[404] <= 19'd0;
		WeightsStore1[405] <= 19'd0;
		WeightsStore1[406] <= 19'd0;
		WeightsStore1[407] <= 19'd0;
		WeightsStore1[408] <= 19'd0;
		WeightsStore1[409] <= 19'd0;
		WeightsStore1[410] <= 19'd0;
		WeightsStore1[411] <= 19'd0;
		WeightsStore1[412] <= 19'd0;
		WeightsStore1[413] <= 19'd0;
		WeightsStore1[414] <= 19'd0;
		WeightsStore1[415] <= 19'd0;
		WeightsStore1[416] <= 19'd0;
		WeightsStore1[417] <= 19'd0;
		WeightsStore1[418] <= 19'd0;
		WeightsStore1[419] <= 19'd0;
		WeightsStore1[420] <= 19'd0;
		WeightsStore1[421] <= 19'd0;
		WeightsStore1[422] <= 19'd0;
		WeightsStore1[423] <= 19'd0;
		WeightsStore1[424] <= 19'd0;
		WeightsStore1[425] <= 19'd0;
		WeightsStore1[426] <= 19'd0;
		WeightsStore1[427] <= 19'd0;
		WeightsStore1[428] <= 19'd0;
		WeightsStore1[429] <= 19'd0;
		WeightsStore1[430] <= 19'd0;
		WeightsStore1[431] <= 19'd0;
		WeightsStore1[432] <= 19'd0;
		WeightsStore1[433] <= 19'd0;
		WeightsStore1[434] <= 19'd0;
		WeightsStore1[435] <= 19'd0;
		WeightsStore1[436] <= 19'd0;
		WeightsStore1[437] <= 19'd0;
		WeightsStore1[438] <= 19'd0;
		WeightsStore1[439] <= 19'd0;
		WeightsStore1[440] <= 19'd0;
		WeightsStore1[441] <= 19'd0;
		WeightsStore1[442] <= 19'd0;
		WeightsStore1[443] <= 19'd0;
		WeightsStore1[444] <= 19'd0;
		WeightsStore1[445] <= 19'd0;
		WeightsStore1[446] <= 19'd0;
		WeightsStore1[447] <= 19'd0;
		WeightsStore1[448] <= 19'd0;
		WeightsStore1[449] <= 19'd0;
		WeightsStore1[450] <= 19'd0;
		WeightsStore1[451] <= 19'd0;
		WeightsStore1[452] <= 19'd0;
		WeightsStore1[453] <= 19'd0;
		WeightsStore1[454] <= 19'd0;
		WeightsStore1[455] <= 19'd0;
		WeightsStore1[456] <= 19'd0;
		WeightsStore1[457] <= 19'd0;
		WeightsStore1[458] <= 19'd0;
		WeightsStore1[459] <= 19'd0;
		WeightsStore1[460] <= 19'd0;
		WeightsStore1[461] <= 19'd0;
		WeightsStore1[462] <= 19'd0;
		WeightsStore1[463] <= 19'd0;
		WeightsStore1[464] <= 19'd0;
		WeightsStore1[465] <= 19'd0;
		WeightsStore1[466] <= 19'd0;
		WeightsStore1[467] <= 19'd0;
		WeightsStore1[468] <= 19'd0;
		WeightsStore1[469] <= 19'd0;
		WeightsStore1[470] <= 19'd0;
		WeightsStore1[471] <= 19'd0;
		WeightsStore1[472] <= 19'd0;
		WeightsStore1[473] <= 19'd0;
		WeightsStore1[474] <= 19'd0;
		WeightsStore1[475] <= 19'd0;
		WeightsStore1[476] <= 19'd0;
		WeightsStore1[477] <= 19'd0;
		WeightsStore1[478] <= 19'd0;
		WeightsStore1[479] <= 19'd0;
		WeightsStore1[480] <= 19'd0;
		WeightsStore1[481] <= 19'd0;
		WeightsStore1[482] <= 19'd0;
		WeightsStore1[483] <= 19'd0;
		WeightsStore1[484] <= 19'd0;
		WeightsStore1[485] <= 19'd0;
		WeightsStore1[486] <= 19'd0;
		WeightsStore1[487] <= 19'd0;
		WeightsStore1[488] <= 19'd0;
		WeightsStore1[489] <= 19'd0;
		WeightsStore1[490] <= 19'd0;
		WeightsStore1[491] <= 19'd0;
		WeightsStore1[492] <= 19'd0;
		WeightsStore1[493] <= 19'd0;
		WeightsStore1[494] <= 19'd0;
		WeightsStore1[495] <= 19'd0;
		WeightsStore1[496] <= 19'd0;
		WeightsStore1[497] <= 19'd0;
		WeightsStore1[498] <= 19'd0;
		WeightsStore1[499] <= 19'd0;
		WeightsStore1[500] <= 19'd0;
		WeightsStore1[501] <= 19'd0;
		WeightsStore1[502] <= 19'd0;
		WeightsStore1[503] <= 19'd0;
		WeightsStore1[504] <= 19'd0;
		WeightsStore1[505] <= 19'd0;
		WeightsStore1[506] <= 19'd0;
		WeightsStore1[507] <= 19'd0;
		WeightsStore1[508] <= 19'd0;
		WeightsStore1[509] <= 19'd0;
		WeightsStore1[510] <= 19'd0;
		WeightsStore1[511] <= 19'd0;
		WeightsStore1[512] <= 19'd0;
		WeightsStore1[513] <= 19'd0;
		WeightsStore1[514] <= 19'd0;
		WeightsStore1[515] <= 19'd0;
		WeightsStore1[516] <= 19'd0;
		WeightsStore1[517] <= 19'd0;
		WeightsStore1[518] <= 19'd0;
		WeightsStore1[519] <= 19'd0;
		WeightsStore1[520] <= 19'd0;
		WeightsStore1[521] <= 19'd0;
		WeightsStore1[522] <= 19'd0;
		WeightsStore1[523] <= 19'd0;
		WeightsStore1[524] <= 19'd0;
		WeightsStore1[525] <= 19'd0;
		WeightsStore1[526] <= 19'd0;
		WeightsStore1[527] <= 19'd0;
		WeightsStore1[528] <= 19'd0;
		WeightsStore1[529] <= 19'd0;
		WeightsStore1[530] <= 19'd0;
		WeightsStore1[531] <= 19'd0;
		WeightsStore1[532] <= 19'd0;
		WeightsStore1[533] <= 19'd0;
		WeightsStore1[534] <= 19'd0;
		WeightsStore1[535] <= 19'd0;
		WeightsStore1[536] <= 19'd0;
		WeightsStore1[537] <= 19'd0;
		WeightsStore1[538] <= 19'd0;
		WeightsStore1[539] <= 19'd0;
		WeightsStore1[540] <= 19'd0;
		WeightsStore1[541] <= 19'd0;
		WeightsStore1[542] <= 19'd0;
		WeightsStore1[543] <= 19'd0;
		WeightsStore1[544] <= 19'd0;
		WeightsStore1[545] <= 19'd0;
		WeightsStore1[546] <= 19'd0;
		WeightsStore1[547] <= 19'd0;
		WeightsStore1[548] <= 19'd0;
		WeightsStore1[549] <= 19'd0;
		WeightsStore1[550] <= 19'd0;
		WeightsStore1[551] <= 19'd0;
		WeightsStore1[552] <= 19'd0;
		WeightsStore1[553] <= 19'd0;
		WeightsStore1[554] <= 19'd0;
		WeightsStore1[555] <= 19'd0;
		WeightsStore1[556] <= 19'd0;
		WeightsStore1[557] <= 19'd0;
		WeightsStore1[558] <= 19'd0;
		WeightsStore1[559] <= 19'd0;
		WeightsStore1[560] <= 19'd0;
		WeightsStore1[561] <= 19'd0;
		WeightsStore1[562] <= 19'd0;
		WeightsStore1[563] <= 19'd0;
		WeightsStore1[564] <= 19'd0;
		WeightsStore1[565] <= 19'd0;
		WeightsStore1[566] <= 19'd0;
		WeightsStore1[567] <= 19'd0;
		WeightsStore1[568] <= 19'd0;
		WeightsStore1[569] <= 19'd0;
		WeightsStore1[570] <= 19'd0;
		WeightsStore1[571] <= 19'd0;
		WeightsStore1[572] <= 19'd0;
		WeightsStore1[573] <= 19'd0;
		WeightsStore1[574] <= 19'd0;
		WeightsStore1[575] <= 19'd0;
		WeightsStore1[576] <= 19'd0;
		WeightsStore1[577] <= 19'd0;
		WeightsStore1[578] <= 19'd0;
		WeightsStore1[579] <= 19'd0;
		WeightsStore1[580] <= 19'd0;
		WeightsStore1[581] <= 19'd0;
		WeightsStore1[582] <= 19'd0;
		WeightsStore1[583] <= 19'd0;
		WeightsStore1[584] <= 19'd0;
		WeightsStore1[585] <= 19'd0;
		WeightsStore1[586] <= 19'd0;
		WeightsStore1[587] <= 19'd0;
		WeightsStore1[588] <= 19'd0;
		WeightsStore1[589] <= 19'd0;
		WeightsStore1[590] <= 19'd0;
		WeightsStore1[591] <= 19'd0;
		WeightsStore1[592] <= 19'd0;
		WeightsStore1[593] <= 19'd0;
		WeightsStore1[594] <= 19'd0;
		WeightsStore1[595] <= 19'd0;
		WeightsStore1[596] <= 19'd0;
		WeightsStore1[597] <= 19'd0;
		WeightsStore1[598] <= 19'd0;
		WeightsStore1[599] <= 19'd0;
		WeightsStore1[600] <= 19'd0;
		WeightsStore1[601] <= 19'd0;
		WeightsStore1[602] <= 19'd0;
		WeightsStore1[603] <= 19'd0;
		WeightsStore1[604] <= 19'd0;
		WeightsStore1[605] <= 19'd0;
		WeightsStore1[606] <= 19'd0;
		WeightsStore1[607] <= 19'd0;
		WeightsStore1[608] <= 19'd0;
		WeightsStore1[609] <= 19'd0;
		WeightsStore1[610] <= 19'd0;
		WeightsStore1[611] <= 19'd0;
		WeightsStore1[612] <= 19'd0;
		WeightsStore1[613] <= 19'd0;
		WeightsStore1[614] <= 19'd0;
		WeightsStore1[615] <= 19'd0;
		WeightsStore1[616] <= 19'd0;
		WeightsStore1[617] <= 19'd0;
		WeightsStore1[618] <= 19'd0;
		WeightsStore1[619] <= 19'd0;
		WeightsStore1[620] <= 19'd0;
		WeightsStore1[621] <= 19'd0;
		WeightsStore1[622] <= 19'd0;
		WeightsStore1[623] <= 19'd0;
		WeightsStore1[624] <= 19'd0;
		WeightsStore1[625] <= 19'd0;
		WeightsStore1[626] <= 19'd0;
		WeightsStore1[627] <= 19'd0;
		WeightsStore1[628] <= 19'd0;
		WeightsStore1[629] <= 19'd0;
		WeightsStore1[630] <= 19'd0;
		WeightsStore1[631] <= 19'd0;
		WeightsStore1[632] <= 19'd0;
		WeightsStore1[633] <= 19'd0;
		WeightsStore1[634] <= 19'd0;
		WeightsStore1[635] <= 19'd0;
		WeightsStore1[636] <= 19'd0;
		WeightsStore1[637] <= 19'd0;
		WeightsStore1[638] <= 19'd0;
		WeightsStore1[639] <= 19'd0;
		WeightsStore1[640] <= 19'd0;
		WeightsStore1[641] <= 19'd0;
		WeightsStore1[642] <= 19'd0;
		WeightsStore1[643] <= 19'd0;
		WeightsStore1[644] <= 19'd0;
		WeightsStore1[645] <= 19'd0;
		WeightsStore1[646] <= 19'd0;
		WeightsStore1[647] <= 19'd0;
		WeightsStore1[648] <= 19'd0;
		WeightsStore1[649] <= 19'd0;
		WeightsStore1[650] <= 19'd0;
		WeightsStore1[651] <= 19'd0;
		WeightsStore1[652] <= 19'd0;
		WeightsStore1[653] <= 19'd0;
		WeightsStore1[654] <= 19'd0;
		WeightsStore1[655] <= 19'd0;
		WeightsStore1[656] <= 19'd0;
		WeightsStore1[657] <= 19'd0;
		WeightsStore1[658] <= 19'd0;
		WeightsStore1[659] <= 19'd0;
		WeightsStore1[660] <= 19'd0;
		WeightsStore1[661] <= 19'd0;
		WeightsStore1[662] <= 19'd0;
		WeightsStore1[663] <= 19'd0;
		WeightsStore1[664] <= 19'd0;
		WeightsStore1[665] <= 19'd0;
		WeightsStore1[666] <= 19'd0;
		WeightsStore1[667] <= 19'd0;
		WeightsStore1[668] <= 19'd0;
		WeightsStore1[669] <= 19'd0;
		WeightsStore1[670] <= 19'd0;
		WeightsStore1[671] <= 19'd0;
		WeightsStore1[672] <= 19'd0;
		WeightsStore1[673] <= 19'd0;
		WeightsStore1[674] <= 19'd0;
		WeightsStore1[675] <= 19'd0;
		WeightsStore1[676] <= 19'd0;
		WeightsStore1[677] <= 19'd0;
		WeightsStore1[678] <= 19'd0;
		WeightsStore1[679] <= 19'd0;
		WeightsStore1[680] <= 19'd0;
		WeightsStore1[681] <= 19'd0;
		WeightsStore1[682] <= 19'd0;
		WeightsStore1[683] <= 19'd0;
		WeightsStore1[684] <= 19'd0;
		WeightsStore1[685] <= 19'd0;
		WeightsStore1[686] <= 19'd0;
		WeightsStore1[687] <= 19'd0;
		WeightsStore1[688] <= 19'd0;
		WeightsStore1[689] <= 19'd0;
		WeightsStore1[690] <= 19'd0;
		WeightsStore1[691] <= 19'd0;
		WeightsStore1[692] <= 19'd0;
		WeightsStore1[693] <= 19'd0;
		WeightsStore1[694] <= 19'd0;
		WeightsStore1[695] <= 19'd0;
		WeightsStore1[696] <= 19'd0;
		WeightsStore1[697] <= 19'd0;
		WeightsStore1[698] <= 19'd0;
		WeightsStore1[699] <= 19'd0;
		WeightsStore1[700] <= 19'd0;
		WeightsStore1[701] <= 19'd0;
		WeightsStore1[702] <= 19'd0;
		WeightsStore1[703] <= 19'd0;
		WeightsStore1[704] <= 19'd0;
		WeightsStore1[705] <= 19'd0;
		WeightsStore1[706] <= 19'd0;
		WeightsStore1[707] <= 19'd0;
		WeightsStore1[708] <= 19'd0;
		WeightsStore1[709] <= 19'd0;
		WeightsStore1[710] <= 19'd0;
		WeightsStore1[711] <= 19'd0;
		WeightsStore1[712] <= 19'd0;
		WeightsStore1[713] <= 19'd0;
		WeightsStore1[714] <= 19'd0;
		WeightsStore1[715] <= 19'd0;
		WeightsStore1[716] <= 19'd0;
		WeightsStore1[717] <= 19'd0;
		WeightsStore1[718] <= 19'd0;
		WeightsStore1[719] <= 19'd0;
		WeightsStore1[720] <= 19'd0;
		WeightsStore1[721] <= 19'd0;
		WeightsStore1[722] <= 19'd0;
		WeightsStore1[723] <= 19'd0;
		WeightsStore1[724] <= 19'd0;
		WeightsStore1[725] <= 19'd0;
		WeightsStore1[726] <= 19'd0;
		WeightsStore1[727] <= 19'd0;
		WeightsStore1[728] <= 19'd0;
		WeightsStore1[729] <= 19'd0;
		WeightsStore1[730] <= 19'd0;
		WeightsStore1[731] <= 19'd0;
		WeightsStore1[732] <= 19'd0;
		WeightsStore1[733] <= 19'd0;
		WeightsStore1[734] <= 19'd0;
		WeightsStore1[735] <= 19'd0;
		WeightsStore1[736] <= 19'd0;
		WeightsStore1[737] <= 19'd0;
		WeightsStore1[738] <= 19'd0;
		WeightsStore1[739] <= 19'd0;
		WeightsStore1[740] <= 19'd0;
		WeightsStore1[741] <= 19'd0;
		WeightsStore1[742] <= 19'd0;
		WeightsStore1[743] <= 19'd0;
		WeightsStore1[744] <= 19'd0;
		WeightsStore1[745] <= 19'd0;
		WeightsStore1[746] <= 19'd0;
		WeightsStore1[747] <= 19'd0;
		WeightsStore1[748] <= 19'd0;
		WeightsStore1[749] <= 19'd0;
		WeightsStore1[750] <= 19'd0;
		WeightsStore1[751] <= 19'd0;
		WeightsStore1[752] <= 19'd0;
		WeightsStore1[753] <= 19'd0;
		WeightsStore1[754] <= 19'd0;
		WeightsStore1[755] <= 19'd0;
		WeightsStore1[756] <= 19'd0;
		WeightsStore1[757] <= 19'd0;
		WeightsStore1[758] <= 19'd0;
		WeightsStore1[759] <= 19'd0;
		WeightsStore1[760] <= 19'd0;
		WeightsStore1[761] <= 19'd0;
		WeightsStore1[762] <= 19'd0;
		WeightsStore1[763] <= 19'd0;
		WeightsStore1[764] <= 19'd0;
		WeightsStore1[765] <= 19'd0;
		WeightsStore1[766] <= 19'd0;
		WeightsStore1[767] <= 19'd0;
		WeightsStore1[768] <= 19'd0;
		WeightsStore1[769] <= 19'd0;
		WeightsStore1[770] <= 19'd0;
		WeightsStore1[771] <= 19'd0;
		WeightsStore1[772] <= 19'd0;
		WeightsStore1[773] <= 19'd0;
		WeightsStore1[774] <= 19'd0;
		WeightsStore1[775] <= 19'd0;
		WeightsStore1[776] <= 19'd0;
		WeightsStore1[777] <= 19'd0;
		WeightsStore1[778] <= 19'd0;
		WeightsStore1[779] <= 19'd0;
		WeightsStore1[780] <= 19'd0;
		WeightsStore1[781] <= 19'd0;
		WeightsStore1[782] <= 19'd0;
		WeightsStore1[783] <= 19'd0;
		WeightsStore1[784] <= 19'd0;
		WeightsStore2[0] <= 19'd0;
		WeightsStore2[1] <= 19'd0;
		WeightsStore2[2] <= 19'd0;
		WeightsStore2[3] <= 19'd0;
		WeightsStore2[4] <= 19'd0;
		WeightsStore2[5] <= 19'd0;
		WeightsStore2[6] <= 19'd0;
		WeightsStore2[7] <= 19'd0;
		WeightsStore2[8] <= 19'd0;
		WeightsStore2[9] <= 19'd0;
		WeightsStore2[10] <= 19'd0;
		WeightsStore2[11] <= 19'd0;
		WeightsStore2[12] <= 19'd0;
		WeightsStore2[13] <= 19'd0;
		WeightsStore2[14] <= 19'd0;
		WeightsStore2[15] <= 19'd0;
		WeightsStore2[16] <= 19'd0;
		WeightsStore2[17] <= 19'd0;
		WeightsStore2[18] <= 19'd0;
		WeightsStore2[19] <= 19'd0;
		WeightsStore2[20] <= 19'd0;
		WeightsStore2[21] <= 19'd0;
		WeightsStore2[22] <= 19'd0;
		WeightsStore2[23] <= 19'd0;
		WeightsStore2[24] <= 19'd0;
		WeightsStore2[25] <= 19'd0;
		WeightsStore2[26] <= 19'd0;
		WeightsStore2[27] <= 19'd0;
		WeightsStore2[28] <= 19'd0;
		WeightsStore2[29] <= 19'd0;
		WeightsStore2[30] <= 19'd0;
		WeightsStore2[31] <= 19'd0;
		WeightsStore2[32] <= 19'd0;
		WeightsStore2[33] <= 19'd0;
		WeightsStore2[34] <= 19'd0;
		WeightsStore2[35] <= 19'd0;
		WeightsStore2[36] <= 19'd0;
		WeightsStore2[37] <= 19'd0;
		WeightsStore2[38] <= 19'd0;
		WeightsStore2[39] <= 19'd0;
		WeightsStore2[40] <= 19'd0;
		WeightsStore2[41] <= 19'd0;
		WeightsStore2[42] <= 19'd0;
		WeightsStore2[43] <= 19'd0;
		WeightsStore2[44] <= 19'd0;
		WeightsStore2[45] <= 19'd0;
		WeightsStore2[46] <= 19'd0;
		WeightsStore2[47] <= 19'd0;
		WeightsStore2[48] <= 19'd0;
		WeightsStore2[49] <= 19'd0;
		WeightsStore2[50] <= 19'd0;
		WeightsStore2[51] <= 19'd0;
		WeightsStore2[52] <= 19'd0;
		WeightsStore2[53] <= 19'd0;
		WeightsStore2[54] <= 19'd0;
		WeightsStore2[55] <= 19'd0;
		WeightsStore2[56] <= 19'd0;
		WeightsStore2[57] <= 19'd0;
		WeightsStore2[58] <= 19'd0;
		WeightsStore2[59] <= 19'd0;
		WeightsStore2[60] <= 19'd0;
		WeightsStore2[61] <= 19'd0;
		WeightsStore2[62] <= 19'd0;
		WeightsStore2[63] <= 19'd0;
		WeightsStore2[64] <= 19'd0;
		WeightsStore2[65] <= 19'd0;
		WeightsStore2[66] <= 19'd0;
		WeightsStore2[67] <= 19'd0;
		WeightsStore2[68] <= 19'd0;
		WeightsStore2[69] <= 19'd0;
		WeightsStore2[70] <= 19'd0;
		WeightsStore2[71] <= 19'd0;
		WeightsStore2[72] <= 19'd0;
		WeightsStore2[73] <= 19'd0;
		WeightsStore2[74] <= 19'd0;
		WeightsStore2[75] <= 19'd0;
		WeightsStore2[76] <= 19'd0;
		WeightsStore2[77] <= 19'd0;
		WeightsStore2[78] <= 19'd0;
		WeightsStore2[79] <= 19'd0;
		WeightsStore2[80] <= 19'd0;
		WeightsStore2[81] <= 19'd0;
		WeightsStore2[82] <= 19'd0;
		WeightsStore2[83] <= 19'd0;
		WeightsStore2[84] <= 19'd0;
		WeightsStore2[85] <= 19'd0;
		WeightsStore2[86] <= 19'd0;
		WeightsStore2[87] <= 19'd0;
		WeightsStore2[88] <= 19'd0;
		WeightsStore2[89] <= 19'd0;
		WeightsStore2[90] <= 19'd0;
		WeightsStore2[91] <= 19'd0;
		WeightsStore2[92] <= 19'd0;
		WeightsStore2[93] <= 19'd0;
		WeightsStore2[94] <= 19'd0;
		WeightsStore2[95] <= 19'd0;
		WeightsStore2[96] <= 19'd0;
		WeightsStore2[97] <= 19'd0;
		WeightsStore2[98] <= 19'd0;
		WeightsStore2[99] <= 19'd0;
		WeightsStore2[100] <= 19'd0;
		WeightsStore2[101] <= 19'd0;
		WeightsStore2[102] <= 19'd0;
		WeightsStore2[103] <= 19'd0;
		WeightsStore2[104] <= 19'd0;
		WeightsStore2[105] <= 19'd0;
		WeightsStore2[106] <= 19'd0;
		WeightsStore2[107] <= 19'd0;
		WeightsStore2[108] <= 19'd0;
		WeightsStore2[109] <= 19'd0;
		WeightsStore2[110] <= 19'd0;
		WeightsStore2[111] <= 19'd0;
		WeightsStore2[112] <= 19'd0;
		WeightsStore2[113] <= 19'd0;
		WeightsStore2[114] <= 19'd0;
		WeightsStore2[115] <= 19'd0;
		WeightsStore2[116] <= 19'd0;
		WeightsStore2[117] <= 19'd0;
		WeightsStore2[118] <= 19'd0;
		WeightsStore2[119] <= 19'd0;
		WeightsStore2[120] <= 19'd0;
		WeightsStore2[121] <= 19'd0;
		WeightsStore2[122] <= 19'd0;
		WeightsStore2[123] <= 19'd0;
		WeightsStore2[124] <= 19'd0;
		WeightsStore2[125] <= 19'd0;
		WeightsStore2[126] <= 19'd0;
		WeightsStore2[127] <= 19'd0;
		WeightsStore2[128] <= 19'd0;
		WeightsStore2[129] <= 19'd0;
		WeightsStore2[130] <= 19'd0;
		WeightsStore2[131] <= 19'd0;
		WeightsStore2[132] <= 19'd0;
		WeightsStore2[133] <= 19'd0;
		WeightsStore2[134] <= 19'd0;
		WeightsStore2[135] <= 19'd0;
		WeightsStore2[136] <= 19'd0;
		WeightsStore2[137] <= 19'd0;
		WeightsStore2[138] <= 19'd0;
		WeightsStore2[139] <= 19'd0;
		WeightsStore2[140] <= 19'd0;
		WeightsStore2[141] <= 19'd0;
		WeightsStore2[142] <= 19'd0;
		WeightsStore2[143] <= 19'd0;
		WeightsStore2[144] <= 19'd0;
		WeightsStore2[145] <= 19'd0;
		WeightsStore2[146] <= 19'd0;
		WeightsStore2[147] <= 19'd0;
		WeightsStore2[148] <= 19'd0;
		WeightsStore2[149] <= 19'd0;
		WeightsStore2[150] <= 19'd0;
		WeightsStore2[151] <= 19'd0;
		WeightsStore2[152] <= 19'd0;
		WeightsStore2[153] <= 19'd0;
		WeightsStore2[154] <= 19'd0;
		WeightsStore2[155] <= 19'd0;
		WeightsStore2[156] <= 19'd0;
		WeightsStore2[157] <= 19'd0;
		WeightsStore2[158] <= 19'd0;
		WeightsStore2[159] <= 19'd0;
		WeightsStore2[160] <= 19'd0;
		WeightsStore2[161] <= 19'd0;
		WeightsStore2[162] <= 19'd0;
		WeightsStore2[163] <= 19'd0;
		WeightsStore2[164] <= 19'd0;
		WeightsStore2[165] <= 19'd0;
		WeightsStore2[166] <= 19'd0;
		WeightsStore2[167] <= 19'd0;
		WeightsStore2[168] <= 19'd0;
		WeightsStore2[169] <= 19'd0;
		WeightsStore2[170] <= 19'd0;
		WeightsStore2[171] <= 19'd0;
		WeightsStore2[172] <= 19'd0;
		WeightsStore2[173] <= 19'd0;
		WeightsStore2[174] <= 19'd0;
		WeightsStore2[175] <= 19'd0;
		WeightsStore2[176] <= 19'd0;
		WeightsStore2[177] <= 19'd0;
		WeightsStore2[178] <= 19'd0;
		WeightsStore2[179] <= 19'd0;
		WeightsStore2[180] <= 19'd0;
		WeightsStore2[181] <= 19'd0;
		WeightsStore2[182] <= 19'd0;
		WeightsStore2[183] <= 19'd0;
		WeightsStore2[184] <= 19'd0;
		WeightsStore2[185] <= 19'd0;
		WeightsStore2[186] <= 19'd0;
		WeightsStore2[187] <= 19'd0;
		WeightsStore2[188] <= 19'd0;
		WeightsStore2[189] <= 19'd0;
		WeightsStore2[190] <= 19'd0;
		WeightsStore2[191] <= 19'd0;
		WeightsStore2[192] <= 19'd0;
		WeightsStore2[193] <= 19'd0;
		WeightsStore2[194] <= 19'd0;
		WeightsStore2[195] <= 19'd0;
		WeightsStore2[196] <= 19'd0;
		WeightsStore2[197] <= 19'd0;
		WeightsStore2[198] <= 19'd0;
		WeightsStore2[199] <= 19'd0;
		WeightsStore2[200] <= 19'd0;
		WeightsStore2[201] <= 19'd0;
		WeightsStore2[202] <= 19'd0;
		WeightsStore2[203] <= 19'd0;
		WeightsStore2[204] <= 19'd0;
		WeightsStore2[205] <= 19'd0;
		WeightsStore2[206] <= 19'd0;
		WeightsStore2[207] <= 19'd0;
		WeightsStore2[208] <= 19'd0;
		WeightsStore2[209] <= 19'd0;
		WeightsStore2[210] <= 19'd0;
		WeightsStore2[211] <= 19'd0;
		WeightsStore2[212] <= 19'd0;
		WeightsStore2[213] <= 19'd0;
		WeightsStore2[214] <= 19'd0;
		WeightsStore2[215] <= 19'd0;
		WeightsStore2[216] <= 19'd0;
		WeightsStore2[217] <= 19'd0;
		WeightsStore2[218] <= 19'd0;
		WeightsStore2[219] <= 19'd0;
		WeightsStore2[220] <= 19'd0;
		WeightsStore2[221] <= 19'd0;
		WeightsStore2[222] <= 19'd0;
		WeightsStore2[223] <= 19'd0;
		WeightsStore2[224] <= 19'd0;
		WeightsStore2[225] <= 19'd0;
		WeightsStore2[226] <= 19'd0;
		WeightsStore2[227] <= 19'd0;
		WeightsStore2[228] <= 19'd0;
		WeightsStore2[229] <= 19'd0;
		WeightsStore2[230] <= 19'd0;
		WeightsStore2[231] <= 19'd0;
		WeightsStore2[232] <= 19'd0;
		WeightsStore2[233] <= 19'd0;
		WeightsStore2[234] <= 19'd0;
		WeightsStore2[235] <= 19'd0;
		WeightsStore2[236] <= 19'd0;
		WeightsStore2[237] <= 19'd0;
		WeightsStore2[238] <= 19'd0;
		WeightsStore2[239] <= 19'd0;
		WeightsStore2[240] <= 19'd0;
		WeightsStore2[241] <= 19'd0;
		WeightsStore2[242] <= 19'd0;
		WeightsStore2[243] <= 19'd0;
		WeightsStore2[244] <= 19'd0;
		WeightsStore2[245] <= 19'd0;
		WeightsStore2[246] <= 19'd0;
		WeightsStore2[247] <= 19'd0;
		WeightsStore2[248] <= 19'd0;
		WeightsStore2[249] <= 19'd0;
		WeightsStore2[250] <= 19'd0;
		WeightsStore2[251] <= 19'd0;
		WeightsStore2[252] <= 19'd0;
		WeightsStore2[253] <= 19'd0;
		WeightsStore2[254] <= 19'd0;
		WeightsStore2[255] <= 19'd0;
		WeightsStore2[256] <= 19'd0;
		WeightsStore2[257] <= 19'd0;
		WeightsStore2[258] <= 19'd0;
		WeightsStore2[259] <= 19'd0;
		WeightsStore2[260] <= 19'd0;
		WeightsStore2[261] <= 19'd0;
		WeightsStore2[262] <= 19'd0;
		WeightsStore2[263] <= 19'd0;
		WeightsStore2[264] <= 19'd0;
		WeightsStore2[265] <= 19'd0;
		WeightsStore2[266] <= 19'd0;
		WeightsStore2[267] <= 19'd0;
		WeightsStore2[268] <= 19'd0;
		WeightsStore2[269] <= 19'd0;
		WeightsStore2[270] <= 19'd0;
		WeightsStore2[271] <= 19'd0;
		WeightsStore2[272] <= 19'd0;
		WeightsStore2[273] <= 19'd0;
		WeightsStore2[274] <= 19'd0;
		WeightsStore2[275] <= 19'd0;
		WeightsStore2[276] <= 19'd0;
		WeightsStore2[277] <= 19'd0;
		WeightsStore2[278] <= 19'd0;
		WeightsStore2[279] <= 19'd0;
		WeightsStore2[280] <= 19'd0;
		WeightsStore2[281] <= 19'd0;
		WeightsStore2[282] <= 19'd0;
		WeightsStore2[283] <= 19'd0;
		WeightsStore2[284] <= 19'd0;
		WeightsStore2[285] <= 19'd0;
		WeightsStore2[286] <= 19'd0;
		WeightsStore2[287] <= 19'd0;
		WeightsStore2[288] <= 19'd0;
		WeightsStore2[289] <= 19'd0;
		WeightsStore2[290] <= 19'd0;
		WeightsStore2[291] <= 19'd0;
		WeightsStore2[292] <= 19'd0;
		WeightsStore2[293] <= 19'd0;
		WeightsStore2[294] <= 19'd0;
		WeightsStore2[295] <= 19'd0;
		WeightsStore2[296] <= 19'd0;
		WeightsStore2[297] <= 19'd0;
		WeightsStore2[298] <= 19'd0;
		WeightsStore2[299] <= 19'd0;
		WeightsStore2[300] <= 19'd0;
		WeightsStore2[301] <= 19'd0;
		WeightsStore2[302] <= 19'd0;
		WeightsStore2[303] <= 19'd0;
		WeightsStore2[304] <= 19'd0;
		WeightsStore2[305] <= 19'd0;
		WeightsStore2[306] <= 19'd0;
		WeightsStore2[307] <= 19'd0;
		WeightsStore2[308] <= 19'd0;
		WeightsStore2[309] <= 19'd0;
		WeightsStore2[310] <= 19'd0;
		WeightsStore2[311] <= 19'd0;
		WeightsStore2[312] <= 19'd0;
		WeightsStore2[313] <= 19'd0;
		WeightsStore2[314] <= 19'd0;
		WeightsStore2[315] <= 19'd0;
		WeightsStore2[316] <= 19'd0;
		WeightsStore2[317] <= 19'd0;
		WeightsStore2[318] <= 19'd0;
		WeightsStore2[319] <= 19'd0;
		WeightsStore2[320] <= 19'd0;
		WeightsStore2[321] <= 19'd0;
		WeightsStore2[322] <= 19'd0;
		WeightsStore2[323] <= 19'd0;
		WeightsStore2[324] <= 19'd0;
		WeightsStore2[325] <= 19'd0;
		WeightsStore2[326] <= 19'd0;
		WeightsStore2[327] <= 19'd0;
		WeightsStore2[328] <= 19'd0;
		WeightsStore2[329] <= 19'd0;
		WeightsStore2[330] <= 19'd0;
		WeightsStore2[331] <= 19'd0;
		WeightsStore2[332] <= 19'd0;
		WeightsStore2[333] <= 19'd0;
		WeightsStore2[334] <= 19'd0;
		WeightsStore2[335] <= 19'd0;
		WeightsStore2[336] <= 19'd0;
		WeightsStore2[337] <= 19'd0;
		WeightsStore2[338] <= 19'd0;
		WeightsStore2[339] <= 19'd0;
		WeightsStore2[340] <= 19'd0;
		WeightsStore2[341] <= 19'd0;
		WeightsStore2[342] <= 19'd0;
		WeightsStore2[343] <= 19'd0;
		WeightsStore2[344] <= 19'd0;
		WeightsStore2[345] <= 19'd0;
		WeightsStore2[346] <= 19'd0;
		WeightsStore2[347] <= 19'd0;
		WeightsStore2[348] <= 19'd0;
		WeightsStore2[349] <= 19'd0;
		WeightsStore2[350] <= 19'd0;
		WeightsStore2[351] <= 19'd0;
		WeightsStore2[352] <= 19'd0;
		WeightsStore2[353] <= 19'd0;
		WeightsStore2[354] <= 19'd0;
		WeightsStore2[355] <= 19'd0;
		WeightsStore2[356] <= 19'd0;
		WeightsStore2[357] <= 19'd0;
		WeightsStore2[358] <= 19'd0;
		WeightsStore2[359] <= 19'd0;
		WeightsStore2[360] <= 19'd0;
		WeightsStore2[361] <= 19'd0;
		WeightsStore2[362] <= 19'd0;
		WeightsStore2[363] <= 19'd0;
		WeightsStore2[364] <= 19'd0;
		WeightsStore2[365] <= 19'd0;
		WeightsStore2[366] <= 19'd0;
		WeightsStore2[367] <= 19'd0;
		WeightsStore2[368] <= 19'd0;
		WeightsStore2[369] <= 19'd0;
		WeightsStore2[370] <= 19'd0;
		WeightsStore2[371] <= 19'd0;
		WeightsStore2[372] <= 19'd0;
		WeightsStore2[373] <= 19'd0;
		WeightsStore2[374] <= 19'd0;
		WeightsStore2[375] <= 19'd0;
		WeightsStore2[376] <= 19'd0;
		WeightsStore2[377] <= 19'd0;
		WeightsStore2[378] <= 19'd0;
		WeightsStore2[379] <= 19'd0;
		WeightsStore2[380] <= 19'd0;
		WeightsStore2[381] <= 19'd0;
		WeightsStore2[382] <= 19'd0;
		WeightsStore2[383] <= 19'd0;
		WeightsStore2[384] <= 19'd0;
		WeightsStore2[385] <= 19'd0;
		WeightsStore2[386] <= 19'd0;
		WeightsStore2[387] <= 19'd0;
		WeightsStore2[388] <= 19'd0;
		WeightsStore2[389] <= 19'd0;
		WeightsStore2[390] <= 19'd0;
		WeightsStore2[391] <= 19'd0;
		WeightsStore2[392] <= 19'd0;
		WeightsStore2[393] <= 19'd0;
		WeightsStore2[394] <= 19'd0;
		WeightsStore2[395] <= 19'd0;
		WeightsStore2[396] <= 19'd0;
		WeightsStore2[397] <= 19'd0;
		WeightsStore2[398] <= 19'd0;
		WeightsStore2[399] <= 19'd0;
		WeightsStore2[400] <= 19'd0;
		WeightsStore2[401] <= 19'd0;
		WeightsStore2[402] <= 19'd0;
		WeightsStore2[403] <= 19'd0;
		WeightsStore2[404] <= 19'd0;
		WeightsStore2[405] <= 19'd0;
		WeightsStore2[406] <= 19'd0;
		WeightsStore2[407] <= 19'd0;
		WeightsStore2[408] <= 19'd0;
		WeightsStore2[409] <= 19'd0;
		WeightsStore2[410] <= 19'd0;
		WeightsStore2[411] <= 19'd0;
		WeightsStore2[412] <= 19'd0;
		WeightsStore2[413] <= 19'd0;
		WeightsStore2[414] <= 19'd0;
		WeightsStore2[415] <= 19'd0;
		WeightsStore2[416] <= 19'd0;
		WeightsStore2[417] <= 19'd0;
		WeightsStore2[418] <= 19'd0;
		WeightsStore2[419] <= 19'd0;
		WeightsStore2[420] <= 19'd0;
		WeightsStore2[421] <= 19'd0;
		WeightsStore2[422] <= 19'd0;
		WeightsStore2[423] <= 19'd0;
		WeightsStore2[424] <= 19'd0;
		WeightsStore2[425] <= 19'd0;
		WeightsStore2[426] <= 19'd0;
		WeightsStore2[427] <= 19'd0;
		WeightsStore2[428] <= 19'd0;
		WeightsStore2[429] <= 19'd0;
		WeightsStore2[430] <= 19'd0;
		WeightsStore2[431] <= 19'd0;
		WeightsStore2[432] <= 19'd0;
		WeightsStore2[433] <= 19'd0;
		WeightsStore2[434] <= 19'd0;
		WeightsStore2[435] <= 19'd0;
		WeightsStore2[436] <= 19'd0;
		WeightsStore2[437] <= 19'd0;
		WeightsStore2[438] <= 19'd0;
		WeightsStore2[439] <= 19'd0;
		WeightsStore2[440] <= 19'd0;
		WeightsStore2[441] <= 19'd0;
		WeightsStore2[442] <= 19'd0;
		WeightsStore2[443] <= 19'd0;
		WeightsStore2[444] <= 19'd0;
		WeightsStore2[445] <= 19'd0;
		WeightsStore2[446] <= 19'd0;
		WeightsStore2[447] <= 19'd0;
		WeightsStore2[448] <= 19'd0;
		WeightsStore2[449] <= 19'd0;
		WeightsStore2[450] <= 19'd0;
		WeightsStore2[451] <= 19'd0;
		WeightsStore2[452] <= 19'd0;
		WeightsStore2[453] <= 19'd0;
		WeightsStore2[454] <= 19'd0;
		WeightsStore2[455] <= 19'd0;
		WeightsStore2[456] <= 19'd0;
		WeightsStore2[457] <= 19'd0;
		WeightsStore2[458] <= 19'd0;
		WeightsStore2[459] <= 19'd0;
		WeightsStore2[460] <= 19'd0;
		WeightsStore2[461] <= 19'd0;
		WeightsStore2[462] <= 19'd0;
		WeightsStore2[463] <= 19'd0;
		WeightsStore2[464] <= 19'd0;
		WeightsStore2[465] <= 19'd0;
		WeightsStore2[466] <= 19'd0;
		WeightsStore2[467] <= 19'd0;
		WeightsStore2[468] <= 19'd0;
		WeightsStore2[469] <= 19'd0;
		WeightsStore2[470] <= 19'd0;
		WeightsStore2[471] <= 19'd0;
		WeightsStore2[472] <= 19'd0;
		WeightsStore2[473] <= 19'd0;
		WeightsStore2[474] <= 19'd0;
		WeightsStore2[475] <= 19'd0;
		WeightsStore2[476] <= 19'd0;
		WeightsStore2[477] <= 19'd0;
		WeightsStore2[478] <= 19'd0;
		WeightsStore2[479] <= 19'd0;
		WeightsStore2[480] <= 19'd0;
		WeightsStore2[481] <= 19'd0;
		WeightsStore2[482] <= 19'd0;
		WeightsStore2[483] <= 19'd0;
		WeightsStore2[484] <= 19'd0;
		WeightsStore2[485] <= 19'd0;
		WeightsStore2[486] <= 19'd0;
		WeightsStore2[487] <= 19'd0;
		WeightsStore2[488] <= 19'd0;
		WeightsStore2[489] <= 19'd0;
		WeightsStore2[490] <= 19'd0;
		WeightsStore2[491] <= 19'd0;
		WeightsStore2[492] <= 19'd0;
		WeightsStore2[493] <= 19'd0;
		WeightsStore2[494] <= 19'd0;
		WeightsStore2[495] <= 19'd0;
		WeightsStore2[496] <= 19'd0;
		WeightsStore2[497] <= 19'd0;
		WeightsStore2[498] <= 19'd0;
		WeightsStore2[499] <= 19'd0;
		WeightsStore2[500] <= 19'd0;
		WeightsStore2[501] <= 19'd0;
		WeightsStore2[502] <= 19'd0;
		WeightsStore2[503] <= 19'd0;
		WeightsStore2[504] <= 19'd0;
		WeightsStore2[505] <= 19'd0;
		WeightsStore2[506] <= 19'd0;
		WeightsStore2[507] <= 19'd0;
		WeightsStore2[508] <= 19'd0;
		WeightsStore2[509] <= 19'd0;
		WeightsStore2[510] <= 19'd0;
		WeightsStore2[511] <= 19'd0;
		WeightsStore2[512] <= 19'd0;
		WeightsStore2[513] <= 19'd0;
		WeightsStore2[514] <= 19'd0;
		WeightsStore2[515] <= 19'd0;
		WeightsStore2[516] <= 19'd0;
		WeightsStore2[517] <= 19'd0;
		WeightsStore2[518] <= 19'd0;
		WeightsStore2[519] <= 19'd0;
		WeightsStore2[520] <= 19'd0;
		WeightsStore2[521] <= 19'd0;
		WeightsStore2[522] <= 19'd0;
		WeightsStore2[523] <= 19'd0;
		WeightsStore2[524] <= 19'd0;
		WeightsStore2[525] <= 19'd0;
		WeightsStore2[526] <= 19'd0;
		WeightsStore2[527] <= 19'd0;
		WeightsStore2[528] <= 19'd0;
		WeightsStore2[529] <= 19'd0;
		WeightsStore2[530] <= 19'd0;
		WeightsStore2[531] <= 19'd0;
		WeightsStore2[532] <= 19'd0;
		WeightsStore2[533] <= 19'd0;
		WeightsStore2[534] <= 19'd0;
		WeightsStore2[535] <= 19'd0;
		WeightsStore2[536] <= 19'd0;
		WeightsStore2[537] <= 19'd0;
		WeightsStore2[538] <= 19'd0;
		WeightsStore2[539] <= 19'd0;
		WeightsStore2[540] <= 19'd0;
		WeightsStore2[541] <= 19'd0;
		WeightsStore2[542] <= 19'd0;
		WeightsStore2[543] <= 19'd0;
		WeightsStore2[544] <= 19'd0;
		WeightsStore2[545] <= 19'd0;
		WeightsStore2[546] <= 19'd0;
		WeightsStore2[547] <= 19'd0;
		WeightsStore2[548] <= 19'd0;
		WeightsStore2[549] <= 19'd0;
		WeightsStore2[550] <= 19'd0;
		WeightsStore2[551] <= 19'd0;
		WeightsStore2[552] <= 19'd0;
		WeightsStore2[553] <= 19'd0;
		WeightsStore2[554] <= 19'd0;
		WeightsStore2[555] <= 19'd0;
		WeightsStore2[556] <= 19'd0;
		WeightsStore2[557] <= 19'd0;
		WeightsStore2[558] <= 19'd0;
		WeightsStore2[559] <= 19'd0;
		WeightsStore2[560] <= 19'd0;
		WeightsStore2[561] <= 19'd0;
		WeightsStore2[562] <= 19'd0;
		WeightsStore2[563] <= 19'd0;
		WeightsStore2[564] <= 19'd0;
		WeightsStore2[565] <= 19'd0;
		WeightsStore2[566] <= 19'd0;
		WeightsStore2[567] <= 19'd0;
		WeightsStore2[568] <= 19'd0;
		WeightsStore2[569] <= 19'd0;
		WeightsStore2[570] <= 19'd0;
		WeightsStore2[571] <= 19'd0;
		WeightsStore2[572] <= 19'd0;
		WeightsStore2[573] <= 19'd0;
		WeightsStore2[574] <= 19'd0;
		WeightsStore2[575] <= 19'd0;
		WeightsStore2[576] <= 19'd0;
		WeightsStore2[577] <= 19'd0;
		WeightsStore2[578] <= 19'd0;
		WeightsStore2[579] <= 19'd0;
		WeightsStore2[580] <= 19'd0;
		WeightsStore2[581] <= 19'd0;
		WeightsStore2[582] <= 19'd0;
		WeightsStore2[583] <= 19'd0;
		WeightsStore2[584] <= 19'd0;
		WeightsStore2[585] <= 19'd0;
		WeightsStore2[586] <= 19'd0;
		WeightsStore2[587] <= 19'd0;
		WeightsStore2[588] <= 19'd0;
		WeightsStore2[589] <= 19'd0;
		WeightsStore2[590] <= 19'd0;
		WeightsStore2[591] <= 19'd0;
		WeightsStore2[592] <= 19'd0;
		WeightsStore2[593] <= 19'd0;
		WeightsStore2[594] <= 19'd0;
		WeightsStore2[595] <= 19'd0;
		WeightsStore2[596] <= 19'd0;
		WeightsStore2[597] <= 19'd0;
		WeightsStore2[598] <= 19'd0;
		WeightsStore2[599] <= 19'd0;
		WeightsStore2[600] <= 19'd0;
		WeightsStore2[601] <= 19'd0;
		WeightsStore2[602] <= 19'd0;
		WeightsStore2[603] <= 19'd0;
		WeightsStore2[604] <= 19'd0;
		WeightsStore2[605] <= 19'd0;
		WeightsStore2[606] <= 19'd0;
		WeightsStore2[607] <= 19'd0;
		WeightsStore2[608] <= 19'd0;
		WeightsStore2[609] <= 19'd0;
		WeightsStore2[610] <= 19'd0;
		WeightsStore2[611] <= 19'd0;
		WeightsStore2[612] <= 19'd0;
		WeightsStore2[613] <= 19'd0;
		WeightsStore2[614] <= 19'd0;
		WeightsStore2[615] <= 19'd0;
		WeightsStore2[616] <= 19'd0;
		WeightsStore2[617] <= 19'd0;
		WeightsStore2[618] <= 19'd0;
		WeightsStore2[619] <= 19'd0;
		WeightsStore2[620] <= 19'd0;
		WeightsStore2[621] <= 19'd0;
		WeightsStore2[622] <= 19'd0;
		WeightsStore2[623] <= 19'd0;
		WeightsStore2[624] <= 19'd0;
		WeightsStore2[625] <= 19'd0;
		WeightsStore2[626] <= 19'd0;
		WeightsStore2[627] <= 19'd0;
		WeightsStore2[628] <= 19'd0;
		WeightsStore2[629] <= 19'd0;
		WeightsStore2[630] <= 19'd0;
		WeightsStore2[631] <= 19'd0;
		WeightsStore2[632] <= 19'd0;
		WeightsStore2[633] <= 19'd0;
		WeightsStore2[634] <= 19'd0;
		WeightsStore2[635] <= 19'd0;
		WeightsStore2[636] <= 19'd0;
		WeightsStore2[637] <= 19'd0;
		WeightsStore2[638] <= 19'd0;
		WeightsStore2[639] <= 19'd0;
		WeightsStore2[640] <= 19'd0;
		WeightsStore2[641] <= 19'd0;
		WeightsStore2[642] <= 19'd0;
		WeightsStore2[643] <= 19'd0;
		WeightsStore2[644] <= 19'd0;
		WeightsStore2[645] <= 19'd0;
		WeightsStore2[646] <= 19'd0;
		WeightsStore2[647] <= 19'd0;
		WeightsStore2[648] <= 19'd0;
		WeightsStore2[649] <= 19'd0;
		WeightsStore2[650] <= 19'd0;
		WeightsStore2[651] <= 19'd0;
		WeightsStore2[652] <= 19'd0;
		WeightsStore2[653] <= 19'd0;
		WeightsStore2[654] <= 19'd0;
		WeightsStore2[655] <= 19'd0;
		WeightsStore2[656] <= 19'd0;
		WeightsStore2[657] <= 19'd0;
		WeightsStore2[658] <= 19'd0;
		WeightsStore2[659] <= 19'd0;
		WeightsStore2[660] <= 19'd0;
		WeightsStore2[661] <= 19'd0;
		WeightsStore2[662] <= 19'd0;
		WeightsStore2[663] <= 19'd0;
		WeightsStore2[664] <= 19'd0;
		WeightsStore2[665] <= 19'd0;
		WeightsStore2[666] <= 19'd0;
		WeightsStore2[667] <= 19'd0;
		WeightsStore2[668] <= 19'd0;
		WeightsStore2[669] <= 19'd0;
		WeightsStore2[670] <= 19'd0;
		WeightsStore2[671] <= 19'd0;
		WeightsStore2[672] <= 19'd0;
		WeightsStore2[673] <= 19'd0;
		WeightsStore2[674] <= 19'd0;
		WeightsStore2[675] <= 19'd0;
		WeightsStore2[676] <= 19'd0;
		WeightsStore2[677] <= 19'd0;
		WeightsStore2[678] <= 19'd0;
		WeightsStore2[679] <= 19'd0;
		WeightsStore2[680] <= 19'd0;
		WeightsStore2[681] <= 19'd0;
		WeightsStore2[682] <= 19'd0;
		WeightsStore2[683] <= 19'd0;
		WeightsStore2[684] <= 19'd0;
		WeightsStore2[685] <= 19'd0;
		WeightsStore2[686] <= 19'd0;
		WeightsStore2[687] <= 19'd0;
		WeightsStore2[688] <= 19'd0;
		WeightsStore2[689] <= 19'd0;
		WeightsStore2[690] <= 19'd0;
		WeightsStore2[691] <= 19'd0;
		WeightsStore2[692] <= 19'd0;
		WeightsStore2[693] <= 19'd0;
		WeightsStore2[694] <= 19'd0;
		WeightsStore2[695] <= 19'd0;
		WeightsStore2[696] <= 19'd0;
		WeightsStore2[697] <= 19'd0;
		WeightsStore2[698] <= 19'd0;
		WeightsStore2[699] <= 19'd0;
		WeightsStore2[700] <= 19'd0;
		WeightsStore2[701] <= 19'd0;
		WeightsStore2[702] <= 19'd0;
		WeightsStore2[703] <= 19'd0;
		WeightsStore2[704] <= 19'd0;
		WeightsStore2[705] <= 19'd0;
		WeightsStore2[706] <= 19'd0;
		WeightsStore2[707] <= 19'd0;
		WeightsStore2[708] <= 19'd0;
		WeightsStore2[709] <= 19'd0;
		WeightsStore2[710] <= 19'd0;
		WeightsStore2[711] <= 19'd0;
		WeightsStore2[712] <= 19'd0;
		WeightsStore2[713] <= 19'd0;
		WeightsStore2[714] <= 19'd0;
		WeightsStore2[715] <= 19'd0;
		WeightsStore2[716] <= 19'd0;
		WeightsStore2[717] <= 19'd0;
		WeightsStore2[718] <= 19'd0;
		WeightsStore2[719] <= 19'd0;
		WeightsStore2[720] <= 19'd0;
		WeightsStore2[721] <= 19'd0;
		WeightsStore2[722] <= 19'd0;
		WeightsStore2[723] <= 19'd0;
		WeightsStore2[724] <= 19'd0;
		WeightsStore2[725] <= 19'd0;
		WeightsStore2[726] <= 19'd0;
		WeightsStore2[727] <= 19'd0;
		WeightsStore2[728] <= 19'd0;
		WeightsStore2[729] <= 19'd0;
		WeightsStore2[730] <= 19'd0;
		WeightsStore2[731] <= 19'd0;
		WeightsStore2[732] <= 19'd0;
		WeightsStore2[733] <= 19'd0;
		WeightsStore2[734] <= 19'd0;
		WeightsStore2[735] <= 19'd0;
		WeightsStore2[736] <= 19'd0;
		WeightsStore2[737] <= 19'd0;
		WeightsStore2[738] <= 19'd0;
		WeightsStore2[739] <= 19'd0;
		WeightsStore2[740] <= 19'd0;
		WeightsStore2[741] <= 19'd0;
		WeightsStore2[742] <= 19'd0;
		WeightsStore2[743] <= 19'd0;
		WeightsStore2[744] <= 19'd0;
		WeightsStore2[745] <= 19'd0;
		WeightsStore2[746] <= 19'd0;
		WeightsStore2[747] <= 19'd0;
		WeightsStore2[748] <= 19'd0;
		WeightsStore2[749] <= 19'd0;
		WeightsStore2[750] <= 19'd0;
		WeightsStore2[751] <= 19'd0;
		WeightsStore2[752] <= 19'd0;
		WeightsStore2[753] <= 19'd0;
		WeightsStore2[754] <= 19'd0;
		WeightsStore2[755] <= 19'd0;
		WeightsStore2[756] <= 19'd0;
		WeightsStore2[757] <= 19'd0;
		WeightsStore2[758] <= 19'd0;
		WeightsStore2[759] <= 19'd0;
		WeightsStore2[760] <= 19'd0;
		WeightsStore2[761] <= 19'd0;
		WeightsStore2[762] <= 19'd0;
		WeightsStore2[763] <= 19'd0;
		WeightsStore2[764] <= 19'd0;
		WeightsStore2[765] <= 19'd0;
		WeightsStore2[766] <= 19'd0;
		WeightsStore2[767] <= 19'd0;
		WeightsStore2[768] <= 19'd0;
		WeightsStore2[769] <= 19'd0;
		WeightsStore2[770] <= 19'd0;
		WeightsStore2[771] <= 19'd0;
		WeightsStore2[772] <= 19'd0;
		WeightsStore2[773] <= 19'd0;
		WeightsStore2[774] <= 19'd0;
		WeightsStore2[775] <= 19'd0;
		WeightsStore2[776] <= 19'd0;
		WeightsStore2[777] <= 19'd0;
		WeightsStore2[778] <= 19'd0;
		WeightsStore2[779] <= 19'd0;
		WeightsStore2[780] <= 19'd0;
		WeightsStore2[781] <= 19'd0;
		WeightsStore2[782] <= 19'd0;
		WeightsStore2[783] <= 19'd0;
		WeightsStore2[784] <= 19'd0;
		WeightsStore3[0] <= 19'd0;
		WeightsStore3[1] <= 19'd0;
		WeightsStore3[2] <= 19'd0;
		WeightsStore3[3] <= 19'd0;
		WeightsStore3[4] <= 19'd0;
		WeightsStore3[5] <= 19'd0;
		WeightsStore3[6] <= 19'd0;
		WeightsStore3[7] <= 19'd0;
		WeightsStore3[8] <= 19'd0;
		WeightsStore3[9] <= 19'd0;
		WeightsStore3[10] <= 19'd0;
		WeightsStore3[11] <= 19'd0;
		WeightsStore3[12] <= 19'd0;
		WeightsStore3[13] <= 19'd0;
		WeightsStore3[14] <= 19'd0;
		WeightsStore3[15] <= 19'd0;
		WeightsStore3[16] <= 19'd0;
		WeightsStore3[17] <= 19'd0;
		WeightsStore3[18] <= 19'd0;
		WeightsStore3[19] <= 19'd0;
		WeightsStore3[20] <= 19'd0;
		WeightsStore3[21] <= 19'd0;
		WeightsStore3[22] <= 19'd0;
		WeightsStore3[23] <= 19'd0;
		WeightsStore3[24] <= 19'd0;
		WeightsStore3[25] <= 19'd0;
		WeightsStore3[26] <= 19'd0;
		WeightsStore3[27] <= 19'd0;
		WeightsStore3[28] <= 19'd0;
		WeightsStore3[29] <= 19'd0;
		WeightsStore3[30] <= 19'd0;
		WeightsStore3[31] <= 19'd0;
		WeightsStore3[32] <= 19'd0;
		WeightsStore3[33] <= 19'd0;
		WeightsStore3[34] <= 19'd0;
		WeightsStore3[35] <= 19'd0;
		WeightsStore3[36] <= 19'd0;
		WeightsStore3[37] <= 19'd0;
		WeightsStore3[38] <= 19'd0;
		WeightsStore3[39] <= 19'd0;
		WeightsStore3[40] <= 19'd0;
		WeightsStore3[41] <= 19'd0;
		WeightsStore3[42] <= 19'd0;
		WeightsStore3[43] <= 19'd0;
		WeightsStore3[44] <= 19'd0;
		WeightsStore3[45] <= 19'd0;
		WeightsStore3[46] <= 19'd0;
		WeightsStore3[47] <= 19'd0;
		WeightsStore3[48] <= 19'd0;
		WeightsStore3[49] <= 19'd0;
		WeightsStore3[50] <= 19'd0;
		WeightsStore3[51] <= 19'd0;
		WeightsStore3[52] <= 19'd0;
		WeightsStore3[53] <= 19'd0;
		WeightsStore3[54] <= 19'd0;
		WeightsStore3[55] <= 19'd0;
		WeightsStore3[56] <= 19'd0;
		WeightsStore3[57] <= 19'd0;
		WeightsStore3[58] <= 19'd0;
		WeightsStore3[59] <= 19'd0;
		WeightsStore3[60] <= 19'd0;
		WeightsStore3[61] <= 19'd0;
		WeightsStore3[62] <= 19'd0;
		WeightsStore3[63] <= 19'd0;
		WeightsStore3[64] <= 19'd0;
		WeightsStore3[65] <= 19'd0;
		WeightsStore3[66] <= 19'd0;
		WeightsStore3[67] <= 19'd0;
		WeightsStore3[68] <= 19'd0;
		WeightsStore3[69] <= 19'd0;
		WeightsStore3[70] <= 19'd0;
		WeightsStore3[71] <= 19'd0;
		WeightsStore3[72] <= 19'd0;
		WeightsStore3[73] <= 19'd0;
		WeightsStore3[74] <= 19'd0;
		WeightsStore3[75] <= 19'd0;
		WeightsStore3[76] <= 19'd0;
		WeightsStore3[77] <= 19'd0;
		WeightsStore3[78] <= 19'd0;
		WeightsStore3[79] <= 19'd0;
		WeightsStore3[80] <= 19'd0;
		WeightsStore3[81] <= 19'd0;
		WeightsStore3[82] <= 19'd0;
		WeightsStore3[83] <= 19'd0;
		WeightsStore3[84] <= 19'd0;
		WeightsStore3[85] <= 19'd0;
		WeightsStore3[86] <= 19'd0;
		WeightsStore3[87] <= 19'd0;
		WeightsStore3[88] <= 19'd0;
		WeightsStore3[89] <= 19'd0;
		WeightsStore3[90] <= 19'd0;
		WeightsStore3[91] <= 19'd0;
		WeightsStore3[92] <= 19'd0;
		WeightsStore3[93] <= 19'd0;
		WeightsStore3[94] <= 19'd0;
		WeightsStore3[95] <= 19'd0;
		WeightsStore3[96] <= 19'd0;
		WeightsStore3[97] <= 19'd0;
		WeightsStore3[98] <= 19'd0;
		WeightsStore3[99] <= 19'd0;
		WeightsStore3[100] <= 19'd0;
		WeightsStore3[101] <= 19'd0;
		WeightsStore3[102] <= 19'd0;
		WeightsStore3[103] <= 19'd0;
		WeightsStore3[104] <= 19'd0;
		WeightsStore3[105] <= 19'd0;
		WeightsStore3[106] <= 19'd0;
		WeightsStore3[107] <= 19'd0;
		WeightsStore3[108] <= 19'd0;
		WeightsStore3[109] <= 19'd0;
		WeightsStore3[110] <= 19'd0;
		WeightsStore3[111] <= 19'd0;
		WeightsStore3[112] <= 19'd0;
		WeightsStore3[113] <= 19'd0;
		WeightsStore3[114] <= 19'd0;
		WeightsStore3[115] <= 19'd0;
		WeightsStore3[116] <= 19'd0;
		WeightsStore3[117] <= 19'd0;
		WeightsStore3[118] <= 19'd0;
		WeightsStore3[119] <= 19'd0;
		WeightsStore3[120] <= 19'd0;
		WeightsStore3[121] <= 19'd0;
		WeightsStore3[122] <= 19'd0;
		WeightsStore3[123] <= 19'd0;
		WeightsStore3[124] <= 19'd0;
		WeightsStore3[125] <= 19'd0;
		WeightsStore3[126] <= 19'd0;
		WeightsStore3[127] <= 19'd0;
		WeightsStore3[128] <= 19'd0;
		WeightsStore3[129] <= 19'd0;
		WeightsStore3[130] <= 19'd0;
		WeightsStore3[131] <= 19'd0;
		WeightsStore3[132] <= 19'd0;
		WeightsStore3[133] <= 19'd0;
		WeightsStore3[134] <= 19'd0;
		WeightsStore3[135] <= 19'd0;
		WeightsStore3[136] <= 19'd0;
		WeightsStore3[137] <= 19'd0;
		WeightsStore3[138] <= 19'd0;
		WeightsStore3[139] <= 19'd0;
		WeightsStore3[140] <= 19'd0;
		WeightsStore3[141] <= 19'd0;
		WeightsStore3[142] <= 19'd0;
		WeightsStore3[143] <= 19'd0;
		WeightsStore3[144] <= 19'd0;
		WeightsStore3[145] <= 19'd0;
		WeightsStore3[146] <= 19'd0;
		WeightsStore3[147] <= 19'd0;
		WeightsStore3[148] <= 19'd0;
		WeightsStore3[149] <= 19'd0;
		WeightsStore3[150] <= 19'd0;
		WeightsStore3[151] <= 19'd0;
		WeightsStore3[152] <= 19'd0;
		WeightsStore3[153] <= 19'd0;
		WeightsStore3[154] <= 19'd0;
		WeightsStore3[155] <= 19'd0;
		WeightsStore3[156] <= 19'd0;
		WeightsStore3[157] <= 19'd0;
		WeightsStore3[158] <= 19'd0;
		WeightsStore3[159] <= 19'd0;
		WeightsStore3[160] <= 19'd0;
		WeightsStore3[161] <= 19'd0;
		WeightsStore3[162] <= 19'd0;
		WeightsStore3[163] <= 19'd0;
		WeightsStore3[164] <= 19'd0;
		WeightsStore3[165] <= 19'd0;
		WeightsStore3[166] <= 19'd0;
		WeightsStore3[167] <= 19'd0;
		WeightsStore3[168] <= 19'd0;
		WeightsStore3[169] <= 19'd0;
		WeightsStore3[170] <= 19'd0;
		WeightsStore3[171] <= 19'd0;
		WeightsStore3[172] <= 19'd0;
		WeightsStore3[173] <= 19'd0;
		WeightsStore3[174] <= 19'd0;
		WeightsStore3[175] <= 19'd0;
		WeightsStore3[176] <= 19'd0;
		WeightsStore3[177] <= 19'd0;
		WeightsStore3[178] <= 19'd0;
		WeightsStore3[179] <= 19'd0;
		WeightsStore3[180] <= 19'd0;
		WeightsStore3[181] <= 19'd0;
		WeightsStore3[182] <= 19'd0;
		WeightsStore3[183] <= 19'd0;
		WeightsStore3[184] <= 19'd0;
		WeightsStore3[185] <= 19'd0;
		WeightsStore3[186] <= 19'd0;
		WeightsStore3[187] <= 19'd0;
		WeightsStore3[188] <= 19'd0;
		WeightsStore3[189] <= 19'd0;
		WeightsStore3[190] <= 19'd0;
		WeightsStore3[191] <= 19'd0;
		WeightsStore3[192] <= 19'd0;
		WeightsStore3[193] <= 19'd0;
		WeightsStore3[194] <= 19'd0;
		WeightsStore3[195] <= 19'd0;
		WeightsStore3[196] <= 19'd0;
		WeightsStore3[197] <= 19'd0;
		WeightsStore3[198] <= 19'd0;
		WeightsStore3[199] <= 19'd0;
		WeightsStore3[200] <= 19'd0;
		WeightsStore3[201] <= 19'd0;
		WeightsStore3[202] <= 19'd0;
		WeightsStore3[203] <= 19'd0;
		WeightsStore3[204] <= 19'd0;
		WeightsStore3[205] <= 19'd0;
		WeightsStore3[206] <= 19'd0;
		WeightsStore3[207] <= 19'd0;
		WeightsStore3[208] <= 19'd0;
		WeightsStore3[209] <= 19'd0;
		WeightsStore3[210] <= 19'd0;
		WeightsStore3[211] <= 19'd0;
		WeightsStore3[212] <= 19'd0;
		WeightsStore3[213] <= 19'd0;
		WeightsStore3[214] <= 19'd0;
		WeightsStore3[215] <= 19'd0;
		WeightsStore3[216] <= 19'd0;
		WeightsStore3[217] <= 19'd0;
		WeightsStore3[218] <= 19'd0;
		WeightsStore3[219] <= 19'd0;
		WeightsStore3[220] <= 19'd0;
		WeightsStore3[221] <= 19'd0;
		WeightsStore3[222] <= 19'd0;
		WeightsStore3[223] <= 19'd0;
		WeightsStore3[224] <= 19'd0;
		WeightsStore3[225] <= 19'd0;
		WeightsStore3[226] <= 19'd0;
		WeightsStore3[227] <= 19'd0;
		WeightsStore3[228] <= 19'd0;
		WeightsStore3[229] <= 19'd0;
		WeightsStore3[230] <= 19'd0;
		WeightsStore3[231] <= 19'd0;
		WeightsStore3[232] <= 19'd0;
		WeightsStore3[233] <= 19'd0;
		WeightsStore3[234] <= 19'd0;
		WeightsStore3[235] <= 19'd0;
		WeightsStore3[236] <= 19'd0;
		WeightsStore3[237] <= 19'd0;
		WeightsStore3[238] <= 19'd0;
		WeightsStore3[239] <= 19'd0;
		WeightsStore3[240] <= 19'd0;
		WeightsStore3[241] <= 19'd0;
		WeightsStore3[242] <= 19'd0;
		WeightsStore3[243] <= 19'd0;
		WeightsStore3[244] <= 19'd0;
		WeightsStore3[245] <= 19'd0;
		WeightsStore3[246] <= 19'd0;
		WeightsStore3[247] <= 19'd0;
		WeightsStore3[248] <= 19'd0;
		WeightsStore3[249] <= 19'd0;
		WeightsStore3[250] <= 19'd0;
		WeightsStore3[251] <= 19'd0;
		WeightsStore3[252] <= 19'd0;
		WeightsStore3[253] <= 19'd0;
		WeightsStore3[254] <= 19'd0;
		WeightsStore3[255] <= 19'd0;
		WeightsStore3[256] <= 19'd0;
		WeightsStore3[257] <= 19'd0;
		WeightsStore3[258] <= 19'd0;
		WeightsStore3[259] <= 19'd0;
		WeightsStore3[260] <= 19'd0;
		WeightsStore3[261] <= 19'd0;
		WeightsStore3[262] <= 19'd0;
		WeightsStore3[263] <= 19'd0;
		WeightsStore3[264] <= 19'd0;
		WeightsStore3[265] <= 19'd0;
		WeightsStore3[266] <= 19'd0;
		WeightsStore3[267] <= 19'd0;
		WeightsStore3[268] <= 19'd0;
		WeightsStore3[269] <= 19'd0;
		WeightsStore3[270] <= 19'd0;
		WeightsStore3[271] <= 19'd0;
		WeightsStore3[272] <= 19'd0;
		WeightsStore3[273] <= 19'd0;
		WeightsStore3[274] <= 19'd0;
		WeightsStore3[275] <= 19'd0;
		WeightsStore3[276] <= 19'd0;
		WeightsStore3[277] <= 19'd0;
		WeightsStore3[278] <= 19'd0;
		WeightsStore3[279] <= 19'd0;
		WeightsStore3[280] <= 19'd0;
		WeightsStore3[281] <= 19'd0;
		WeightsStore3[282] <= 19'd0;
		WeightsStore3[283] <= 19'd0;
		WeightsStore3[284] <= 19'd0;
		WeightsStore3[285] <= 19'd0;
		WeightsStore3[286] <= 19'd0;
		WeightsStore3[287] <= 19'd0;
		WeightsStore3[288] <= 19'd0;
		WeightsStore3[289] <= 19'd0;
		WeightsStore3[290] <= 19'd0;
		WeightsStore3[291] <= 19'd0;
		WeightsStore3[292] <= 19'd0;
		WeightsStore3[293] <= 19'd0;
		WeightsStore3[294] <= 19'd0;
		WeightsStore3[295] <= 19'd0;
		WeightsStore3[296] <= 19'd0;
		WeightsStore3[297] <= 19'd0;
		WeightsStore3[298] <= 19'd0;
		WeightsStore3[299] <= 19'd0;
		WeightsStore3[300] <= 19'd0;
		WeightsStore3[301] <= 19'd0;
		WeightsStore3[302] <= 19'd0;
		WeightsStore3[303] <= 19'd0;
		WeightsStore3[304] <= 19'd0;
		WeightsStore3[305] <= 19'd0;
		WeightsStore3[306] <= 19'd0;
		WeightsStore3[307] <= 19'd0;
		WeightsStore3[308] <= 19'd0;
		WeightsStore3[309] <= 19'd0;
		WeightsStore3[310] <= 19'd0;
		WeightsStore3[311] <= 19'd0;
		WeightsStore3[312] <= 19'd0;
		WeightsStore3[313] <= 19'd0;
		WeightsStore3[314] <= 19'd0;
		WeightsStore3[315] <= 19'd0;
		WeightsStore3[316] <= 19'd0;
		WeightsStore3[317] <= 19'd0;
		WeightsStore3[318] <= 19'd0;
		WeightsStore3[319] <= 19'd0;
		WeightsStore3[320] <= 19'd0;
		WeightsStore3[321] <= 19'd0;
		WeightsStore3[322] <= 19'd0;
		WeightsStore3[323] <= 19'd0;
		WeightsStore3[324] <= 19'd0;
		WeightsStore3[325] <= 19'd0;
		WeightsStore3[326] <= 19'd0;
		WeightsStore3[327] <= 19'd0;
		WeightsStore3[328] <= 19'd0;
		WeightsStore3[329] <= 19'd0;
		WeightsStore3[330] <= 19'd0;
		WeightsStore3[331] <= 19'd0;
		WeightsStore3[332] <= 19'd0;
		WeightsStore3[333] <= 19'd0;
		WeightsStore3[334] <= 19'd0;
		WeightsStore3[335] <= 19'd0;
		WeightsStore3[336] <= 19'd0;
		WeightsStore3[337] <= 19'd0;
		WeightsStore3[338] <= 19'd0;
		WeightsStore3[339] <= 19'd0;
		WeightsStore3[340] <= 19'd0;
		WeightsStore3[341] <= 19'd0;
		WeightsStore3[342] <= 19'd0;
		WeightsStore3[343] <= 19'd0;
		WeightsStore3[344] <= 19'd0;
		WeightsStore3[345] <= 19'd0;
		WeightsStore3[346] <= 19'd0;
		WeightsStore3[347] <= 19'd0;
		WeightsStore3[348] <= 19'd0;
		WeightsStore3[349] <= 19'd0;
		WeightsStore3[350] <= 19'd0;
		WeightsStore3[351] <= 19'd0;
		WeightsStore3[352] <= 19'd0;
		WeightsStore3[353] <= 19'd0;
		WeightsStore3[354] <= 19'd0;
		WeightsStore3[355] <= 19'd0;
		WeightsStore3[356] <= 19'd0;
		WeightsStore3[357] <= 19'd0;
		WeightsStore3[358] <= 19'd0;
		WeightsStore3[359] <= 19'd0;
		WeightsStore3[360] <= 19'd0;
		WeightsStore3[361] <= 19'd0;
		WeightsStore3[362] <= 19'd0;
		WeightsStore3[363] <= 19'd0;
		WeightsStore3[364] <= 19'd0;
		WeightsStore3[365] <= 19'd0;
		WeightsStore3[366] <= 19'd0;
		WeightsStore3[367] <= 19'd0;
		WeightsStore3[368] <= 19'd0;
		WeightsStore3[369] <= 19'd0;
		WeightsStore3[370] <= 19'd0;
		WeightsStore3[371] <= 19'd0;
		WeightsStore3[372] <= 19'd0;
		WeightsStore3[373] <= 19'd0;
		WeightsStore3[374] <= 19'd0;
		WeightsStore3[375] <= 19'd0;
		WeightsStore3[376] <= 19'd0;
		WeightsStore3[377] <= 19'd0;
		WeightsStore3[378] <= 19'd0;
		WeightsStore3[379] <= 19'd0;
		WeightsStore3[380] <= 19'd0;
		WeightsStore3[381] <= 19'd0;
		WeightsStore3[382] <= 19'd0;
		WeightsStore3[383] <= 19'd0;
		WeightsStore3[384] <= 19'd0;
		WeightsStore3[385] <= 19'd0;
		WeightsStore3[386] <= 19'd0;
		WeightsStore3[387] <= 19'd0;
		WeightsStore3[388] <= 19'd0;
		WeightsStore3[389] <= 19'd0;
		WeightsStore3[390] <= 19'd0;
		WeightsStore3[391] <= 19'd0;
		WeightsStore3[392] <= 19'd0;
		WeightsStore3[393] <= 19'd0;
		WeightsStore3[394] <= 19'd0;
		WeightsStore3[395] <= 19'd0;
		WeightsStore3[396] <= 19'd0;
		WeightsStore3[397] <= 19'd0;
		WeightsStore3[398] <= 19'd0;
		WeightsStore3[399] <= 19'd0;
		WeightsStore3[400] <= 19'd0;
		WeightsStore3[401] <= 19'd0;
		WeightsStore3[402] <= 19'd0;
		WeightsStore3[403] <= 19'd0;
		WeightsStore3[404] <= 19'd0;
		WeightsStore3[405] <= 19'd0;
		WeightsStore3[406] <= 19'd0;
		WeightsStore3[407] <= 19'd0;
		WeightsStore3[408] <= 19'd0;
		WeightsStore3[409] <= 19'd0;
		WeightsStore3[410] <= 19'd0;
		WeightsStore3[411] <= 19'd0;
		WeightsStore3[412] <= 19'd0;
		WeightsStore3[413] <= 19'd0;
		WeightsStore3[414] <= 19'd0;
		WeightsStore3[415] <= 19'd0;
		WeightsStore3[416] <= 19'd0;
		WeightsStore3[417] <= 19'd0;
		WeightsStore3[418] <= 19'd0;
		WeightsStore3[419] <= 19'd0;
		WeightsStore3[420] <= 19'd0;
		WeightsStore3[421] <= 19'd0;
		WeightsStore3[422] <= 19'd0;
		WeightsStore3[423] <= 19'd0;
		WeightsStore3[424] <= 19'd0;
		WeightsStore3[425] <= 19'd0;
		WeightsStore3[426] <= 19'd0;
		WeightsStore3[427] <= 19'd0;
		WeightsStore3[428] <= 19'd0;
		WeightsStore3[429] <= 19'd0;
		WeightsStore3[430] <= 19'd0;
		WeightsStore3[431] <= 19'd0;
		WeightsStore3[432] <= 19'd0;
		WeightsStore3[433] <= 19'd0;
		WeightsStore3[434] <= 19'd0;
		WeightsStore3[435] <= 19'd0;
		WeightsStore3[436] <= 19'd0;
		WeightsStore3[437] <= 19'd0;
		WeightsStore3[438] <= 19'd0;
		WeightsStore3[439] <= 19'd0;
		WeightsStore3[440] <= 19'd0;
		WeightsStore3[441] <= 19'd0;
		WeightsStore3[442] <= 19'd0;
		WeightsStore3[443] <= 19'd0;
		WeightsStore3[444] <= 19'd0;
		WeightsStore3[445] <= 19'd0;
		WeightsStore3[446] <= 19'd0;
		WeightsStore3[447] <= 19'd0;
		WeightsStore3[448] <= 19'd0;
		WeightsStore3[449] <= 19'd0;
		WeightsStore3[450] <= 19'd0;
		WeightsStore3[451] <= 19'd0;
		WeightsStore3[452] <= 19'd0;
		WeightsStore3[453] <= 19'd0;
		WeightsStore3[454] <= 19'd0;
		WeightsStore3[455] <= 19'd0;
		WeightsStore3[456] <= 19'd0;
		WeightsStore3[457] <= 19'd0;
		WeightsStore3[458] <= 19'd0;
		WeightsStore3[459] <= 19'd0;
		WeightsStore3[460] <= 19'd0;
		WeightsStore3[461] <= 19'd0;
		WeightsStore3[462] <= 19'd0;
		WeightsStore3[463] <= 19'd0;
		WeightsStore3[464] <= 19'd0;
		WeightsStore3[465] <= 19'd0;
		WeightsStore3[466] <= 19'd0;
		WeightsStore3[467] <= 19'd0;
		WeightsStore3[468] <= 19'd0;
		WeightsStore3[469] <= 19'd0;
		WeightsStore3[470] <= 19'd0;
		WeightsStore3[471] <= 19'd0;
		WeightsStore3[472] <= 19'd0;
		WeightsStore3[473] <= 19'd0;
		WeightsStore3[474] <= 19'd0;
		WeightsStore3[475] <= 19'd0;
		WeightsStore3[476] <= 19'd0;
		WeightsStore3[477] <= 19'd0;
		WeightsStore3[478] <= 19'd0;
		WeightsStore3[479] <= 19'd0;
		WeightsStore3[480] <= 19'd0;
		WeightsStore3[481] <= 19'd0;
		WeightsStore3[482] <= 19'd0;
		WeightsStore3[483] <= 19'd0;
		WeightsStore3[484] <= 19'd0;
		WeightsStore3[485] <= 19'd0;
		WeightsStore3[486] <= 19'd0;
		WeightsStore3[487] <= 19'd0;
		WeightsStore3[488] <= 19'd0;
		WeightsStore3[489] <= 19'd0;
		WeightsStore3[490] <= 19'd0;
		WeightsStore3[491] <= 19'd0;
		WeightsStore3[492] <= 19'd0;
		WeightsStore3[493] <= 19'd0;
		WeightsStore3[494] <= 19'd0;
		WeightsStore3[495] <= 19'd0;
		WeightsStore3[496] <= 19'd0;
		WeightsStore3[497] <= 19'd0;
		WeightsStore3[498] <= 19'd0;
		WeightsStore3[499] <= 19'd0;
		WeightsStore3[500] <= 19'd0;
		WeightsStore3[501] <= 19'd0;
		WeightsStore3[502] <= 19'd0;
		WeightsStore3[503] <= 19'd0;
		WeightsStore3[504] <= 19'd0;
		WeightsStore3[505] <= 19'd0;
		WeightsStore3[506] <= 19'd0;
		WeightsStore3[507] <= 19'd0;
		WeightsStore3[508] <= 19'd0;
		WeightsStore3[509] <= 19'd0;
		WeightsStore3[510] <= 19'd0;
		WeightsStore3[511] <= 19'd0;
		WeightsStore3[512] <= 19'd0;
		WeightsStore3[513] <= 19'd0;
		WeightsStore3[514] <= 19'd0;
		WeightsStore3[515] <= 19'd0;
		WeightsStore3[516] <= 19'd0;
		WeightsStore3[517] <= 19'd0;
		WeightsStore3[518] <= 19'd0;
		WeightsStore3[519] <= 19'd0;
		WeightsStore3[520] <= 19'd0;
		WeightsStore3[521] <= 19'd0;
		WeightsStore3[522] <= 19'd0;
		WeightsStore3[523] <= 19'd0;
		WeightsStore3[524] <= 19'd0;
		WeightsStore3[525] <= 19'd0;
		WeightsStore3[526] <= 19'd0;
		WeightsStore3[527] <= 19'd0;
		WeightsStore3[528] <= 19'd0;
		WeightsStore3[529] <= 19'd0;
		WeightsStore3[530] <= 19'd0;
		WeightsStore3[531] <= 19'd0;
		WeightsStore3[532] <= 19'd0;
		WeightsStore3[533] <= 19'd0;
		WeightsStore3[534] <= 19'd0;
		WeightsStore3[535] <= 19'd0;
		WeightsStore3[536] <= 19'd0;
		WeightsStore3[537] <= 19'd0;
		WeightsStore3[538] <= 19'd0;
		WeightsStore3[539] <= 19'd0;
		WeightsStore3[540] <= 19'd0;
		WeightsStore3[541] <= 19'd0;
		WeightsStore3[542] <= 19'd0;
		WeightsStore3[543] <= 19'd0;
		WeightsStore3[544] <= 19'd0;
		WeightsStore3[545] <= 19'd0;
		WeightsStore3[546] <= 19'd0;
		WeightsStore3[547] <= 19'd0;
		WeightsStore3[548] <= 19'd0;
		WeightsStore3[549] <= 19'd0;
		WeightsStore3[550] <= 19'd0;
		WeightsStore3[551] <= 19'd0;
		WeightsStore3[552] <= 19'd0;
		WeightsStore3[553] <= 19'd0;
		WeightsStore3[554] <= 19'd0;
		WeightsStore3[555] <= 19'd0;
		WeightsStore3[556] <= 19'd0;
		WeightsStore3[557] <= 19'd0;
		WeightsStore3[558] <= 19'd0;
		WeightsStore3[559] <= 19'd0;
		WeightsStore3[560] <= 19'd0;
		WeightsStore3[561] <= 19'd0;
		WeightsStore3[562] <= 19'd0;
		WeightsStore3[563] <= 19'd0;
		WeightsStore3[564] <= 19'd0;
		WeightsStore3[565] <= 19'd0;
		WeightsStore3[566] <= 19'd0;
		WeightsStore3[567] <= 19'd0;
		WeightsStore3[568] <= 19'd0;
		WeightsStore3[569] <= 19'd0;
		WeightsStore3[570] <= 19'd0;
		WeightsStore3[571] <= 19'd0;
		WeightsStore3[572] <= 19'd0;
		WeightsStore3[573] <= 19'd0;
		WeightsStore3[574] <= 19'd0;
		WeightsStore3[575] <= 19'd0;
		WeightsStore3[576] <= 19'd0;
		WeightsStore3[577] <= 19'd0;
		WeightsStore3[578] <= 19'd0;
		WeightsStore3[579] <= 19'd0;
		WeightsStore3[580] <= 19'd0;
		WeightsStore3[581] <= 19'd0;
		WeightsStore3[582] <= 19'd0;
		WeightsStore3[583] <= 19'd0;
		WeightsStore3[584] <= 19'd0;
		WeightsStore3[585] <= 19'd0;
		WeightsStore3[586] <= 19'd0;
		WeightsStore3[587] <= 19'd0;
		WeightsStore3[588] <= 19'd0;
		WeightsStore3[589] <= 19'd0;
		WeightsStore3[590] <= 19'd0;
		WeightsStore3[591] <= 19'd0;
		WeightsStore3[592] <= 19'd0;
		WeightsStore3[593] <= 19'd0;
		WeightsStore3[594] <= 19'd0;
		WeightsStore3[595] <= 19'd0;
		WeightsStore3[596] <= 19'd0;
		WeightsStore3[597] <= 19'd0;
		WeightsStore3[598] <= 19'd0;
		WeightsStore3[599] <= 19'd0;
		WeightsStore3[600] <= 19'd0;
		WeightsStore3[601] <= 19'd0;
		WeightsStore3[602] <= 19'd0;
		WeightsStore3[603] <= 19'd0;
		WeightsStore3[604] <= 19'd0;
		WeightsStore3[605] <= 19'd0;
		WeightsStore3[606] <= 19'd0;
		WeightsStore3[607] <= 19'd0;
		WeightsStore3[608] <= 19'd0;
		WeightsStore3[609] <= 19'd0;
		WeightsStore3[610] <= 19'd0;
		WeightsStore3[611] <= 19'd0;
		WeightsStore3[612] <= 19'd0;
		WeightsStore3[613] <= 19'd0;
		WeightsStore3[614] <= 19'd0;
		WeightsStore3[615] <= 19'd0;
		WeightsStore3[616] <= 19'd0;
		WeightsStore3[617] <= 19'd0;
		WeightsStore3[618] <= 19'd0;
		WeightsStore3[619] <= 19'd0;
		WeightsStore3[620] <= 19'd0;
		WeightsStore3[621] <= 19'd0;
		WeightsStore3[622] <= 19'd0;
		WeightsStore3[623] <= 19'd0;
		WeightsStore3[624] <= 19'd0;
		WeightsStore3[625] <= 19'd0;
		WeightsStore3[626] <= 19'd0;
		WeightsStore3[627] <= 19'd0;
		WeightsStore3[628] <= 19'd0;
		WeightsStore3[629] <= 19'd0;
		WeightsStore3[630] <= 19'd0;
		WeightsStore3[631] <= 19'd0;
		WeightsStore3[632] <= 19'd0;
		WeightsStore3[633] <= 19'd0;
		WeightsStore3[634] <= 19'd0;
		WeightsStore3[635] <= 19'd0;
		WeightsStore3[636] <= 19'd0;
		WeightsStore3[637] <= 19'd0;
		WeightsStore3[638] <= 19'd0;
		WeightsStore3[639] <= 19'd0;
		WeightsStore3[640] <= 19'd0;
		WeightsStore3[641] <= 19'd0;
		WeightsStore3[642] <= 19'd0;
		WeightsStore3[643] <= 19'd0;
		WeightsStore3[644] <= 19'd0;
		WeightsStore3[645] <= 19'd0;
		WeightsStore3[646] <= 19'd0;
		WeightsStore3[647] <= 19'd0;
		WeightsStore3[648] <= 19'd0;
		WeightsStore3[649] <= 19'd0;
		WeightsStore3[650] <= 19'd0;
		WeightsStore3[651] <= 19'd0;
		WeightsStore3[652] <= 19'd0;
		WeightsStore3[653] <= 19'd0;
		WeightsStore3[654] <= 19'd0;
		WeightsStore3[655] <= 19'd0;
		WeightsStore3[656] <= 19'd0;
		WeightsStore3[657] <= 19'd0;
		WeightsStore3[658] <= 19'd0;
		WeightsStore3[659] <= 19'd0;
		WeightsStore3[660] <= 19'd0;
		WeightsStore3[661] <= 19'd0;
		WeightsStore3[662] <= 19'd0;
		WeightsStore3[663] <= 19'd0;
		WeightsStore3[664] <= 19'd0;
		WeightsStore3[665] <= 19'd0;
		WeightsStore3[666] <= 19'd0;
		WeightsStore3[667] <= 19'd0;
		WeightsStore3[668] <= 19'd0;
		WeightsStore3[669] <= 19'd0;
		WeightsStore3[670] <= 19'd0;
		WeightsStore3[671] <= 19'd0;
		WeightsStore3[672] <= 19'd0;
		WeightsStore3[673] <= 19'd0;
		WeightsStore3[674] <= 19'd0;
		WeightsStore3[675] <= 19'd0;
		WeightsStore3[676] <= 19'd0;
		WeightsStore3[677] <= 19'd0;
		WeightsStore3[678] <= 19'd0;
		WeightsStore3[679] <= 19'd0;
		WeightsStore3[680] <= 19'd0;
		WeightsStore3[681] <= 19'd0;
		WeightsStore3[682] <= 19'd0;
		WeightsStore3[683] <= 19'd0;
		WeightsStore3[684] <= 19'd0;
		WeightsStore3[685] <= 19'd0;
		WeightsStore3[686] <= 19'd0;
		WeightsStore3[687] <= 19'd0;
		WeightsStore3[688] <= 19'd0;
		WeightsStore3[689] <= 19'd0;
		WeightsStore3[690] <= 19'd0;
		WeightsStore3[691] <= 19'd0;
		WeightsStore3[692] <= 19'd0;
		WeightsStore3[693] <= 19'd0;
		WeightsStore3[694] <= 19'd0;
		WeightsStore3[695] <= 19'd0;
		WeightsStore3[696] <= 19'd0;
		WeightsStore3[697] <= 19'd0;
		WeightsStore3[698] <= 19'd0;
		WeightsStore3[699] <= 19'd0;
		WeightsStore3[700] <= 19'd0;
		WeightsStore3[701] <= 19'd0;
		WeightsStore3[702] <= 19'd0;
		WeightsStore3[703] <= 19'd0;
		WeightsStore3[704] <= 19'd0;
		WeightsStore3[705] <= 19'd0;
		WeightsStore3[706] <= 19'd0;
		WeightsStore3[707] <= 19'd0;
		WeightsStore3[708] <= 19'd0;
		WeightsStore3[709] <= 19'd0;
		WeightsStore3[710] <= 19'd0;
		WeightsStore3[711] <= 19'd0;
		WeightsStore3[712] <= 19'd0;
		WeightsStore3[713] <= 19'd0;
		WeightsStore3[714] <= 19'd0;
		WeightsStore3[715] <= 19'd0;
		WeightsStore3[716] <= 19'd0;
		WeightsStore3[717] <= 19'd0;
		WeightsStore3[718] <= 19'd0;
		WeightsStore3[719] <= 19'd0;
		WeightsStore3[720] <= 19'd0;
		WeightsStore3[721] <= 19'd0;
		WeightsStore3[722] <= 19'd0;
		WeightsStore3[723] <= 19'd0;
		WeightsStore3[724] <= 19'd0;
		WeightsStore3[725] <= 19'd0;
		WeightsStore3[726] <= 19'd0;
		WeightsStore3[727] <= 19'd0;
		WeightsStore3[728] <= 19'd0;
		WeightsStore3[729] <= 19'd0;
		WeightsStore3[730] <= 19'd0;
		WeightsStore3[731] <= 19'd0;
		WeightsStore3[732] <= 19'd0;
		WeightsStore3[733] <= 19'd0;
		WeightsStore3[734] <= 19'd0;
		WeightsStore3[735] <= 19'd0;
		WeightsStore3[736] <= 19'd0;
		WeightsStore3[737] <= 19'd0;
		WeightsStore3[738] <= 19'd0;
		WeightsStore3[739] <= 19'd0;
		WeightsStore3[740] <= 19'd0;
		WeightsStore3[741] <= 19'd0;
		WeightsStore3[742] <= 19'd0;
		WeightsStore3[743] <= 19'd0;
		WeightsStore3[744] <= 19'd0;
		WeightsStore3[745] <= 19'd0;
		WeightsStore3[746] <= 19'd0;
		WeightsStore3[747] <= 19'd0;
		WeightsStore3[748] <= 19'd0;
		WeightsStore3[749] <= 19'd0;
		WeightsStore3[750] <= 19'd0;
		WeightsStore3[751] <= 19'd0;
		WeightsStore3[752] <= 19'd0;
		WeightsStore3[753] <= 19'd0;
		WeightsStore3[754] <= 19'd0;
		WeightsStore3[755] <= 19'd0;
		WeightsStore3[756] <= 19'd0;
		WeightsStore3[757] <= 19'd0;
		WeightsStore3[758] <= 19'd0;
		WeightsStore3[759] <= 19'd0;
		WeightsStore3[760] <= 19'd0;
		WeightsStore3[761] <= 19'd0;
		WeightsStore3[762] <= 19'd0;
		WeightsStore3[763] <= 19'd0;
		WeightsStore3[764] <= 19'd0;
		WeightsStore3[765] <= 19'd0;
		WeightsStore3[766] <= 19'd0;
		WeightsStore3[767] <= 19'd0;
		WeightsStore3[768] <= 19'd0;
		WeightsStore3[769] <= 19'd0;
		WeightsStore3[770] <= 19'd0;
		WeightsStore3[771] <= 19'd0;
		WeightsStore3[772] <= 19'd0;
		WeightsStore3[773] <= 19'd0;
		WeightsStore3[774] <= 19'd0;
		WeightsStore3[775] <= 19'd0;
		WeightsStore3[776] <= 19'd0;
		WeightsStore3[777] <= 19'd0;
		WeightsStore3[778] <= 19'd0;
		WeightsStore3[779] <= 19'd0;
		WeightsStore3[780] <= 19'd0;
		WeightsStore3[781] <= 19'd0;
		WeightsStore3[782] <= 19'd0;
		WeightsStore3[783] <= 19'd0;
		WeightsStore3[784] <= 19'd0;
		WeightsStore4[0] <= 19'd0;
		WeightsStore4[1] <= 19'd0;
		WeightsStore4[2] <= 19'd0;
		WeightsStore4[3] <= 19'd0;
		WeightsStore4[4] <= 19'd0;
		WeightsStore4[5] <= 19'd0;
		WeightsStore4[6] <= 19'd0;
		WeightsStore4[7] <= 19'd0;
		WeightsStore4[8] <= 19'd0;
		WeightsStore4[9] <= 19'd0;
		WeightsStore4[10] <= 19'd0;
		WeightsStore4[11] <= 19'd0;
		WeightsStore4[12] <= 19'd0;
		WeightsStore4[13] <= 19'd0;
		WeightsStore4[14] <= 19'd0;
		WeightsStore4[15] <= 19'd0;
		WeightsStore4[16] <= 19'd0;
		WeightsStore4[17] <= 19'd0;
		WeightsStore4[18] <= 19'd0;
		WeightsStore4[19] <= 19'd0;
		WeightsStore4[20] <= 19'd0;
		WeightsStore4[21] <= 19'd0;
		WeightsStore4[22] <= 19'd0;
		WeightsStore4[23] <= 19'd0;
		WeightsStore4[24] <= 19'd0;
		WeightsStore4[25] <= 19'd0;
		WeightsStore4[26] <= 19'd0;
		WeightsStore4[27] <= 19'd0;
		WeightsStore4[28] <= 19'd0;
		WeightsStore4[29] <= 19'd0;
		WeightsStore4[30] <= 19'd0;
		WeightsStore4[31] <= 19'd0;
		WeightsStore4[32] <= 19'd0;
		WeightsStore4[33] <= 19'd0;
		WeightsStore4[34] <= 19'd0;
		WeightsStore4[35] <= 19'd0;
		WeightsStore4[36] <= 19'd0;
		WeightsStore4[37] <= 19'd0;
		WeightsStore4[38] <= 19'd0;
		WeightsStore4[39] <= 19'd0;
		WeightsStore4[40] <= 19'd0;
		WeightsStore4[41] <= 19'd0;
		WeightsStore4[42] <= 19'd0;
		WeightsStore4[43] <= 19'd0;
		WeightsStore4[44] <= 19'd0;
		WeightsStore4[45] <= 19'd0;
		WeightsStore4[46] <= 19'd0;
		WeightsStore4[47] <= 19'd0;
		WeightsStore4[48] <= 19'd0;
		WeightsStore4[49] <= 19'd0;
		WeightsStore4[50] <= 19'd0;
		WeightsStore4[51] <= 19'd0;
		WeightsStore4[52] <= 19'd0;
		WeightsStore4[53] <= 19'd0;
		WeightsStore4[54] <= 19'd0;
		WeightsStore4[55] <= 19'd0;
		WeightsStore4[56] <= 19'd0;
		WeightsStore4[57] <= 19'd0;
		WeightsStore4[58] <= 19'd0;
		WeightsStore4[59] <= 19'd0;
		WeightsStore4[60] <= 19'd0;
		WeightsStore4[61] <= 19'd0;
		WeightsStore4[62] <= 19'd0;
		WeightsStore4[63] <= 19'd0;
		WeightsStore4[64] <= 19'd0;
		WeightsStore4[65] <= 19'd0;
		WeightsStore4[66] <= 19'd0;
		WeightsStore4[67] <= 19'd0;
		WeightsStore4[68] <= 19'd0;
		WeightsStore4[69] <= 19'd0;
		WeightsStore4[70] <= 19'd0;
		WeightsStore4[71] <= 19'd0;
		WeightsStore4[72] <= 19'd0;
		WeightsStore4[73] <= 19'd0;
		WeightsStore4[74] <= 19'd0;
		WeightsStore4[75] <= 19'd0;
		WeightsStore4[76] <= 19'd0;
		WeightsStore4[77] <= 19'd0;
		WeightsStore4[78] <= 19'd0;
		WeightsStore4[79] <= 19'd0;
		WeightsStore4[80] <= 19'd0;
		WeightsStore4[81] <= 19'd0;
		WeightsStore4[82] <= 19'd0;
		WeightsStore4[83] <= 19'd0;
		WeightsStore4[84] <= 19'd0;
		WeightsStore4[85] <= 19'd0;
		WeightsStore4[86] <= 19'd0;
		WeightsStore4[87] <= 19'd0;
		WeightsStore4[88] <= 19'd0;
		WeightsStore4[89] <= 19'd0;
		WeightsStore4[90] <= 19'd0;
		WeightsStore4[91] <= 19'd0;
		WeightsStore4[92] <= 19'd0;
		WeightsStore4[93] <= 19'd0;
		WeightsStore4[94] <= 19'd0;
		WeightsStore4[95] <= 19'd0;
		WeightsStore4[96] <= 19'd0;
		WeightsStore4[97] <= 19'd0;
		WeightsStore4[98] <= 19'd0;
		WeightsStore4[99] <= 19'd0;
		WeightsStore4[100] <= 19'd0;
		WeightsStore4[101] <= 19'd0;
		WeightsStore4[102] <= 19'd0;
		WeightsStore4[103] <= 19'd0;
		WeightsStore4[104] <= 19'd0;
		WeightsStore4[105] <= 19'd0;
		WeightsStore4[106] <= 19'd0;
		WeightsStore4[107] <= 19'd0;
		WeightsStore4[108] <= 19'd0;
		WeightsStore4[109] <= 19'd0;
		WeightsStore4[110] <= 19'd0;
		WeightsStore4[111] <= 19'd0;
		WeightsStore4[112] <= 19'd0;
		WeightsStore4[113] <= 19'd0;
		WeightsStore4[114] <= 19'd0;
		WeightsStore4[115] <= 19'd0;
		WeightsStore4[116] <= 19'd0;
		WeightsStore4[117] <= 19'd0;
		WeightsStore4[118] <= 19'd0;
		WeightsStore4[119] <= 19'd0;
		WeightsStore4[120] <= 19'd0;
		WeightsStore4[121] <= 19'd0;
		WeightsStore4[122] <= 19'd0;
		WeightsStore4[123] <= 19'd0;
		WeightsStore4[124] <= 19'd0;
		WeightsStore4[125] <= 19'd0;
		WeightsStore4[126] <= 19'd0;
		WeightsStore4[127] <= 19'd0;
		WeightsStore4[128] <= 19'd0;
		WeightsStore4[129] <= 19'd0;
		WeightsStore4[130] <= 19'd0;
		WeightsStore4[131] <= 19'd0;
		WeightsStore4[132] <= 19'd0;
		WeightsStore4[133] <= 19'd0;
		WeightsStore4[134] <= 19'd0;
		WeightsStore4[135] <= 19'd0;
		WeightsStore4[136] <= 19'd0;
		WeightsStore4[137] <= 19'd0;
		WeightsStore4[138] <= 19'd0;
		WeightsStore4[139] <= 19'd0;
		WeightsStore4[140] <= 19'd0;
		WeightsStore4[141] <= 19'd0;
		WeightsStore4[142] <= 19'd0;
		WeightsStore4[143] <= 19'd0;
		WeightsStore4[144] <= 19'd0;
		WeightsStore4[145] <= 19'd0;
		WeightsStore4[146] <= 19'd0;
		WeightsStore4[147] <= 19'd0;
		WeightsStore4[148] <= 19'd0;
		WeightsStore4[149] <= 19'd0;
		WeightsStore4[150] <= 19'd0;
		WeightsStore4[151] <= 19'd0;
		WeightsStore4[152] <= 19'd0;
		WeightsStore4[153] <= 19'd0;
		WeightsStore4[154] <= 19'd0;
		WeightsStore4[155] <= 19'd0;
		WeightsStore4[156] <= 19'd0;
		WeightsStore4[157] <= 19'd0;
		WeightsStore4[158] <= 19'd0;
		WeightsStore4[159] <= 19'd0;
		WeightsStore4[160] <= 19'd0;
		WeightsStore4[161] <= 19'd0;
		WeightsStore4[162] <= 19'd0;
		WeightsStore4[163] <= 19'd0;
		WeightsStore4[164] <= 19'd0;
		WeightsStore4[165] <= 19'd0;
		WeightsStore4[166] <= 19'd0;
		WeightsStore4[167] <= 19'd0;
		WeightsStore4[168] <= 19'd0;
		WeightsStore4[169] <= 19'd0;
		WeightsStore4[170] <= 19'd0;
		WeightsStore4[171] <= 19'd0;
		WeightsStore4[172] <= 19'd0;
		WeightsStore4[173] <= 19'd0;
		WeightsStore4[174] <= 19'd0;
		WeightsStore4[175] <= 19'd0;
		WeightsStore4[176] <= 19'd0;
		WeightsStore4[177] <= 19'd0;
		WeightsStore4[178] <= 19'd0;
		WeightsStore4[179] <= 19'd0;
		WeightsStore4[180] <= 19'd0;
		WeightsStore4[181] <= 19'd0;
		WeightsStore4[182] <= 19'd0;
		WeightsStore4[183] <= 19'd0;
		WeightsStore4[184] <= 19'd0;
		WeightsStore4[185] <= 19'd0;
		WeightsStore4[186] <= 19'd0;
		WeightsStore4[187] <= 19'd0;
		WeightsStore4[188] <= 19'd0;
		WeightsStore4[189] <= 19'd0;
		WeightsStore4[190] <= 19'd0;
		WeightsStore4[191] <= 19'd0;
		WeightsStore4[192] <= 19'd0;
		WeightsStore4[193] <= 19'd0;
		WeightsStore4[194] <= 19'd0;
		WeightsStore4[195] <= 19'd0;
		WeightsStore4[196] <= 19'd0;
		WeightsStore4[197] <= 19'd0;
		WeightsStore4[198] <= 19'd0;
		WeightsStore4[199] <= 19'd0;
		WeightsStore4[200] <= 19'd0;
		WeightsStore4[201] <= 19'd0;
		WeightsStore4[202] <= 19'd0;
		WeightsStore4[203] <= 19'd0;
		WeightsStore4[204] <= 19'd0;
		WeightsStore4[205] <= 19'd0;
		WeightsStore4[206] <= 19'd0;
		WeightsStore4[207] <= 19'd0;
		WeightsStore4[208] <= 19'd0;
		WeightsStore4[209] <= 19'd0;
		WeightsStore4[210] <= 19'd0;
		WeightsStore4[211] <= 19'd0;
		WeightsStore4[212] <= 19'd0;
		WeightsStore4[213] <= 19'd0;
		WeightsStore4[214] <= 19'd0;
		WeightsStore4[215] <= 19'd0;
		WeightsStore4[216] <= 19'd0;
		WeightsStore4[217] <= 19'd0;
		WeightsStore4[218] <= 19'd0;
		WeightsStore4[219] <= 19'd0;
		WeightsStore4[220] <= 19'd0;
		WeightsStore4[221] <= 19'd0;
		WeightsStore4[222] <= 19'd0;
		WeightsStore4[223] <= 19'd0;
		WeightsStore4[224] <= 19'd0;
		WeightsStore4[225] <= 19'd0;
		WeightsStore4[226] <= 19'd0;
		WeightsStore4[227] <= 19'd0;
		WeightsStore4[228] <= 19'd0;
		WeightsStore4[229] <= 19'd0;
		WeightsStore4[230] <= 19'd0;
		WeightsStore4[231] <= 19'd0;
		WeightsStore4[232] <= 19'd0;
		WeightsStore4[233] <= 19'd0;
		WeightsStore4[234] <= 19'd0;
		WeightsStore4[235] <= 19'd0;
		WeightsStore4[236] <= 19'd0;
		WeightsStore4[237] <= 19'd0;
		WeightsStore4[238] <= 19'd0;
		WeightsStore4[239] <= 19'd0;
		WeightsStore4[240] <= 19'd0;
		WeightsStore4[241] <= 19'd0;
		WeightsStore4[242] <= 19'd0;
		WeightsStore4[243] <= 19'd0;
		WeightsStore4[244] <= 19'd0;
		WeightsStore4[245] <= 19'd0;
		WeightsStore4[246] <= 19'd0;
		WeightsStore4[247] <= 19'd0;
		WeightsStore4[248] <= 19'd0;
		WeightsStore4[249] <= 19'd0;
		WeightsStore4[250] <= 19'd0;
		WeightsStore4[251] <= 19'd0;
		WeightsStore4[252] <= 19'd0;
		WeightsStore4[253] <= 19'd0;
		WeightsStore4[254] <= 19'd0;
		WeightsStore4[255] <= 19'd0;
		WeightsStore4[256] <= 19'd0;
		WeightsStore4[257] <= 19'd0;
		WeightsStore4[258] <= 19'd0;
		WeightsStore4[259] <= 19'd0;
		WeightsStore4[260] <= 19'd0;
		WeightsStore4[261] <= 19'd0;
		WeightsStore4[262] <= 19'd0;
		WeightsStore4[263] <= 19'd0;
		WeightsStore4[264] <= 19'd0;
		WeightsStore4[265] <= 19'd0;
		WeightsStore4[266] <= 19'd0;
		WeightsStore4[267] <= 19'd0;
		WeightsStore4[268] <= 19'd0;
		WeightsStore4[269] <= 19'd0;
		WeightsStore4[270] <= 19'd0;
		WeightsStore4[271] <= 19'd0;
		WeightsStore4[272] <= 19'd0;
		WeightsStore4[273] <= 19'd0;
		WeightsStore4[274] <= 19'd0;
		WeightsStore4[275] <= 19'd0;
		WeightsStore4[276] <= 19'd0;
		WeightsStore4[277] <= 19'd0;
		WeightsStore4[278] <= 19'd0;
		WeightsStore4[279] <= 19'd0;
		WeightsStore4[280] <= 19'd0;
		WeightsStore4[281] <= 19'd0;
		WeightsStore4[282] <= 19'd0;
		WeightsStore4[283] <= 19'd0;
		WeightsStore4[284] <= 19'd0;
		WeightsStore4[285] <= 19'd0;
		WeightsStore4[286] <= 19'd0;
		WeightsStore4[287] <= 19'd0;
		WeightsStore4[288] <= 19'd0;
		WeightsStore4[289] <= 19'd0;
		WeightsStore4[290] <= 19'd0;
		WeightsStore4[291] <= 19'd0;
		WeightsStore4[292] <= 19'd0;
		WeightsStore4[293] <= 19'd0;
		WeightsStore4[294] <= 19'd0;
		WeightsStore4[295] <= 19'd0;
		WeightsStore4[296] <= 19'd0;
		WeightsStore4[297] <= 19'd0;
		WeightsStore4[298] <= 19'd0;
		WeightsStore4[299] <= 19'd0;
		WeightsStore4[300] <= 19'd0;
		WeightsStore4[301] <= 19'd0;
		WeightsStore4[302] <= 19'd0;
		WeightsStore4[303] <= 19'd0;
		WeightsStore4[304] <= 19'd0;
		WeightsStore4[305] <= 19'd0;
		WeightsStore4[306] <= 19'd0;
		WeightsStore4[307] <= 19'd0;
		WeightsStore4[308] <= 19'd0;
		WeightsStore4[309] <= 19'd0;
		WeightsStore4[310] <= 19'd0;
		WeightsStore4[311] <= 19'd0;
		WeightsStore4[312] <= 19'd0;
		WeightsStore4[313] <= 19'd0;
		WeightsStore4[314] <= 19'd0;
		WeightsStore4[315] <= 19'd0;
		WeightsStore4[316] <= 19'd0;
		WeightsStore4[317] <= 19'd0;
		WeightsStore4[318] <= 19'd0;
		WeightsStore4[319] <= 19'd0;
		WeightsStore4[320] <= 19'd0;
		WeightsStore4[321] <= 19'd0;
		WeightsStore4[322] <= 19'd0;
		WeightsStore4[323] <= 19'd0;
		WeightsStore4[324] <= 19'd0;
		WeightsStore4[325] <= 19'd0;
		WeightsStore4[326] <= 19'd0;
		WeightsStore4[327] <= 19'd0;
		WeightsStore4[328] <= 19'd0;
		WeightsStore4[329] <= 19'd0;
		WeightsStore4[330] <= 19'd0;
		WeightsStore4[331] <= 19'd0;
		WeightsStore4[332] <= 19'd0;
		WeightsStore4[333] <= 19'd0;
		WeightsStore4[334] <= 19'd0;
		WeightsStore4[335] <= 19'd0;
		WeightsStore4[336] <= 19'd0;
		WeightsStore4[337] <= 19'd0;
		WeightsStore4[338] <= 19'd0;
		WeightsStore4[339] <= 19'd0;
		WeightsStore4[340] <= 19'd0;
		WeightsStore4[341] <= 19'd0;
		WeightsStore4[342] <= 19'd0;
		WeightsStore4[343] <= 19'd0;
		WeightsStore4[344] <= 19'd0;
		WeightsStore4[345] <= 19'd0;
		WeightsStore4[346] <= 19'd0;
		WeightsStore4[347] <= 19'd0;
		WeightsStore4[348] <= 19'd0;
		WeightsStore4[349] <= 19'd0;
		WeightsStore4[350] <= 19'd0;
		WeightsStore4[351] <= 19'd0;
		WeightsStore4[352] <= 19'd0;
		WeightsStore4[353] <= 19'd0;
		WeightsStore4[354] <= 19'd0;
		WeightsStore4[355] <= 19'd0;
		WeightsStore4[356] <= 19'd0;
		WeightsStore4[357] <= 19'd0;
		WeightsStore4[358] <= 19'd0;
		WeightsStore4[359] <= 19'd0;
		WeightsStore4[360] <= 19'd0;
		WeightsStore4[361] <= 19'd0;
		WeightsStore4[362] <= 19'd0;
		WeightsStore4[363] <= 19'd0;
		WeightsStore4[364] <= 19'd0;
		WeightsStore4[365] <= 19'd0;
		WeightsStore4[366] <= 19'd0;
		WeightsStore4[367] <= 19'd0;
		WeightsStore4[368] <= 19'd0;
		WeightsStore4[369] <= 19'd0;
		WeightsStore4[370] <= 19'd0;
		WeightsStore4[371] <= 19'd0;
		WeightsStore4[372] <= 19'd0;
		WeightsStore4[373] <= 19'd0;
		WeightsStore4[374] <= 19'd0;
		WeightsStore4[375] <= 19'd0;
		WeightsStore4[376] <= 19'd0;
		WeightsStore4[377] <= 19'd0;
		WeightsStore4[378] <= 19'd0;
		WeightsStore4[379] <= 19'd0;
		WeightsStore4[380] <= 19'd0;
		WeightsStore4[381] <= 19'd0;
		WeightsStore4[382] <= 19'd0;
		WeightsStore4[383] <= 19'd0;
		WeightsStore4[384] <= 19'd0;
		WeightsStore4[385] <= 19'd0;
		WeightsStore4[386] <= 19'd0;
		WeightsStore4[387] <= 19'd0;
		WeightsStore4[388] <= 19'd0;
		WeightsStore4[389] <= 19'd0;
		WeightsStore4[390] <= 19'd0;
		WeightsStore4[391] <= 19'd0;
		WeightsStore4[392] <= 19'd0;
		WeightsStore4[393] <= 19'd0;
		WeightsStore4[394] <= 19'd0;
		WeightsStore4[395] <= 19'd0;
		WeightsStore4[396] <= 19'd0;
		WeightsStore4[397] <= 19'd0;
		WeightsStore4[398] <= 19'd0;
		WeightsStore4[399] <= 19'd0;
		WeightsStore4[400] <= 19'd0;
		WeightsStore4[401] <= 19'd0;
		WeightsStore4[402] <= 19'd0;
		WeightsStore4[403] <= 19'd0;
		WeightsStore4[404] <= 19'd0;
		WeightsStore4[405] <= 19'd0;
		WeightsStore4[406] <= 19'd0;
		WeightsStore4[407] <= 19'd0;
		WeightsStore4[408] <= 19'd0;
		WeightsStore4[409] <= 19'd0;
		WeightsStore4[410] <= 19'd0;
		WeightsStore4[411] <= 19'd0;
		WeightsStore4[412] <= 19'd0;
		WeightsStore4[413] <= 19'd0;
		WeightsStore4[414] <= 19'd0;
		WeightsStore4[415] <= 19'd0;
		WeightsStore4[416] <= 19'd0;
		WeightsStore4[417] <= 19'd0;
		WeightsStore4[418] <= 19'd0;
		WeightsStore4[419] <= 19'd0;
		WeightsStore4[420] <= 19'd0;
		WeightsStore4[421] <= 19'd0;
		WeightsStore4[422] <= 19'd0;
		WeightsStore4[423] <= 19'd0;
		WeightsStore4[424] <= 19'd0;
		WeightsStore4[425] <= 19'd0;
		WeightsStore4[426] <= 19'd0;
		WeightsStore4[427] <= 19'd0;
		WeightsStore4[428] <= 19'd0;
		WeightsStore4[429] <= 19'd0;
		WeightsStore4[430] <= 19'd0;
		WeightsStore4[431] <= 19'd0;
		WeightsStore4[432] <= 19'd0;
		WeightsStore4[433] <= 19'd0;
		WeightsStore4[434] <= 19'd0;
		WeightsStore4[435] <= 19'd0;
		WeightsStore4[436] <= 19'd0;
		WeightsStore4[437] <= 19'd0;
		WeightsStore4[438] <= 19'd0;
		WeightsStore4[439] <= 19'd0;
		WeightsStore4[440] <= 19'd0;
		WeightsStore4[441] <= 19'd0;
		WeightsStore4[442] <= 19'd0;
		WeightsStore4[443] <= 19'd0;
		WeightsStore4[444] <= 19'd0;
		WeightsStore4[445] <= 19'd0;
		WeightsStore4[446] <= 19'd0;
		WeightsStore4[447] <= 19'd0;
		WeightsStore4[448] <= 19'd0;
		WeightsStore4[449] <= 19'd0;
		WeightsStore4[450] <= 19'd0;
		WeightsStore4[451] <= 19'd0;
		WeightsStore4[452] <= 19'd0;
		WeightsStore4[453] <= 19'd0;
		WeightsStore4[454] <= 19'd0;
		WeightsStore4[455] <= 19'd0;
		WeightsStore4[456] <= 19'd0;
		WeightsStore4[457] <= 19'd0;
		WeightsStore4[458] <= 19'd0;
		WeightsStore4[459] <= 19'd0;
		WeightsStore4[460] <= 19'd0;
		WeightsStore4[461] <= 19'd0;
		WeightsStore4[462] <= 19'd0;
		WeightsStore4[463] <= 19'd0;
		WeightsStore4[464] <= 19'd0;
		WeightsStore4[465] <= 19'd0;
		WeightsStore4[466] <= 19'd0;
		WeightsStore4[467] <= 19'd0;
		WeightsStore4[468] <= 19'd0;
		WeightsStore4[469] <= 19'd0;
		WeightsStore4[470] <= 19'd0;
		WeightsStore4[471] <= 19'd0;
		WeightsStore4[472] <= 19'd0;
		WeightsStore4[473] <= 19'd0;
		WeightsStore4[474] <= 19'd0;
		WeightsStore4[475] <= 19'd0;
		WeightsStore4[476] <= 19'd0;
		WeightsStore4[477] <= 19'd0;
		WeightsStore4[478] <= 19'd0;
		WeightsStore4[479] <= 19'd0;
		WeightsStore4[480] <= 19'd0;
		WeightsStore4[481] <= 19'd0;
		WeightsStore4[482] <= 19'd0;
		WeightsStore4[483] <= 19'd0;
		WeightsStore4[484] <= 19'd0;
		WeightsStore4[485] <= 19'd0;
		WeightsStore4[486] <= 19'd0;
		WeightsStore4[487] <= 19'd0;
		WeightsStore4[488] <= 19'd0;
		WeightsStore4[489] <= 19'd0;
		WeightsStore4[490] <= 19'd0;
		WeightsStore4[491] <= 19'd0;
		WeightsStore4[492] <= 19'd0;
		WeightsStore4[493] <= 19'd0;
		WeightsStore4[494] <= 19'd0;
		WeightsStore4[495] <= 19'd0;
		WeightsStore4[496] <= 19'd0;
		WeightsStore4[497] <= 19'd0;
		WeightsStore4[498] <= 19'd0;
		WeightsStore4[499] <= 19'd0;
		WeightsStore4[500] <= 19'd0;
		WeightsStore4[501] <= 19'd0;
		WeightsStore4[502] <= 19'd0;
		WeightsStore4[503] <= 19'd0;
		WeightsStore4[504] <= 19'd0;
		WeightsStore4[505] <= 19'd0;
		WeightsStore4[506] <= 19'd0;
		WeightsStore4[507] <= 19'd0;
		WeightsStore4[508] <= 19'd0;
		WeightsStore4[509] <= 19'd0;
		WeightsStore4[510] <= 19'd0;
		WeightsStore4[511] <= 19'd0;
		WeightsStore4[512] <= 19'd0;
		WeightsStore4[513] <= 19'd0;
		WeightsStore4[514] <= 19'd0;
		WeightsStore4[515] <= 19'd0;
		WeightsStore4[516] <= 19'd0;
		WeightsStore4[517] <= 19'd0;
		WeightsStore4[518] <= 19'd0;
		WeightsStore4[519] <= 19'd0;
		WeightsStore4[520] <= 19'd0;
		WeightsStore4[521] <= 19'd0;
		WeightsStore4[522] <= 19'd0;
		WeightsStore4[523] <= 19'd0;
		WeightsStore4[524] <= 19'd0;
		WeightsStore4[525] <= 19'd0;
		WeightsStore4[526] <= 19'd0;
		WeightsStore4[527] <= 19'd0;
		WeightsStore4[528] <= 19'd0;
		WeightsStore4[529] <= 19'd0;
		WeightsStore4[530] <= 19'd0;
		WeightsStore4[531] <= 19'd0;
		WeightsStore4[532] <= 19'd0;
		WeightsStore4[533] <= 19'd0;
		WeightsStore4[534] <= 19'd0;
		WeightsStore4[535] <= 19'd0;
		WeightsStore4[536] <= 19'd0;
		WeightsStore4[537] <= 19'd0;
		WeightsStore4[538] <= 19'd0;
		WeightsStore4[539] <= 19'd0;
		WeightsStore4[540] <= 19'd0;
		WeightsStore4[541] <= 19'd0;
		WeightsStore4[542] <= 19'd0;
		WeightsStore4[543] <= 19'd0;
		WeightsStore4[544] <= 19'd0;
		WeightsStore4[545] <= 19'd0;
		WeightsStore4[546] <= 19'd0;
		WeightsStore4[547] <= 19'd0;
		WeightsStore4[548] <= 19'd0;
		WeightsStore4[549] <= 19'd0;
		WeightsStore4[550] <= 19'd0;
		WeightsStore4[551] <= 19'd0;
		WeightsStore4[552] <= 19'd0;
		WeightsStore4[553] <= 19'd0;
		WeightsStore4[554] <= 19'd0;
		WeightsStore4[555] <= 19'd0;
		WeightsStore4[556] <= 19'd0;
		WeightsStore4[557] <= 19'd0;
		WeightsStore4[558] <= 19'd0;
		WeightsStore4[559] <= 19'd0;
		WeightsStore4[560] <= 19'd0;
		WeightsStore4[561] <= 19'd0;
		WeightsStore4[562] <= 19'd0;
		WeightsStore4[563] <= 19'd0;
		WeightsStore4[564] <= 19'd0;
		WeightsStore4[565] <= 19'd0;
		WeightsStore4[566] <= 19'd0;
		WeightsStore4[567] <= 19'd0;
		WeightsStore4[568] <= 19'd0;
		WeightsStore4[569] <= 19'd0;
		WeightsStore4[570] <= 19'd0;
		WeightsStore4[571] <= 19'd0;
		WeightsStore4[572] <= 19'd0;
		WeightsStore4[573] <= 19'd0;
		WeightsStore4[574] <= 19'd0;
		WeightsStore4[575] <= 19'd0;
		WeightsStore4[576] <= 19'd0;
		WeightsStore4[577] <= 19'd0;
		WeightsStore4[578] <= 19'd0;
		WeightsStore4[579] <= 19'd0;
		WeightsStore4[580] <= 19'd0;
		WeightsStore4[581] <= 19'd0;
		WeightsStore4[582] <= 19'd0;
		WeightsStore4[583] <= 19'd0;
		WeightsStore4[584] <= 19'd0;
		WeightsStore4[585] <= 19'd0;
		WeightsStore4[586] <= 19'd0;
		WeightsStore4[587] <= 19'd0;
		WeightsStore4[588] <= 19'd0;
		WeightsStore4[589] <= 19'd0;
		WeightsStore4[590] <= 19'd0;
		WeightsStore4[591] <= 19'd0;
		WeightsStore4[592] <= 19'd0;
		WeightsStore4[593] <= 19'd0;
		WeightsStore4[594] <= 19'd0;
		WeightsStore4[595] <= 19'd0;
		WeightsStore4[596] <= 19'd0;
		WeightsStore4[597] <= 19'd0;
		WeightsStore4[598] <= 19'd0;
		WeightsStore4[599] <= 19'd0;
		WeightsStore4[600] <= 19'd0;
		WeightsStore4[601] <= 19'd0;
		WeightsStore4[602] <= 19'd0;
		WeightsStore4[603] <= 19'd0;
		WeightsStore4[604] <= 19'd0;
		WeightsStore4[605] <= 19'd0;
		WeightsStore4[606] <= 19'd0;
		WeightsStore4[607] <= 19'd0;
		WeightsStore4[608] <= 19'd0;
		WeightsStore4[609] <= 19'd0;
		WeightsStore4[610] <= 19'd0;
		WeightsStore4[611] <= 19'd0;
		WeightsStore4[612] <= 19'd0;
		WeightsStore4[613] <= 19'd0;
		WeightsStore4[614] <= 19'd0;
		WeightsStore4[615] <= 19'd0;
		WeightsStore4[616] <= 19'd0;
		WeightsStore4[617] <= 19'd0;
		WeightsStore4[618] <= 19'd0;
		WeightsStore4[619] <= 19'd0;
		WeightsStore4[620] <= 19'd0;
		WeightsStore4[621] <= 19'd0;
		WeightsStore4[622] <= 19'd0;
		WeightsStore4[623] <= 19'd0;
		WeightsStore4[624] <= 19'd0;
		WeightsStore4[625] <= 19'd0;
		WeightsStore4[626] <= 19'd0;
		WeightsStore4[627] <= 19'd0;
		WeightsStore4[628] <= 19'd0;
		WeightsStore4[629] <= 19'd0;
		WeightsStore4[630] <= 19'd0;
		WeightsStore4[631] <= 19'd0;
		WeightsStore4[632] <= 19'd0;
		WeightsStore4[633] <= 19'd0;
		WeightsStore4[634] <= 19'd0;
		WeightsStore4[635] <= 19'd0;
		WeightsStore4[636] <= 19'd0;
		WeightsStore4[637] <= 19'd0;
		WeightsStore4[638] <= 19'd0;
		WeightsStore4[639] <= 19'd0;
		WeightsStore4[640] <= 19'd0;
		WeightsStore4[641] <= 19'd0;
		WeightsStore4[642] <= 19'd0;
		WeightsStore4[643] <= 19'd0;
		WeightsStore4[644] <= 19'd0;
		WeightsStore4[645] <= 19'd0;
		WeightsStore4[646] <= 19'd0;
		WeightsStore4[647] <= 19'd0;
		WeightsStore4[648] <= 19'd0;
		WeightsStore4[649] <= 19'd0;
		WeightsStore4[650] <= 19'd0;
		WeightsStore4[651] <= 19'd0;
		WeightsStore4[652] <= 19'd0;
		WeightsStore4[653] <= 19'd0;
		WeightsStore4[654] <= 19'd0;
		WeightsStore4[655] <= 19'd0;
		WeightsStore4[656] <= 19'd0;
		WeightsStore4[657] <= 19'd0;
		WeightsStore4[658] <= 19'd0;
		WeightsStore4[659] <= 19'd0;
		WeightsStore4[660] <= 19'd0;
		WeightsStore4[661] <= 19'd0;
		WeightsStore4[662] <= 19'd0;
		WeightsStore4[663] <= 19'd0;
		WeightsStore4[664] <= 19'd0;
		WeightsStore4[665] <= 19'd0;
		WeightsStore4[666] <= 19'd0;
		WeightsStore4[667] <= 19'd0;
		WeightsStore4[668] <= 19'd0;
		WeightsStore4[669] <= 19'd0;
		WeightsStore4[670] <= 19'd0;
		WeightsStore4[671] <= 19'd0;
		WeightsStore4[672] <= 19'd0;
		WeightsStore4[673] <= 19'd0;
		WeightsStore4[674] <= 19'd0;
		WeightsStore4[675] <= 19'd0;
		WeightsStore4[676] <= 19'd0;
		WeightsStore4[677] <= 19'd0;
		WeightsStore4[678] <= 19'd0;
		WeightsStore4[679] <= 19'd0;
		WeightsStore4[680] <= 19'd0;
		WeightsStore4[681] <= 19'd0;
		WeightsStore4[682] <= 19'd0;
		WeightsStore4[683] <= 19'd0;
		WeightsStore4[684] <= 19'd0;
		WeightsStore4[685] <= 19'd0;
		WeightsStore4[686] <= 19'd0;
		WeightsStore4[687] <= 19'd0;
		WeightsStore4[688] <= 19'd0;
		WeightsStore4[689] <= 19'd0;
		WeightsStore4[690] <= 19'd0;
		WeightsStore4[691] <= 19'd0;
		WeightsStore4[692] <= 19'd0;
		WeightsStore4[693] <= 19'd0;
		WeightsStore4[694] <= 19'd0;
		WeightsStore4[695] <= 19'd0;
		WeightsStore4[696] <= 19'd0;
		WeightsStore4[697] <= 19'd0;
		WeightsStore4[698] <= 19'd0;
		WeightsStore4[699] <= 19'd0;
		WeightsStore4[700] <= 19'd0;
		WeightsStore4[701] <= 19'd0;
		WeightsStore4[702] <= 19'd0;
		WeightsStore4[703] <= 19'd0;
		WeightsStore4[704] <= 19'd0;
		WeightsStore4[705] <= 19'd0;
		WeightsStore4[706] <= 19'd0;
		WeightsStore4[707] <= 19'd0;
		WeightsStore4[708] <= 19'd0;
		WeightsStore4[709] <= 19'd0;
		WeightsStore4[710] <= 19'd0;
		WeightsStore4[711] <= 19'd0;
		WeightsStore4[712] <= 19'd0;
		WeightsStore4[713] <= 19'd0;
		WeightsStore4[714] <= 19'd0;
		WeightsStore4[715] <= 19'd0;
		WeightsStore4[716] <= 19'd0;
		WeightsStore4[717] <= 19'd0;
		WeightsStore4[718] <= 19'd0;
		WeightsStore4[719] <= 19'd0;
		WeightsStore4[720] <= 19'd0;
		WeightsStore4[721] <= 19'd0;
		WeightsStore4[722] <= 19'd0;
		WeightsStore4[723] <= 19'd0;
		WeightsStore4[724] <= 19'd0;
		WeightsStore4[725] <= 19'd0;
		WeightsStore4[726] <= 19'd0;
		WeightsStore4[727] <= 19'd0;
		WeightsStore4[728] <= 19'd0;
		WeightsStore4[729] <= 19'd0;
		WeightsStore4[730] <= 19'd0;
		WeightsStore4[731] <= 19'd0;
		WeightsStore4[732] <= 19'd0;
		WeightsStore4[733] <= 19'd0;
		WeightsStore4[734] <= 19'd0;
		WeightsStore4[735] <= 19'd0;
		WeightsStore4[736] <= 19'd0;
		WeightsStore4[737] <= 19'd0;
		WeightsStore4[738] <= 19'd0;
		WeightsStore4[739] <= 19'd0;
		WeightsStore4[740] <= 19'd0;
		WeightsStore4[741] <= 19'd0;
		WeightsStore4[742] <= 19'd0;
		WeightsStore4[743] <= 19'd0;
		WeightsStore4[744] <= 19'd0;
		WeightsStore4[745] <= 19'd0;
		WeightsStore4[746] <= 19'd0;
		WeightsStore4[747] <= 19'd0;
		WeightsStore4[748] <= 19'd0;
		WeightsStore4[749] <= 19'd0;
		WeightsStore4[750] <= 19'd0;
		WeightsStore4[751] <= 19'd0;
		WeightsStore4[752] <= 19'd0;
		WeightsStore4[753] <= 19'd0;
		WeightsStore4[754] <= 19'd0;
		WeightsStore4[755] <= 19'd0;
		WeightsStore4[756] <= 19'd0;
		WeightsStore4[757] <= 19'd0;
		WeightsStore4[758] <= 19'd0;
		WeightsStore4[759] <= 19'd0;
		WeightsStore4[760] <= 19'd0;
		WeightsStore4[761] <= 19'd0;
		WeightsStore4[762] <= 19'd0;
		WeightsStore4[763] <= 19'd0;
		WeightsStore4[764] <= 19'd0;
		WeightsStore4[765] <= 19'd0;
		WeightsStore4[766] <= 19'd0;
		WeightsStore4[767] <= 19'd0;
		WeightsStore4[768] <= 19'd0;
		WeightsStore4[769] <= 19'd0;
		WeightsStore4[770] <= 19'd0;
		WeightsStore4[771] <= 19'd0;
		WeightsStore4[772] <= 19'd0;
		WeightsStore4[773] <= 19'd0;
		WeightsStore4[774] <= 19'd0;
		WeightsStore4[775] <= 19'd0;
		WeightsStore4[776] <= 19'd0;
		WeightsStore4[777] <= 19'd0;
		WeightsStore4[778] <= 19'd0;
		WeightsStore4[779] <= 19'd0;
		WeightsStore4[780] <= 19'd0;
		WeightsStore4[781] <= 19'd0;
		WeightsStore4[782] <= 19'd0;
		WeightsStore4[783] <= 19'd0;
		WeightsStore4[784] <= 19'd0;
		WeightsStore5[0] <= 19'd0;
		WeightsStore5[1] <= 19'd0;
		WeightsStore5[2] <= 19'd0;
		WeightsStore5[3] <= 19'd0;
		WeightsStore5[4] <= 19'd0;
		WeightsStore5[5] <= 19'd0;
		WeightsStore5[6] <= 19'd0;
		WeightsStore5[7] <= 19'd0;
		WeightsStore5[8] <= 19'd0;
		WeightsStore5[9] <= 19'd0;
		WeightsStore5[10] <= 19'd0;
		WeightsStore5[11] <= 19'd0;
		WeightsStore5[12] <= 19'd0;
		WeightsStore5[13] <= 19'd0;
		WeightsStore5[14] <= 19'd0;
		WeightsStore5[15] <= 19'd0;
		WeightsStore5[16] <= 19'd0;
		WeightsStore5[17] <= 19'd0;
		WeightsStore5[18] <= 19'd0;
		WeightsStore5[19] <= 19'd0;
		WeightsStore5[20] <= 19'd0;
		WeightsStore5[21] <= 19'd0;
		WeightsStore5[22] <= 19'd0;
		WeightsStore5[23] <= 19'd0;
		WeightsStore5[24] <= 19'd0;
		WeightsStore5[25] <= 19'd0;
		WeightsStore5[26] <= 19'd0;
		WeightsStore5[27] <= 19'd0;
		WeightsStore5[28] <= 19'd0;
		WeightsStore5[29] <= 19'd0;
		WeightsStore5[30] <= 19'd0;
		WeightsStore5[31] <= 19'd0;
		WeightsStore5[32] <= 19'd0;
		WeightsStore5[33] <= 19'd0;
		WeightsStore5[34] <= 19'd0;
		WeightsStore5[35] <= 19'd0;
		WeightsStore5[36] <= 19'd0;
		WeightsStore5[37] <= 19'd0;
		WeightsStore5[38] <= 19'd0;
		WeightsStore5[39] <= 19'd0;
		WeightsStore5[40] <= 19'd0;
		WeightsStore5[41] <= 19'd0;
		WeightsStore5[42] <= 19'd0;
		WeightsStore5[43] <= 19'd0;
		WeightsStore5[44] <= 19'd0;
		WeightsStore5[45] <= 19'd0;
		WeightsStore5[46] <= 19'd0;
		WeightsStore5[47] <= 19'd0;
		WeightsStore5[48] <= 19'd0;
		WeightsStore5[49] <= 19'd0;
		WeightsStore5[50] <= 19'd0;
		WeightsStore5[51] <= 19'd0;
		WeightsStore5[52] <= 19'd0;
		WeightsStore5[53] <= 19'd0;
		WeightsStore5[54] <= 19'd0;
		WeightsStore5[55] <= 19'd0;
		WeightsStore5[56] <= 19'd0;
		WeightsStore5[57] <= 19'd0;
		WeightsStore5[58] <= 19'd0;
		WeightsStore5[59] <= 19'd0;
		WeightsStore5[60] <= 19'd0;
		WeightsStore5[61] <= 19'd0;
		WeightsStore5[62] <= 19'd0;
		WeightsStore5[63] <= 19'd0;
		WeightsStore5[64] <= 19'd0;
		WeightsStore5[65] <= 19'd0;
		WeightsStore5[66] <= 19'd0;
		WeightsStore5[67] <= 19'd0;
		WeightsStore5[68] <= 19'd0;
		WeightsStore5[69] <= 19'd0;
		WeightsStore5[70] <= 19'd0;
		WeightsStore5[71] <= 19'd0;
		WeightsStore5[72] <= 19'd0;
		WeightsStore5[73] <= 19'd0;
		WeightsStore5[74] <= 19'd0;
		WeightsStore5[75] <= 19'd0;
		WeightsStore5[76] <= 19'd0;
		WeightsStore5[77] <= 19'd0;
		WeightsStore5[78] <= 19'd0;
		WeightsStore5[79] <= 19'd0;
		WeightsStore5[80] <= 19'd0;
		WeightsStore5[81] <= 19'd0;
		WeightsStore5[82] <= 19'd0;
		WeightsStore5[83] <= 19'd0;
		WeightsStore5[84] <= 19'd0;
		WeightsStore5[85] <= 19'd0;
		WeightsStore5[86] <= 19'd0;
		WeightsStore5[87] <= 19'd0;
		WeightsStore5[88] <= 19'd0;
		WeightsStore5[89] <= 19'd0;
		WeightsStore5[90] <= 19'd0;
		WeightsStore5[91] <= 19'd0;
		WeightsStore5[92] <= 19'd0;
		WeightsStore5[93] <= 19'd0;
		WeightsStore5[94] <= 19'd0;
		WeightsStore5[95] <= 19'd0;
		WeightsStore5[96] <= 19'd0;
		WeightsStore5[97] <= 19'd0;
		WeightsStore5[98] <= 19'd0;
		WeightsStore5[99] <= 19'd0;
		WeightsStore5[100] <= 19'd0;
		WeightsStore5[101] <= 19'd0;
		WeightsStore5[102] <= 19'd0;
		WeightsStore5[103] <= 19'd0;
		WeightsStore5[104] <= 19'd0;
		WeightsStore5[105] <= 19'd0;
		WeightsStore5[106] <= 19'd0;
		WeightsStore5[107] <= 19'd0;
		WeightsStore5[108] <= 19'd0;
		WeightsStore5[109] <= 19'd0;
		WeightsStore5[110] <= 19'd0;
		WeightsStore5[111] <= 19'd0;
		WeightsStore5[112] <= 19'd0;
		WeightsStore5[113] <= 19'd0;
		WeightsStore5[114] <= 19'd0;
		WeightsStore5[115] <= 19'd0;
		WeightsStore5[116] <= 19'd0;
		WeightsStore5[117] <= 19'd0;
		WeightsStore5[118] <= 19'd0;
		WeightsStore5[119] <= 19'd0;
		WeightsStore5[120] <= 19'd0;
		WeightsStore5[121] <= 19'd0;
		WeightsStore5[122] <= 19'd0;
		WeightsStore5[123] <= 19'd0;
		WeightsStore5[124] <= 19'd0;
		WeightsStore5[125] <= 19'd0;
		WeightsStore5[126] <= 19'd0;
		WeightsStore5[127] <= 19'd0;
		WeightsStore5[128] <= 19'd0;
		WeightsStore5[129] <= 19'd0;
		WeightsStore5[130] <= 19'd0;
		WeightsStore5[131] <= 19'd0;
		WeightsStore5[132] <= 19'd0;
		WeightsStore5[133] <= 19'd0;
		WeightsStore5[134] <= 19'd0;
		WeightsStore5[135] <= 19'd0;
		WeightsStore5[136] <= 19'd0;
		WeightsStore5[137] <= 19'd0;
		WeightsStore5[138] <= 19'd0;
		WeightsStore5[139] <= 19'd0;
		WeightsStore5[140] <= 19'd0;
		WeightsStore5[141] <= 19'd0;
		WeightsStore5[142] <= 19'd0;
		WeightsStore5[143] <= 19'd0;
		WeightsStore5[144] <= 19'd0;
		WeightsStore5[145] <= 19'd0;
		WeightsStore5[146] <= 19'd0;
		WeightsStore5[147] <= 19'd0;
		WeightsStore5[148] <= 19'd0;
		WeightsStore5[149] <= 19'd0;
		WeightsStore5[150] <= 19'd0;
		WeightsStore5[151] <= 19'd0;
		WeightsStore5[152] <= 19'd0;
		WeightsStore5[153] <= 19'd0;
		WeightsStore5[154] <= 19'd0;
		WeightsStore5[155] <= 19'd0;
		WeightsStore5[156] <= 19'd0;
		WeightsStore5[157] <= 19'd0;
		WeightsStore5[158] <= 19'd0;
		WeightsStore5[159] <= 19'd0;
		WeightsStore5[160] <= 19'd0;
		WeightsStore5[161] <= 19'd0;
		WeightsStore5[162] <= 19'd0;
		WeightsStore5[163] <= 19'd0;
		WeightsStore5[164] <= 19'd0;
		WeightsStore5[165] <= 19'd0;
		WeightsStore5[166] <= 19'd0;
		WeightsStore5[167] <= 19'd0;
		WeightsStore5[168] <= 19'd0;
		WeightsStore5[169] <= 19'd0;
		WeightsStore5[170] <= 19'd0;
		WeightsStore5[171] <= 19'd0;
		WeightsStore5[172] <= 19'd0;
		WeightsStore5[173] <= 19'd0;
		WeightsStore5[174] <= 19'd0;
		WeightsStore5[175] <= 19'd0;
		WeightsStore5[176] <= 19'd0;
		WeightsStore5[177] <= 19'd0;
		WeightsStore5[178] <= 19'd0;
		WeightsStore5[179] <= 19'd0;
		WeightsStore5[180] <= 19'd0;
		WeightsStore5[181] <= 19'd0;
		WeightsStore5[182] <= 19'd0;
		WeightsStore5[183] <= 19'd0;
		WeightsStore5[184] <= 19'd0;
		WeightsStore5[185] <= 19'd0;
		WeightsStore5[186] <= 19'd0;
		WeightsStore5[187] <= 19'd0;
		WeightsStore5[188] <= 19'd0;
		WeightsStore5[189] <= 19'd0;
		WeightsStore5[190] <= 19'd0;
		WeightsStore5[191] <= 19'd0;
		WeightsStore5[192] <= 19'd0;
		WeightsStore5[193] <= 19'd0;
		WeightsStore5[194] <= 19'd0;
		WeightsStore5[195] <= 19'd0;
		WeightsStore5[196] <= 19'd0;
		WeightsStore5[197] <= 19'd0;
		WeightsStore5[198] <= 19'd0;
		WeightsStore5[199] <= 19'd0;
		WeightsStore5[200] <= 19'd0;
		WeightsStore5[201] <= 19'd0;
		WeightsStore5[202] <= 19'd0;
		WeightsStore5[203] <= 19'd0;
		WeightsStore5[204] <= 19'd0;
		WeightsStore5[205] <= 19'd0;
		WeightsStore5[206] <= 19'd0;
		WeightsStore5[207] <= 19'd0;
		WeightsStore5[208] <= 19'd0;
		WeightsStore5[209] <= 19'd0;
		WeightsStore5[210] <= 19'd0;
		WeightsStore5[211] <= 19'd0;
		WeightsStore5[212] <= 19'd0;
		WeightsStore5[213] <= 19'd0;
		WeightsStore5[214] <= 19'd0;
		WeightsStore5[215] <= 19'd0;
		WeightsStore5[216] <= 19'd0;
		WeightsStore5[217] <= 19'd0;
		WeightsStore5[218] <= 19'd0;
		WeightsStore5[219] <= 19'd0;
		WeightsStore5[220] <= 19'd0;
		WeightsStore5[221] <= 19'd0;
		WeightsStore5[222] <= 19'd0;
		WeightsStore5[223] <= 19'd0;
		WeightsStore5[224] <= 19'd0;
		WeightsStore5[225] <= 19'd0;
		WeightsStore5[226] <= 19'd0;
		WeightsStore5[227] <= 19'd0;
		WeightsStore5[228] <= 19'd0;
		WeightsStore5[229] <= 19'd0;
		WeightsStore5[230] <= 19'd0;
		WeightsStore5[231] <= 19'd0;
		WeightsStore5[232] <= 19'd0;
		WeightsStore5[233] <= 19'd0;
		WeightsStore5[234] <= 19'd0;
		WeightsStore5[235] <= 19'd0;
		WeightsStore5[236] <= 19'd0;
		WeightsStore5[237] <= 19'd0;
		WeightsStore5[238] <= 19'd0;
		WeightsStore5[239] <= 19'd0;
		WeightsStore5[240] <= 19'd0;
		WeightsStore5[241] <= 19'd0;
		WeightsStore5[242] <= 19'd0;
		WeightsStore5[243] <= 19'd0;
		WeightsStore5[244] <= 19'd0;
		WeightsStore5[245] <= 19'd0;
		WeightsStore5[246] <= 19'd0;
		WeightsStore5[247] <= 19'd0;
		WeightsStore5[248] <= 19'd0;
		WeightsStore5[249] <= 19'd0;
		WeightsStore5[250] <= 19'd0;
		WeightsStore5[251] <= 19'd0;
		WeightsStore5[252] <= 19'd0;
		WeightsStore5[253] <= 19'd0;
		WeightsStore5[254] <= 19'd0;
		WeightsStore5[255] <= 19'd0;
		WeightsStore5[256] <= 19'd0;
		WeightsStore5[257] <= 19'd0;
		WeightsStore5[258] <= 19'd0;
		WeightsStore5[259] <= 19'd0;
		WeightsStore5[260] <= 19'd0;
		WeightsStore5[261] <= 19'd0;
		WeightsStore5[262] <= 19'd0;
		WeightsStore5[263] <= 19'd0;
		WeightsStore5[264] <= 19'd0;
		WeightsStore5[265] <= 19'd0;
		WeightsStore5[266] <= 19'd0;
		WeightsStore5[267] <= 19'd0;
		WeightsStore5[268] <= 19'd0;
		WeightsStore5[269] <= 19'd0;
		WeightsStore5[270] <= 19'd0;
		WeightsStore5[271] <= 19'd0;
		WeightsStore5[272] <= 19'd0;
		WeightsStore5[273] <= 19'd0;
		WeightsStore5[274] <= 19'd0;
		WeightsStore5[275] <= 19'd0;
		WeightsStore5[276] <= 19'd0;
		WeightsStore5[277] <= 19'd0;
		WeightsStore5[278] <= 19'd0;
		WeightsStore5[279] <= 19'd0;
		WeightsStore5[280] <= 19'd0;
		WeightsStore5[281] <= 19'd0;
		WeightsStore5[282] <= 19'd0;
		WeightsStore5[283] <= 19'd0;
		WeightsStore5[284] <= 19'd0;
		WeightsStore5[285] <= 19'd0;
		WeightsStore5[286] <= 19'd0;
		WeightsStore5[287] <= 19'd0;
		WeightsStore5[288] <= 19'd0;
		WeightsStore5[289] <= 19'd0;
		WeightsStore5[290] <= 19'd0;
		WeightsStore5[291] <= 19'd0;
		WeightsStore5[292] <= 19'd0;
		WeightsStore5[293] <= 19'd0;
		WeightsStore5[294] <= 19'd0;
		WeightsStore5[295] <= 19'd0;
		WeightsStore5[296] <= 19'd0;
		WeightsStore5[297] <= 19'd0;
		WeightsStore5[298] <= 19'd0;
		WeightsStore5[299] <= 19'd0;
		WeightsStore5[300] <= 19'd0;
		WeightsStore5[301] <= 19'd0;
		WeightsStore5[302] <= 19'd0;
		WeightsStore5[303] <= 19'd0;
		WeightsStore5[304] <= 19'd0;
		WeightsStore5[305] <= 19'd0;
		WeightsStore5[306] <= 19'd0;
		WeightsStore5[307] <= 19'd0;
		WeightsStore5[308] <= 19'd0;
		WeightsStore5[309] <= 19'd0;
		WeightsStore5[310] <= 19'd0;
		WeightsStore5[311] <= 19'd0;
		WeightsStore5[312] <= 19'd0;
		WeightsStore5[313] <= 19'd0;
		WeightsStore5[314] <= 19'd0;
		WeightsStore5[315] <= 19'd0;
		WeightsStore5[316] <= 19'd0;
		WeightsStore5[317] <= 19'd0;
		WeightsStore5[318] <= 19'd0;
		WeightsStore5[319] <= 19'd0;
		WeightsStore5[320] <= 19'd0;
		WeightsStore5[321] <= 19'd0;
		WeightsStore5[322] <= 19'd0;
		WeightsStore5[323] <= 19'd0;
		WeightsStore5[324] <= 19'd0;
		WeightsStore5[325] <= 19'd0;
		WeightsStore5[326] <= 19'd0;
		WeightsStore5[327] <= 19'd0;
		WeightsStore5[328] <= 19'd0;
		WeightsStore5[329] <= 19'd0;
		WeightsStore5[330] <= 19'd0;
		WeightsStore5[331] <= 19'd0;
		WeightsStore5[332] <= 19'd0;
		WeightsStore5[333] <= 19'd0;
		WeightsStore5[334] <= 19'd0;
		WeightsStore5[335] <= 19'd0;
		WeightsStore5[336] <= 19'd0;
		WeightsStore5[337] <= 19'd0;
		WeightsStore5[338] <= 19'd0;
		WeightsStore5[339] <= 19'd0;
		WeightsStore5[340] <= 19'd0;
		WeightsStore5[341] <= 19'd0;
		WeightsStore5[342] <= 19'd0;
		WeightsStore5[343] <= 19'd0;
		WeightsStore5[344] <= 19'd0;
		WeightsStore5[345] <= 19'd0;
		WeightsStore5[346] <= 19'd0;
		WeightsStore5[347] <= 19'd0;
		WeightsStore5[348] <= 19'd0;
		WeightsStore5[349] <= 19'd0;
		WeightsStore5[350] <= 19'd0;
		WeightsStore5[351] <= 19'd0;
		WeightsStore5[352] <= 19'd0;
		WeightsStore5[353] <= 19'd0;
		WeightsStore5[354] <= 19'd0;
		WeightsStore5[355] <= 19'd0;
		WeightsStore5[356] <= 19'd0;
		WeightsStore5[357] <= 19'd0;
		WeightsStore5[358] <= 19'd0;
		WeightsStore5[359] <= 19'd0;
		WeightsStore5[360] <= 19'd0;
		WeightsStore5[361] <= 19'd0;
		WeightsStore5[362] <= 19'd0;
		WeightsStore5[363] <= 19'd0;
		WeightsStore5[364] <= 19'd0;
		WeightsStore5[365] <= 19'd0;
		WeightsStore5[366] <= 19'd0;
		WeightsStore5[367] <= 19'd0;
		WeightsStore5[368] <= 19'd0;
		WeightsStore5[369] <= 19'd0;
		WeightsStore5[370] <= 19'd0;
		WeightsStore5[371] <= 19'd0;
		WeightsStore5[372] <= 19'd0;
		WeightsStore5[373] <= 19'd0;
		WeightsStore5[374] <= 19'd0;
		WeightsStore5[375] <= 19'd0;
		WeightsStore5[376] <= 19'd0;
		WeightsStore5[377] <= 19'd0;
		WeightsStore5[378] <= 19'd0;
		WeightsStore5[379] <= 19'd0;
		WeightsStore5[380] <= 19'd0;
		WeightsStore5[381] <= 19'd0;
		WeightsStore5[382] <= 19'd0;
		WeightsStore5[383] <= 19'd0;
		WeightsStore5[384] <= 19'd0;
		WeightsStore5[385] <= 19'd0;
		WeightsStore5[386] <= 19'd0;
		WeightsStore5[387] <= 19'd0;
		WeightsStore5[388] <= 19'd0;
		WeightsStore5[389] <= 19'd0;
		WeightsStore5[390] <= 19'd0;
		WeightsStore5[391] <= 19'd0;
		WeightsStore5[392] <= 19'd0;
		WeightsStore5[393] <= 19'd0;
		WeightsStore5[394] <= 19'd0;
		WeightsStore5[395] <= 19'd0;
		WeightsStore5[396] <= 19'd0;
		WeightsStore5[397] <= 19'd0;
		WeightsStore5[398] <= 19'd0;
		WeightsStore5[399] <= 19'd0;
		WeightsStore5[400] <= 19'd0;
		WeightsStore5[401] <= 19'd0;
		WeightsStore5[402] <= 19'd0;
		WeightsStore5[403] <= 19'd0;
		WeightsStore5[404] <= 19'd0;
		WeightsStore5[405] <= 19'd0;
		WeightsStore5[406] <= 19'd0;
		WeightsStore5[407] <= 19'd0;
		WeightsStore5[408] <= 19'd0;
		WeightsStore5[409] <= 19'd0;
		WeightsStore5[410] <= 19'd0;
		WeightsStore5[411] <= 19'd0;
		WeightsStore5[412] <= 19'd0;
		WeightsStore5[413] <= 19'd0;
		WeightsStore5[414] <= 19'd0;
		WeightsStore5[415] <= 19'd0;
		WeightsStore5[416] <= 19'd0;
		WeightsStore5[417] <= 19'd0;
		WeightsStore5[418] <= 19'd0;
		WeightsStore5[419] <= 19'd0;
		WeightsStore5[420] <= 19'd0;
		WeightsStore5[421] <= 19'd0;
		WeightsStore5[422] <= 19'd0;
		WeightsStore5[423] <= 19'd0;
		WeightsStore5[424] <= 19'd0;
		WeightsStore5[425] <= 19'd0;
		WeightsStore5[426] <= 19'd0;
		WeightsStore5[427] <= 19'd0;
		WeightsStore5[428] <= 19'd0;
		WeightsStore5[429] <= 19'd0;
		WeightsStore5[430] <= 19'd0;
		WeightsStore5[431] <= 19'd0;
		WeightsStore5[432] <= 19'd0;
		WeightsStore5[433] <= 19'd0;
		WeightsStore5[434] <= 19'd0;
		WeightsStore5[435] <= 19'd0;
		WeightsStore5[436] <= 19'd0;
		WeightsStore5[437] <= 19'd0;
		WeightsStore5[438] <= 19'd0;
		WeightsStore5[439] <= 19'd0;
		WeightsStore5[440] <= 19'd0;
		WeightsStore5[441] <= 19'd0;
		WeightsStore5[442] <= 19'd0;
		WeightsStore5[443] <= 19'd0;
		WeightsStore5[444] <= 19'd0;
		WeightsStore5[445] <= 19'd0;
		WeightsStore5[446] <= 19'd0;
		WeightsStore5[447] <= 19'd0;
		WeightsStore5[448] <= 19'd0;
		WeightsStore5[449] <= 19'd0;
		WeightsStore5[450] <= 19'd0;
		WeightsStore5[451] <= 19'd0;
		WeightsStore5[452] <= 19'd0;
		WeightsStore5[453] <= 19'd0;
		WeightsStore5[454] <= 19'd0;
		WeightsStore5[455] <= 19'd0;
		WeightsStore5[456] <= 19'd0;
		WeightsStore5[457] <= 19'd0;
		WeightsStore5[458] <= 19'd0;
		WeightsStore5[459] <= 19'd0;
		WeightsStore5[460] <= 19'd0;
		WeightsStore5[461] <= 19'd0;
		WeightsStore5[462] <= 19'd0;
		WeightsStore5[463] <= 19'd0;
		WeightsStore5[464] <= 19'd0;
		WeightsStore5[465] <= 19'd0;
		WeightsStore5[466] <= 19'd0;
		WeightsStore5[467] <= 19'd0;
		WeightsStore5[468] <= 19'd0;
		WeightsStore5[469] <= 19'd0;
		WeightsStore5[470] <= 19'd0;
		WeightsStore5[471] <= 19'd0;
		WeightsStore5[472] <= 19'd0;
		WeightsStore5[473] <= 19'd0;
		WeightsStore5[474] <= 19'd0;
		WeightsStore5[475] <= 19'd0;
		WeightsStore5[476] <= 19'd0;
		WeightsStore5[477] <= 19'd0;
		WeightsStore5[478] <= 19'd0;
		WeightsStore5[479] <= 19'd0;
		WeightsStore5[480] <= 19'd0;
		WeightsStore5[481] <= 19'd0;
		WeightsStore5[482] <= 19'd0;
		WeightsStore5[483] <= 19'd0;
		WeightsStore5[484] <= 19'd0;
		WeightsStore5[485] <= 19'd0;
		WeightsStore5[486] <= 19'd0;
		WeightsStore5[487] <= 19'd0;
		WeightsStore5[488] <= 19'd0;
		WeightsStore5[489] <= 19'd0;
		WeightsStore5[490] <= 19'd0;
		WeightsStore5[491] <= 19'd0;
		WeightsStore5[492] <= 19'd0;
		WeightsStore5[493] <= 19'd0;
		WeightsStore5[494] <= 19'd0;
		WeightsStore5[495] <= 19'd0;
		WeightsStore5[496] <= 19'd0;
		WeightsStore5[497] <= 19'd0;
		WeightsStore5[498] <= 19'd0;
		WeightsStore5[499] <= 19'd0;
		WeightsStore5[500] <= 19'd0;
		WeightsStore5[501] <= 19'd0;
		WeightsStore5[502] <= 19'd0;
		WeightsStore5[503] <= 19'd0;
		WeightsStore5[504] <= 19'd0;
		WeightsStore5[505] <= 19'd0;
		WeightsStore5[506] <= 19'd0;
		WeightsStore5[507] <= 19'd0;
		WeightsStore5[508] <= 19'd0;
		WeightsStore5[509] <= 19'd0;
		WeightsStore5[510] <= 19'd0;
		WeightsStore5[511] <= 19'd0;
		WeightsStore5[512] <= 19'd0;
		WeightsStore5[513] <= 19'd0;
		WeightsStore5[514] <= 19'd0;
		WeightsStore5[515] <= 19'd0;
		WeightsStore5[516] <= 19'd0;
		WeightsStore5[517] <= 19'd0;
		WeightsStore5[518] <= 19'd0;
		WeightsStore5[519] <= 19'd0;
		WeightsStore5[520] <= 19'd0;
		WeightsStore5[521] <= 19'd0;
		WeightsStore5[522] <= 19'd0;
		WeightsStore5[523] <= 19'd0;
		WeightsStore5[524] <= 19'd0;
		WeightsStore5[525] <= 19'd0;
		WeightsStore5[526] <= 19'd0;
		WeightsStore5[527] <= 19'd0;
		WeightsStore5[528] <= 19'd0;
		WeightsStore5[529] <= 19'd0;
		WeightsStore5[530] <= 19'd0;
		WeightsStore5[531] <= 19'd0;
		WeightsStore5[532] <= 19'd0;
		WeightsStore5[533] <= 19'd0;
		WeightsStore5[534] <= 19'd0;
		WeightsStore5[535] <= 19'd0;
		WeightsStore5[536] <= 19'd0;
		WeightsStore5[537] <= 19'd0;
		WeightsStore5[538] <= 19'd0;
		WeightsStore5[539] <= 19'd0;
		WeightsStore5[540] <= 19'd0;
		WeightsStore5[541] <= 19'd0;
		WeightsStore5[542] <= 19'd0;
		WeightsStore5[543] <= 19'd0;
		WeightsStore5[544] <= 19'd0;
		WeightsStore5[545] <= 19'd0;
		WeightsStore5[546] <= 19'd0;
		WeightsStore5[547] <= 19'd0;
		WeightsStore5[548] <= 19'd0;
		WeightsStore5[549] <= 19'd0;
		WeightsStore5[550] <= 19'd0;
		WeightsStore5[551] <= 19'd0;
		WeightsStore5[552] <= 19'd0;
		WeightsStore5[553] <= 19'd0;
		WeightsStore5[554] <= 19'd0;
		WeightsStore5[555] <= 19'd0;
		WeightsStore5[556] <= 19'd0;
		WeightsStore5[557] <= 19'd0;
		WeightsStore5[558] <= 19'd0;
		WeightsStore5[559] <= 19'd0;
		WeightsStore5[560] <= 19'd0;
		WeightsStore5[561] <= 19'd0;
		WeightsStore5[562] <= 19'd0;
		WeightsStore5[563] <= 19'd0;
		WeightsStore5[564] <= 19'd0;
		WeightsStore5[565] <= 19'd0;
		WeightsStore5[566] <= 19'd0;
		WeightsStore5[567] <= 19'd0;
		WeightsStore5[568] <= 19'd0;
		WeightsStore5[569] <= 19'd0;
		WeightsStore5[570] <= 19'd0;
		WeightsStore5[571] <= 19'd0;
		WeightsStore5[572] <= 19'd0;
		WeightsStore5[573] <= 19'd0;
		WeightsStore5[574] <= 19'd0;
		WeightsStore5[575] <= 19'd0;
		WeightsStore5[576] <= 19'd0;
		WeightsStore5[577] <= 19'd0;
		WeightsStore5[578] <= 19'd0;
		WeightsStore5[579] <= 19'd0;
		WeightsStore5[580] <= 19'd0;
		WeightsStore5[581] <= 19'd0;
		WeightsStore5[582] <= 19'd0;
		WeightsStore5[583] <= 19'd0;
		WeightsStore5[584] <= 19'd0;
		WeightsStore5[585] <= 19'd0;
		WeightsStore5[586] <= 19'd0;
		WeightsStore5[587] <= 19'd0;
		WeightsStore5[588] <= 19'd0;
		WeightsStore5[589] <= 19'd0;
		WeightsStore5[590] <= 19'd0;
		WeightsStore5[591] <= 19'd0;
		WeightsStore5[592] <= 19'd0;
		WeightsStore5[593] <= 19'd0;
		WeightsStore5[594] <= 19'd0;
		WeightsStore5[595] <= 19'd0;
		WeightsStore5[596] <= 19'd0;
		WeightsStore5[597] <= 19'd0;
		WeightsStore5[598] <= 19'd0;
		WeightsStore5[599] <= 19'd0;
		WeightsStore5[600] <= 19'd0;
		WeightsStore5[601] <= 19'd0;
		WeightsStore5[602] <= 19'd0;
		WeightsStore5[603] <= 19'd0;
		WeightsStore5[604] <= 19'd0;
		WeightsStore5[605] <= 19'd0;
		WeightsStore5[606] <= 19'd0;
		WeightsStore5[607] <= 19'd0;
		WeightsStore5[608] <= 19'd0;
		WeightsStore5[609] <= 19'd0;
		WeightsStore5[610] <= 19'd0;
		WeightsStore5[611] <= 19'd0;
		WeightsStore5[612] <= 19'd0;
		WeightsStore5[613] <= 19'd0;
		WeightsStore5[614] <= 19'd0;
		WeightsStore5[615] <= 19'd0;
		WeightsStore5[616] <= 19'd0;
		WeightsStore5[617] <= 19'd0;
		WeightsStore5[618] <= 19'd0;
		WeightsStore5[619] <= 19'd0;
		WeightsStore5[620] <= 19'd0;
		WeightsStore5[621] <= 19'd0;
		WeightsStore5[622] <= 19'd0;
		WeightsStore5[623] <= 19'd0;
		WeightsStore5[624] <= 19'd0;
		WeightsStore5[625] <= 19'd0;
		WeightsStore5[626] <= 19'd0;
		WeightsStore5[627] <= 19'd0;
		WeightsStore5[628] <= 19'd0;
		WeightsStore5[629] <= 19'd0;
		WeightsStore5[630] <= 19'd0;
		WeightsStore5[631] <= 19'd0;
		WeightsStore5[632] <= 19'd0;
		WeightsStore5[633] <= 19'd0;
		WeightsStore5[634] <= 19'd0;
		WeightsStore5[635] <= 19'd0;
		WeightsStore5[636] <= 19'd0;
		WeightsStore5[637] <= 19'd0;
		WeightsStore5[638] <= 19'd0;
		WeightsStore5[639] <= 19'd0;
		WeightsStore5[640] <= 19'd0;
		WeightsStore5[641] <= 19'd0;
		WeightsStore5[642] <= 19'd0;
		WeightsStore5[643] <= 19'd0;
		WeightsStore5[644] <= 19'd0;
		WeightsStore5[645] <= 19'd0;
		WeightsStore5[646] <= 19'd0;
		WeightsStore5[647] <= 19'd0;
		WeightsStore5[648] <= 19'd0;
		WeightsStore5[649] <= 19'd0;
		WeightsStore5[650] <= 19'd0;
		WeightsStore5[651] <= 19'd0;
		WeightsStore5[652] <= 19'd0;
		WeightsStore5[653] <= 19'd0;
		WeightsStore5[654] <= 19'd0;
		WeightsStore5[655] <= 19'd0;
		WeightsStore5[656] <= 19'd0;
		WeightsStore5[657] <= 19'd0;
		WeightsStore5[658] <= 19'd0;
		WeightsStore5[659] <= 19'd0;
		WeightsStore5[660] <= 19'd0;
		WeightsStore5[661] <= 19'd0;
		WeightsStore5[662] <= 19'd0;
		WeightsStore5[663] <= 19'd0;
		WeightsStore5[664] <= 19'd0;
		WeightsStore5[665] <= 19'd0;
		WeightsStore5[666] <= 19'd0;
		WeightsStore5[667] <= 19'd0;
		WeightsStore5[668] <= 19'd0;
		WeightsStore5[669] <= 19'd0;
		WeightsStore5[670] <= 19'd0;
		WeightsStore5[671] <= 19'd0;
		WeightsStore5[672] <= 19'd0;
		WeightsStore5[673] <= 19'd0;
		WeightsStore5[674] <= 19'd0;
		WeightsStore5[675] <= 19'd0;
		WeightsStore5[676] <= 19'd0;
		WeightsStore5[677] <= 19'd0;
		WeightsStore5[678] <= 19'd0;
		WeightsStore5[679] <= 19'd0;
		WeightsStore5[680] <= 19'd0;
		WeightsStore5[681] <= 19'd0;
		WeightsStore5[682] <= 19'd0;
		WeightsStore5[683] <= 19'd0;
		WeightsStore5[684] <= 19'd0;
		WeightsStore5[685] <= 19'd0;
		WeightsStore5[686] <= 19'd0;
		WeightsStore5[687] <= 19'd0;
		WeightsStore5[688] <= 19'd0;
		WeightsStore5[689] <= 19'd0;
		WeightsStore5[690] <= 19'd0;
		WeightsStore5[691] <= 19'd0;
		WeightsStore5[692] <= 19'd0;
		WeightsStore5[693] <= 19'd0;
		WeightsStore5[694] <= 19'd0;
		WeightsStore5[695] <= 19'd0;
		WeightsStore5[696] <= 19'd0;
		WeightsStore5[697] <= 19'd0;
		WeightsStore5[698] <= 19'd0;
		WeightsStore5[699] <= 19'd0;
		WeightsStore5[700] <= 19'd0;
		WeightsStore5[701] <= 19'd0;
		WeightsStore5[702] <= 19'd0;
		WeightsStore5[703] <= 19'd0;
		WeightsStore5[704] <= 19'd0;
		WeightsStore5[705] <= 19'd0;
		WeightsStore5[706] <= 19'd0;
		WeightsStore5[707] <= 19'd0;
		WeightsStore5[708] <= 19'd0;
		WeightsStore5[709] <= 19'd0;
		WeightsStore5[710] <= 19'd0;
		WeightsStore5[711] <= 19'd0;
		WeightsStore5[712] <= 19'd0;
		WeightsStore5[713] <= 19'd0;
		WeightsStore5[714] <= 19'd0;
		WeightsStore5[715] <= 19'd0;
		WeightsStore5[716] <= 19'd0;
		WeightsStore5[717] <= 19'd0;
		WeightsStore5[718] <= 19'd0;
		WeightsStore5[719] <= 19'd0;
		WeightsStore5[720] <= 19'd0;
		WeightsStore5[721] <= 19'd0;
		WeightsStore5[722] <= 19'd0;
		WeightsStore5[723] <= 19'd0;
		WeightsStore5[724] <= 19'd0;
		WeightsStore5[725] <= 19'd0;
		WeightsStore5[726] <= 19'd0;
		WeightsStore5[727] <= 19'd0;
		WeightsStore5[728] <= 19'd0;
		WeightsStore5[729] <= 19'd0;
		WeightsStore5[730] <= 19'd0;
		WeightsStore5[731] <= 19'd0;
		WeightsStore5[732] <= 19'd0;
		WeightsStore5[733] <= 19'd0;
		WeightsStore5[734] <= 19'd0;
		WeightsStore5[735] <= 19'd0;
		WeightsStore5[736] <= 19'd0;
		WeightsStore5[737] <= 19'd0;
		WeightsStore5[738] <= 19'd0;
		WeightsStore5[739] <= 19'd0;
		WeightsStore5[740] <= 19'd0;
		WeightsStore5[741] <= 19'd0;
		WeightsStore5[742] <= 19'd0;
		WeightsStore5[743] <= 19'd0;
		WeightsStore5[744] <= 19'd0;
		WeightsStore5[745] <= 19'd0;
		WeightsStore5[746] <= 19'd0;
		WeightsStore5[747] <= 19'd0;
		WeightsStore5[748] <= 19'd0;
		WeightsStore5[749] <= 19'd0;
		WeightsStore5[750] <= 19'd0;
		WeightsStore5[751] <= 19'd0;
		WeightsStore5[752] <= 19'd0;
		WeightsStore5[753] <= 19'd0;
		WeightsStore5[754] <= 19'd0;
		WeightsStore5[755] <= 19'd0;
		WeightsStore5[756] <= 19'd0;
		WeightsStore5[757] <= 19'd0;
		WeightsStore5[758] <= 19'd0;
		WeightsStore5[759] <= 19'd0;
		WeightsStore5[760] <= 19'd0;
		WeightsStore5[761] <= 19'd0;
		WeightsStore5[762] <= 19'd0;
		WeightsStore5[763] <= 19'd0;
		WeightsStore5[764] <= 19'd0;
		WeightsStore5[765] <= 19'd0;
		WeightsStore5[766] <= 19'd0;
		WeightsStore5[767] <= 19'd0;
		WeightsStore5[768] <= 19'd0;
		WeightsStore5[769] <= 19'd0;
		WeightsStore5[770] <= 19'd0;
		WeightsStore5[771] <= 19'd0;
		WeightsStore5[772] <= 19'd0;
		WeightsStore5[773] <= 19'd0;
		WeightsStore5[774] <= 19'd0;
		WeightsStore5[775] <= 19'd0;
		WeightsStore5[776] <= 19'd0;
		WeightsStore5[777] <= 19'd0;
		WeightsStore5[778] <= 19'd0;
		WeightsStore5[779] <= 19'd0;
		WeightsStore5[780] <= 19'd0;
		WeightsStore5[781] <= 19'd0;
		WeightsStore5[782] <= 19'd0;
		WeightsStore5[783] <= 19'd0;
		WeightsStore5[784] <= 19'd0;
		WeightsStore6[0] <= 19'd0;
		WeightsStore6[1] <= 19'd0;
		WeightsStore6[2] <= 19'd0;
		WeightsStore6[3] <= 19'd0;
		WeightsStore6[4] <= 19'd0;
		WeightsStore6[5] <= 19'd0;
		WeightsStore6[6] <= 19'd0;
		WeightsStore6[7] <= 19'd0;
		WeightsStore6[8] <= 19'd0;
		WeightsStore6[9] <= 19'd0;
		WeightsStore6[10] <= 19'd0;
		WeightsStore6[11] <= 19'd0;
		WeightsStore6[12] <= 19'd0;
		WeightsStore6[13] <= 19'd0;
		WeightsStore6[14] <= 19'd0;
		WeightsStore6[15] <= 19'd0;
		WeightsStore6[16] <= 19'd0;
		WeightsStore6[17] <= 19'd0;
		WeightsStore6[18] <= 19'd0;
		WeightsStore6[19] <= 19'd0;
		WeightsStore6[20] <= 19'd0;
		WeightsStore6[21] <= 19'd0;
		WeightsStore6[22] <= 19'd0;
		WeightsStore6[23] <= 19'd0;
		WeightsStore6[24] <= 19'd0;
		WeightsStore6[25] <= 19'd0;
		WeightsStore6[26] <= 19'd0;
		WeightsStore6[27] <= 19'd0;
		WeightsStore6[28] <= 19'd0;
		WeightsStore6[29] <= 19'd0;
		WeightsStore6[30] <= 19'd0;
		WeightsStore6[31] <= 19'd0;
		WeightsStore6[32] <= 19'd0;
		WeightsStore6[33] <= 19'd0;
		WeightsStore6[34] <= 19'd0;
		WeightsStore6[35] <= 19'd0;
		WeightsStore6[36] <= 19'd0;
		WeightsStore6[37] <= 19'd0;
		WeightsStore6[38] <= 19'd0;
		WeightsStore6[39] <= 19'd0;
		WeightsStore6[40] <= 19'd0;
		WeightsStore6[41] <= 19'd0;
		WeightsStore6[42] <= 19'd0;
		WeightsStore6[43] <= 19'd0;
		WeightsStore6[44] <= 19'd0;
		WeightsStore6[45] <= 19'd0;
		WeightsStore6[46] <= 19'd0;
		WeightsStore6[47] <= 19'd0;
		WeightsStore6[48] <= 19'd0;
		WeightsStore6[49] <= 19'd0;
		WeightsStore6[50] <= 19'd0;
		WeightsStore6[51] <= 19'd0;
		WeightsStore6[52] <= 19'd0;
		WeightsStore6[53] <= 19'd0;
		WeightsStore6[54] <= 19'd0;
		WeightsStore6[55] <= 19'd0;
		WeightsStore6[56] <= 19'd0;
		WeightsStore6[57] <= 19'd0;
		WeightsStore6[58] <= 19'd0;
		WeightsStore6[59] <= 19'd0;
		WeightsStore6[60] <= 19'd0;
		WeightsStore6[61] <= 19'd0;
		WeightsStore6[62] <= 19'd0;
		WeightsStore6[63] <= 19'd0;
		WeightsStore6[64] <= 19'd0;
		WeightsStore6[65] <= 19'd0;
		WeightsStore6[66] <= 19'd0;
		WeightsStore6[67] <= 19'd0;
		WeightsStore6[68] <= 19'd0;
		WeightsStore6[69] <= 19'd0;
		WeightsStore6[70] <= 19'd0;
		WeightsStore6[71] <= 19'd0;
		WeightsStore6[72] <= 19'd0;
		WeightsStore6[73] <= 19'd0;
		WeightsStore6[74] <= 19'd0;
		WeightsStore6[75] <= 19'd0;
		WeightsStore6[76] <= 19'd0;
		WeightsStore6[77] <= 19'd0;
		WeightsStore6[78] <= 19'd0;
		WeightsStore6[79] <= 19'd0;
		WeightsStore6[80] <= 19'd0;
		WeightsStore6[81] <= 19'd0;
		WeightsStore6[82] <= 19'd0;
		WeightsStore6[83] <= 19'd0;
		WeightsStore6[84] <= 19'd0;
		WeightsStore6[85] <= 19'd0;
		WeightsStore6[86] <= 19'd0;
		WeightsStore6[87] <= 19'd0;
		WeightsStore6[88] <= 19'd0;
		WeightsStore6[89] <= 19'd0;
		WeightsStore6[90] <= 19'd0;
		WeightsStore6[91] <= 19'd0;
		WeightsStore6[92] <= 19'd0;
		WeightsStore6[93] <= 19'd0;
		WeightsStore6[94] <= 19'd0;
		WeightsStore6[95] <= 19'd0;
		WeightsStore6[96] <= 19'd0;
		WeightsStore6[97] <= 19'd0;
		WeightsStore6[98] <= 19'd0;
		WeightsStore6[99] <= 19'd0;
		WeightsStore6[100] <= 19'd0;
		WeightsStore6[101] <= 19'd0;
		WeightsStore6[102] <= 19'd0;
		WeightsStore6[103] <= 19'd0;
		WeightsStore6[104] <= 19'd0;
		WeightsStore6[105] <= 19'd0;
		WeightsStore6[106] <= 19'd0;
		WeightsStore6[107] <= 19'd0;
		WeightsStore6[108] <= 19'd0;
		WeightsStore6[109] <= 19'd0;
		WeightsStore6[110] <= 19'd0;
		WeightsStore6[111] <= 19'd0;
		WeightsStore6[112] <= 19'd0;
		WeightsStore6[113] <= 19'd0;
		WeightsStore6[114] <= 19'd0;
		WeightsStore6[115] <= 19'd0;
		WeightsStore6[116] <= 19'd0;
		WeightsStore6[117] <= 19'd0;
		WeightsStore6[118] <= 19'd0;
		WeightsStore6[119] <= 19'd0;
		WeightsStore6[120] <= 19'd0;
		WeightsStore6[121] <= 19'd0;
		WeightsStore6[122] <= 19'd0;
		WeightsStore6[123] <= 19'd0;
		WeightsStore6[124] <= 19'd0;
		WeightsStore6[125] <= 19'd0;
		WeightsStore6[126] <= 19'd0;
		WeightsStore6[127] <= 19'd0;
		WeightsStore6[128] <= 19'd0;
		WeightsStore6[129] <= 19'd0;
		WeightsStore6[130] <= 19'd0;
		WeightsStore6[131] <= 19'd0;
		WeightsStore6[132] <= 19'd0;
		WeightsStore6[133] <= 19'd0;
		WeightsStore6[134] <= 19'd0;
		WeightsStore6[135] <= 19'd0;
		WeightsStore6[136] <= 19'd0;
		WeightsStore6[137] <= 19'd0;
		WeightsStore6[138] <= 19'd0;
		WeightsStore6[139] <= 19'd0;
		WeightsStore6[140] <= 19'd0;
		WeightsStore6[141] <= 19'd0;
		WeightsStore6[142] <= 19'd0;
		WeightsStore6[143] <= 19'd0;
		WeightsStore6[144] <= 19'd0;
		WeightsStore6[145] <= 19'd0;
		WeightsStore6[146] <= 19'd0;
		WeightsStore6[147] <= 19'd0;
		WeightsStore6[148] <= 19'd0;
		WeightsStore6[149] <= 19'd0;
		WeightsStore6[150] <= 19'd0;
		WeightsStore6[151] <= 19'd0;
		WeightsStore6[152] <= 19'd0;
		WeightsStore6[153] <= 19'd0;
		WeightsStore6[154] <= 19'd0;
		WeightsStore6[155] <= 19'd0;
		WeightsStore6[156] <= 19'd0;
		WeightsStore6[157] <= 19'd0;
		WeightsStore6[158] <= 19'd0;
		WeightsStore6[159] <= 19'd0;
		WeightsStore6[160] <= 19'd0;
		WeightsStore6[161] <= 19'd0;
		WeightsStore6[162] <= 19'd0;
		WeightsStore6[163] <= 19'd0;
		WeightsStore6[164] <= 19'd0;
		WeightsStore6[165] <= 19'd0;
		WeightsStore6[166] <= 19'd0;
		WeightsStore6[167] <= 19'd0;
		WeightsStore6[168] <= 19'd0;
		WeightsStore6[169] <= 19'd0;
		WeightsStore6[170] <= 19'd0;
		WeightsStore6[171] <= 19'd0;
		WeightsStore6[172] <= 19'd0;
		WeightsStore6[173] <= 19'd0;
		WeightsStore6[174] <= 19'd0;
		WeightsStore6[175] <= 19'd0;
		WeightsStore6[176] <= 19'd0;
		WeightsStore6[177] <= 19'd0;
		WeightsStore6[178] <= 19'd0;
		WeightsStore6[179] <= 19'd0;
		WeightsStore6[180] <= 19'd0;
		WeightsStore6[181] <= 19'd0;
		WeightsStore6[182] <= 19'd0;
		WeightsStore6[183] <= 19'd0;
		WeightsStore6[184] <= 19'd0;
		WeightsStore6[185] <= 19'd0;
		WeightsStore6[186] <= 19'd0;
		WeightsStore6[187] <= 19'd0;
		WeightsStore6[188] <= 19'd0;
		WeightsStore6[189] <= 19'd0;
		WeightsStore6[190] <= 19'd0;
		WeightsStore6[191] <= 19'd0;
		WeightsStore6[192] <= 19'd0;
		WeightsStore6[193] <= 19'd0;
		WeightsStore6[194] <= 19'd0;
		WeightsStore6[195] <= 19'd0;
		WeightsStore6[196] <= 19'd0;
		WeightsStore6[197] <= 19'd0;
		WeightsStore6[198] <= 19'd0;
		WeightsStore6[199] <= 19'd0;
		WeightsStore6[200] <= 19'd0;
		WeightsStore6[201] <= 19'd0;
		WeightsStore6[202] <= 19'd0;
		WeightsStore6[203] <= 19'd0;
		WeightsStore6[204] <= 19'd0;
		WeightsStore6[205] <= 19'd0;
		WeightsStore6[206] <= 19'd0;
		WeightsStore6[207] <= 19'd0;
		WeightsStore6[208] <= 19'd0;
		WeightsStore6[209] <= 19'd0;
		WeightsStore6[210] <= 19'd0;
		WeightsStore6[211] <= 19'd0;
		WeightsStore6[212] <= 19'd0;
		WeightsStore6[213] <= 19'd0;
		WeightsStore6[214] <= 19'd0;
		WeightsStore6[215] <= 19'd0;
		WeightsStore6[216] <= 19'd0;
		WeightsStore6[217] <= 19'd0;
		WeightsStore6[218] <= 19'd0;
		WeightsStore6[219] <= 19'd0;
		WeightsStore6[220] <= 19'd0;
		WeightsStore6[221] <= 19'd0;
		WeightsStore6[222] <= 19'd0;
		WeightsStore6[223] <= 19'd0;
		WeightsStore6[224] <= 19'd0;
		WeightsStore6[225] <= 19'd0;
		WeightsStore6[226] <= 19'd0;
		WeightsStore6[227] <= 19'd0;
		WeightsStore6[228] <= 19'd0;
		WeightsStore6[229] <= 19'd0;
		WeightsStore6[230] <= 19'd0;
		WeightsStore6[231] <= 19'd0;
		WeightsStore6[232] <= 19'd0;
		WeightsStore6[233] <= 19'd0;
		WeightsStore6[234] <= 19'd0;
		WeightsStore6[235] <= 19'd0;
		WeightsStore6[236] <= 19'd0;
		WeightsStore6[237] <= 19'd0;
		WeightsStore6[238] <= 19'd0;
		WeightsStore6[239] <= 19'd0;
		WeightsStore6[240] <= 19'd0;
		WeightsStore6[241] <= 19'd0;
		WeightsStore6[242] <= 19'd0;
		WeightsStore6[243] <= 19'd0;
		WeightsStore6[244] <= 19'd0;
		WeightsStore6[245] <= 19'd0;
		WeightsStore6[246] <= 19'd0;
		WeightsStore6[247] <= 19'd0;
		WeightsStore6[248] <= 19'd0;
		WeightsStore6[249] <= 19'd0;
		WeightsStore6[250] <= 19'd0;
		WeightsStore6[251] <= 19'd0;
		WeightsStore6[252] <= 19'd0;
		WeightsStore6[253] <= 19'd0;
		WeightsStore6[254] <= 19'd0;
		WeightsStore6[255] <= 19'd0;
		WeightsStore6[256] <= 19'd0;
		WeightsStore6[257] <= 19'd0;
		WeightsStore6[258] <= 19'd0;
		WeightsStore6[259] <= 19'd0;
		WeightsStore6[260] <= 19'd0;
		WeightsStore6[261] <= 19'd0;
		WeightsStore6[262] <= 19'd0;
		WeightsStore6[263] <= 19'd0;
		WeightsStore6[264] <= 19'd0;
		WeightsStore6[265] <= 19'd0;
		WeightsStore6[266] <= 19'd0;
		WeightsStore6[267] <= 19'd0;
		WeightsStore6[268] <= 19'd0;
		WeightsStore6[269] <= 19'd0;
		WeightsStore6[270] <= 19'd0;
		WeightsStore6[271] <= 19'd0;
		WeightsStore6[272] <= 19'd0;
		WeightsStore6[273] <= 19'd0;
		WeightsStore6[274] <= 19'd0;
		WeightsStore6[275] <= 19'd0;
		WeightsStore6[276] <= 19'd0;
		WeightsStore6[277] <= 19'd0;
		WeightsStore6[278] <= 19'd0;
		WeightsStore6[279] <= 19'd0;
		WeightsStore6[280] <= 19'd0;
		WeightsStore6[281] <= 19'd0;
		WeightsStore6[282] <= 19'd0;
		WeightsStore6[283] <= 19'd0;
		WeightsStore6[284] <= 19'd0;
		WeightsStore6[285] <= 19'd0;
		WeightsStore6[286] <= 19'd0;
		WeightsStore6[287] <= 19'd0;
		WeightsStore6[288] <= 19'd0;
		WeightsStore6[289] <= 19'd0;
		WeightsStore6[290] <= 19'd0;
		WeightsStore6[291] <= 19'd0;
		WeightsStore6[292] <= 19'd0;
		WeightsStore6[293] <= 19'd0;
		WeightsStore6[294] <= 19'd0;
		WeightsStore6[295] <= 19'd0;
		WeightsStore6[296] <= 19'd0;
		WeightsStore6[297] <= 19'd0;
		WeightsStore6[298] <= 19'd0;
		WeightsStore6[299] <= 19'd0;
		WeightsStore6[300] <= 19'd0;
		WeightsStore6[301] <= 19'd0;
		WeightsStore6[302] <= 19'd0;
		WeightsStore6[303] <= 19'd0;
		WeightsStore6[304] <= 19'd0;
		WeightsStore6[305] <= 19'd0;
		WeightsStore6[306] <= 19'd0;
		WeightsStore6[307] <= 19'd0;
		WeightsStore6[308] <= 19'd0;
		WeightsStore6[309] <= 19'd0;
		WeightsStore6[310] <= 19'd0;
		WeightsStore6[311] <= 19'd0;
		WeightsStore6[312] <= 19'd0;
		WeightsStore6[313] <= 19'd0;
		WeightsStore6[314] <= 19'd0;
		WeightsStore6[315] <= 19'd0;
		WeightsStore6[316] <= 19'd0;
		WeightsStore6[317] <= 19'd0;
		WeightsStore6[318] <= 19'd0;
		WeightsStore6[319] <= 19'd0;
		WeightsStore6[320] <= 19'd0;
		WeightsStore6[321] <= 19'd0;
		WeightsStore6[322] <= 19'd0;
		WeightsStore6[323] <= 19'd0;
		WeightsStore6[324] <= 19'd0;
		WeightsStore6[325] <= 19'd0;
		WeightsStore6[326] <= 19'd0;
		WeightsStore6[327] <= 19'd0;
		WeightsStore6[328] <= 19'd0;
		WeightsStore6[329] <= 19'd0;
		WeightsStore6[330] <= 19'd0;
		WeightsStore6[331] <= 19'd0;
		WeightsStore6[332] <= 19'd0;
		WeightsStore6[333] <= 19'd0;
		WeightsStore6[334] <= 19'd0;
		WeightsStore6[335] <= 19'd0;
		WeightsStore6[336] <= 19'd0;
		WeightsStore6[337] <= 19'd0;
		WeightsStore6[338] <= 19'd0;
		WeightsStore6[339] <= 19'd0;
		WeightsStore6[340] <= 19'd0;
		WeightsStore6[341] <= 19'd0;
		WeightsStore6[342] <= 19'd0;
		WeightsStore6[343] <= 19'd0;
		WeightsStore6[344] <= 19'd0;
		WeightsStore6[345] <= 19'd0;
		WeightsStore6[346] <= 19'd0;
		WeightsStore6[347] <= 19'd0;
		WeightsStore6[348] <= 19'd0;
		WeightsStore6[349] <= 19'd0;
		WeightsStore6[350] <= 19'd0;
		WeightsStore6[351] <= 19'd0;
		WeightsStore6[352] <= 19'd0;
		WeightsStore6[353] <= 19'd0;
		WeightsStore6[354] <= 19'd0;
		WeightsStore6[355] <= 19'd0;
		WeightsStore6[356] <= 19'd0;
		WeightsStore6[357] <= 19'd0;
		WeightsStore6[358] <= 19'd0;
		WeightsStore6[359] <= 19'd0;
		WeightsStore6[360] <= 19'd0;
		WeightsStore6[361] <= 19'd0;
		WeightsStore6[362] <= 19'd0;
		WeightsStore6[363] <= 19'd0;
		WeightsStore6[364] <= 19'd0;
		WeightsStore6[365] <= 19'd0;
		WeightsStore6[366] <= 19'd0;
		WeightsStore6[367] <= 19'd0;
		WeightsStore6[368] <= 19'd0;
		WeightsStore6[369] <= 19'd0;
		WeightsStore6[370] <= 19'd0;
		WeightsStore6[371] <= 19'd0;
		WeightsStore6[372] <= 19'd0;
		WeightsStore6[373] <= 19'd0;
		WeightsStore6[374] <= 19'd0;
		WeightsStore6[375] <= 19'd0;
		WeightsStore6[376] <= 19'd0;
		WeightsStore6[377] <= 19'd0;
		WeightsStore6[378] <= 19'd0;
		WeightsStore6[379] <= 19'd0;
		WeightsStore6[380] <= 19'd0;
		WeightsStore6[381] <= 19'd0;
		WeightsStore6[382] <= 19'd0;
		WeightsStore6[383] <= 19'd0;
		WeightsStore6[384] <= 19'd0;
		WeightsStore6[385] <= 19'd0;
		WeightsStore6[386] <= 19'd0;
		WeightsStore6[387] <= 19'd0;
		WeightsStore6[388] <= 19'd0;
		WeightsStore6[389] <= 19'd0;
		WeightsStore6[390] <= 19'd0;
		WeightsStore6[391] <= 19'd0;
		WeightsStore6[392] <= 19'd0;
		WeightsStore6[393] <= 19'd0;
		WeightsStore6[394] <= 19'd0;
		WeightsStore6[395] <= 19'd0;
		WeightsStore6[396] <= 19'd0;
		WeightsStore6[397] <= 19'd0;
		WeightsStore6[398] <= 19'd0;
		WeightsStore6[399] <= 19'd0;
		WeightsStore6[400] <= 19'd0;
		WeightsStore6[401] <= 19'd0;
		WeightsStore6[402] <= 19'd0;
		WeightsStore6[403] <= 19'd0;
		WeightsStore6[404] <= 19'd0;
		WeightsStore6[405] <= 19'd0;
		WeightsStore6[406] <= 19'd0;
		WeightsStore6[407] <= 19'd0;
		WeightsStore6[408] <= 19'd0;
		WeightsStore6[409] <= 19'd0;
		WeightsStore6[410] <= 19'd0;
		WeightsStore6[411] <= 19'd0;
		WeightsStore6[412] <= 19'd0;
		WeightsStore6[413] <= 19'd0;
		WeightsStore6[414] <= 19'd0;
		WeightsStore6[415] <= 19'd0;
		WeightsStore6[416] <= 19'd0;
		WeightsStore6[417] <= 19'd0;
		WeightsStore6[418] <= 19'd0;
		WeightsStore6[419] <= 19'd0;
		WeightsStore6[420] <= 19'd0;
		WeightsStore6[421] <= 19'd0;
		WeightsStore6[422] <= 19'd0;
		WeightsStore6[423] <= 19'd0;
		WeightsStore6[424] <= 19'd0;
		WeightsStore6[425] <= 19'd0;
		WeightsStore6[426] <= 19'd0;
		WeightsStore6[427] <= 19'd0;
		WeightsStore6[428] <= 19'd0;
		WeightsStore6[429] <= 19'd0;
		WeightsStore6[430] <= 19'd0;
		WeightsStore6[431] <= 19'd0;
		WeightsStore6[432] <= 19'd0;
		WeightsStore6[433] <= 19'd0;
		WeightsStore6[434] <= 19'd0;
		WeightsStore6[435] <= 19'd0;
		WeightsStore6[436] <= 19'd0;
		WeightsStore6[437] <= 19'd0;
		WeightsStore6[438] <= 19'd0;
		WeightsStore6[439] <= 19'd0;
		WeightsStore6[440] <= 19'd0;
		WeightsStore6[441] <= 19'd0;
		WeightsStore6[442] <= 19'd0;
		WeightsStore6[443] <= 19'd0;
		WeightsStore6[444] <= 19'd0;
		WeightsStore6[445] <= 19'd0;
		WeightsStore6[446] <= 19'd0;
		WeightsStore6[447] <= 19'd0;
		WeightsStore6[448] <= 19'd0;
		WeightsStore6[449] <= 19'd0;
		WeightsStore6[450] <= 19'd0;
		WeightsStore6[451] <= 19'd0;
		WeightsStore6[452] <= 19'd0;
		WeightsStore6[453] <= 19'd0;
		WeightsStore6[454] <= 19'd0;
		WeightsStore6[455] <= 19'd0;
		WeightsStore6[456] <= 19'd0;
		WeightsStore6[457] <= 19'd0;
		WeightsStore6[458] <= 19'd0;
		WeightsStore6[459] <= 19'd0;
		WeightsStore6[460] <= 19'd0;
		WeightsStore6[461] <= 19'd0;
		WeightsStore6[462] <= 19'd0;
		WeightsStore6[463] <= 19'd0;
		WeightsStore6[464] <= 19'd0;
		WeightsStore6[465] <= 19'd0;
		WeightsStore6[466] <= 19'd0;
		WeightsStore6[467] <= 19'd0;
		WeightsStore6[468] <= 19'd0;
		WeightsStore6[469] <= 19'd0;
		WeightsStore6[470] <= 19'd0;
		WeightsStore6[471] <= 19'd0;
		WeightsStore6[472] <= 19'd0;
		WeightsStore6[473] <= 19'd0;
		WeightsStore6[474] <= 19'd0;
		WeightsStore6[475] <= 19'd0;
		WeightsStore6[476] <= 19'd0;
		WeightsStore6[477] <= 19'd0;
		WeightsStore6[478] <= 19'd0;
		WeightsStore6[479] <= 19'd0;
		WeightsStore6[480] <= 19'd0;
		WeightsStore6[481] <= 19'd0;
		WeightsStore6[482] <= 19'd0;
		WeightsStore6[483] <= 19'd0;
		WeightsStore6[484] <= 19'd0;
		WeightsStore6[485] <= 19'd0;
		WeightsStore6[486] <= 19'd0;
		WeightsStore6[487] <= 19'd0;
		WeightsStore6[488] <= 19'd0;
		WeightsStore6[489] <= 19'd0;
		WeightsStore6[490] <= 19'd0;
		WeightsStore6[491] <= 19'd0;
		WeightsStore6[492] <= 19'd0;
		WeightsStore6[493] <= 19'd0;
		WeightsStore6[494] <= 19'd0;
		WeightsStore6[495] <= 19'd0;
		WeightsStore6[496] <= 19'd0;
		WeightsStore6[497] <= 19'd0;
		WeightsStore6[498] <= 19'd0;
		WeightsStore6[499] <= 19'd0;
		WeightsStore6[500] <= 19'd0;
		WeightsStore6[501] <= 19'd0;
		WeightsStore6[502] <= 19'd0;
		WeightsStore6[503] <= 19'd0;
		WeightsStore6[504] <= 19'd0;
		WeightsStore6[505] <= 19'd0;
		WeightsStore6[506] <= 19'd0;
		WeightsStore6[507] <= 19'd0;
		WeightsStore6[508] <= 19'd0;
		WeightsStore6[509] <= 19'd0;
		WeightsStore6[510] <= 19'd0;
		WeightsStore6[511] <= 19'd0;
		WeightsStore6[512] <= 19'd0;
		WeightsStore6[513] <= 19'd0;
		WeightsStore6[514] <= 19'd0;
		WeightsStore6[515] <= 19'd0;
		WeightsStore6[516] <= 19'd0;
		WeightsStore6[517] <= 19'd0;
		WeightsStore6[518] <= 19'd0;
		WeightsStore6[519] <= 19'd0;
		WeightsStore6[520] <= 19'd0;
		WeightsStore6[521] <= 19'd0;
		WeightsStore6[522] <= 19'd0;
		WeightsStore6[523] <= 19'd0;
		WeightsStore6[524] <= 19'd0;
		WeightsStore6[525] <= 19'd0;
		WeightsStore6[526] <= 19'd0;
		WeightsStore6[527] <= 19'd0;
		WeightsStore6[528] <= 19'd0;
		WeightsStore6[529] <= 19'd0;
		WeightsStore6[530] <= 19'd0;
		WeightsStore6[531] <= 19'd0;
		WeightsStore6[532] <= 19'd0;
		WeightsStore6[533] <= 19'd0;
		WeightsStore6[534] <= 19'd0;
		WeightsStore6[535] <= 19'd0;
		WeightsStore6[536] <= 19'd0;
		WeightsStore6[537] <= 19'd0;
		WeightsStore6[538] <= 19'd0;
		WeightsStore6[539] <= 19'd0;
		WeightsStore6[540] <= 19'd0;
		WeightsStore6[541] <= 19'd0;
		WeightsStore6[542] <= 19'd0;
		WeightsStore6[543] <= 19'd0;
		WeightsStore6[544] <= 19'd0;
		WeightsStore6[545] <= 19'd0;
		WeightsStore6[546] <= 19'd0;
		WeightsStore6[547] <= 19'd0;
		WeightsStore6[548] <= 19'd0;
		WeightsStore6[549] <= 19'd0;
		WeightsStore6[550] <= 19'd0;
		WeightsStore6[551] <= 19'd0;
		WeightsStore6[552] <= 19'd0;
		WeightsStore6[553] <= 19'd0;
		WeightsStore6[554] <= 19'd0;
		WeightsStore6[555] <= 19'd0;
		WeightsStore6[556] <= 19'd0;
		WeightsStore6[557] <= 19'd0;
		WeightsStore6[558] <= 19'd0;
		WeightsStore6[559] <= 19'd0;
		WeightsStore6[560] <= 19'd0;
		WeightsStore6[561] <= 19'd0;
		WeightsStore6[562] <= 19'd0;
		WeightsStore6[563] <= 19'd0;
		WeightsStore6[564] <= 19'd0;
		WeightsStore6[565] <= 19'd0;
		WeightsStore6[566] <= 19'd0;
		WeightsStore6[567] <= 19'd0;
		WeightsStore6[568] <= 19'd0;
		WeightsStore6[569] <= 19'd0;
		WeightsStore6[570] <= 19'd0;
		WeightsStore6[571] <= 19'd0;
		WeightsStore6[572] <= 19'd0;
		WeightsStore6[573] <= 19'd0;
		WeightsStore6[574] <= 19'd0;
		WeightsStore6[575] <= 19'd0;
		WeightsStore6[576] <= 19'd0;
		WeightsStore6[577] <= 19'd0;
		WeightsStore6[578] <= 19'd0;
		WeightsStore6[579] <= 19'd0;
		WeightsStore6[580] <= 19'd0;
		WeightsStore6[581] <= 19'd0;
		WeightsStore6[582] <= 19'd0;
		WeightsStore6[583] <= 19'd0;
		WeightsStore6[584] <= 19'd0;
		WeightsStore6[585] <= 19'd0;
		WeightsStore6[586] <= 19'd0;
		WeightsStore6[587] <= 19'd0;
		WeightsStore6[588] <= 19'd0;
		WeightsStore6[589] <= 19'd0;
		WeightsStore6[590] <= 19'd0;
		WeightsStore6[591] <= 19'd0;
		WeightsStore6[592] <= 19'd0;
		WeightsStore6[593] <= 19'd0;
		WeightsStore6[594] <= 19'd0;
		WeightsStore6[595] <= 19'd0;
		WeightsStore6[596] <= 19'd0;
		WeightsStore6[597] <= 19'd0;
		WeightsStore6[598] <= 19'd0;
		WeightsStore6[599] <= 19'd0;
		WeightsStore6[600] <= 19'd0;
		WeightsStore6[601] <= 19'd0;
		WeightsStore6[602] <= 19'd0;
		WeightsStore6[603] <= 19'd0;
		WeightsStore6[604] <= 19'd0;
		WeightsStore6[605] <= 19'd0;
		WeightsStore6[606] <= 19'd0;
		WeightsStore6[607] <= 19'd0;
		WeightsStore6[608] <= 19'd0;
		WeightsStore6[609] <= 19'd0;
		WeightsStore6[610] <= 19'd0;
		WeightsStore6[611] <= 19'd0;
		WeightsStore6[612] <= 19'd0;
		WeightsStore6[613] <= 19'd0;
		WeightsStore6[614] <= 19'd0;
		WeightsStore6[615] <= 19'd0;
		WeightsStore6[616] <= 19'd0;
		WeightsStore6[617] <= 19'd0;
		WeightsStore6[618] <= 19'd0;
		WeightsStore6[619] <= 19'd0;
		WeightsStore6[620] <= 19'd0;
		WeightsStore6[621] <= 19'd0;
		WeightsStore6[622] <= 19'd0;
		WeightsStore6[623] <= 19'd0;
		WeightsStore6[624] <= 19'd0;
		WeightsStore6[625] <= 19'd0;
		WeightsStore6[626] <= 19'd0;
		WeightsStore6[627] <= 19'd0;
		WeightsStore6[628] <= 19'd0;
		WeightsStore6[629] <= 19'd0;
		WeightsStore6[630] <= 19'd0;
		WeightsStore6[631] <= 19'd0;
		WeightsStore6[632] <= 19'd0;
		WeightsStore6[633] <= 19'd0;
		WeightsStore6[634] <= 19'd0;
		WeightsStore6[635] <= 19'd0;
		WeightsStore6[636] <= 19'd0;
		WeightsStore6[637] <= 19'd0;
		WeightsStore6[638] <= 19'd0;
		WeightsStore6[639] <= 19'd0;
		WeightsStore6[640] <= 19'd0;
		WeightsStore6[641] <= 19'd0;
		WeightsStore6[642] <= 19'd0;
		WeightsStore6[643] <= 19'd0;
		WeightsStore6[644] <= 19'd0;
		WeightsStore6[645] <= 19'd0;
		WeightsStore6[646] <= 19'd0;
		WeightsStore6[647] <= 19'd0;
		WeightsStore6[648] <= 19'd0;
		WeightsStore6[649] <= 19'd0;
		WeightsStore6[650] <= 19'd0;
		WeightsStore6[651] <= 19'd0;
		WeightsStore6[652] <= 19'd0;
		WeightsStore6[653] <= 19'd0;
		WeightsStore6[654] <= 19'd0;
		WeightsStore6[655] <= 19'd0;
		WeightsStore6[656] <= 19'd0;
		WeightsStore6[657] <= 19'd0;
		WeightsStore6[658] <= 19'd0;
		WeightsStore6[659] <= 19'd0;
		WeightsStore6[660] <= 19'd0;
		WeightsStore6[661] <= 19'd0;
		WeightsStore6[662] <= 19'd0;
		WeightsStore6[663] <= 19'd0;
		WeightsStore6[664] <= 19'd0;
		WeightsStore6[665] <= 19'd0;
		WeightsStore6[666] <= 19'd0;
		WeightsStore6[667] <= 19'd0;
		WeightsStore6[668] <= 19'd0;
		WeightsStore6[669] <= 19'd0;
		WeightsStore6[670] <= 19'd0;
		WeightsStore6[671] <= 19'd0;
		WeightsStore6[672] <= 19'd0;
		WeightsStore6[673] <= 19'd0;
		WeightsStore6[674] <= 19'd0;
		WeightsStore6[675] <= 19'd0;
		WeightsStore6[676] <= 19'd0;
		WeightsStore6[677] <= 19'd0;
		WeightsStore6[678] <= 19'd0;
		WeightsStore6[679] <= 19'd0;
		WeightsStore6[680] <= 19'd0;
		WeightsStore6[681] <= 19'd0;
		WeightsStore6[682] <= 19'd0;
		WeightsStore6[683] <= 19'd0;
		WeightsStore6[684] <= 19'd0;
		WeightsStore6[685] <= 19'd0;
		WeightsStore6[686] <= 19'd0;
		WeightsStore6[687] <= 19'd0;
		WeightsStore6[688] <= 19'd0;
		WeightsStore6[689] <= 19'd0;
		WeightsStore6[690] <= 19'd0;
		WeightsStore6[691] <= 19'd0;
		WeightsStore6[692] <= 19'd0;
		WeightsStore6[693] <= 19'd0;
		WeightsStore6[694] <= 19'd0;
		WeightsStore6[695] <= 19'd0;
		WeightsStore6[696] <= 19'd0;
		WeightsStore6[697] <= 19'd0;
		WeightsStore6[698] <= 19'd0;
		WeightsStore6[699] <= 19'd0;
		WeightsStore6[700] <= 19'd0;
		WeightsStore6[701] <= 19'd0;
		WeightsStore6[702] <= 19'd0;
		WeightsStore6[703] <= 19'd0;
		WeightsStore6[704] <= 19'd0;
		WeightsStore6[705] <= 19'd0;
		WeightsStore6[706] <= 19'd0;
		WeightsStore6[707] <= 19'd0;
		WeightsStore6[708] <= 19'd0;
		WeightsStore6[709] <= 19'd0;
		WeightsStore6[710] <= 19'd0;
		WeightsStore6[711] <= 19'd0;
		WeightsStore6[712] <= 19'd0;
		WeightsStore6[713] <= 19'd0;
		WeightsStore6[714] <= 19'd0;
		WeightsStore6[715] <= 19'd0;
		WeightsStore6[716] <= 19'd0;
		WeightsStore6[717] <= 19'd0;
		WeightsStore6[718] <= 19'd0;
		WeightsStore6[719] <= 19'd0;
		WeightsStore6[720] <= 19'd0;
		WeightsStore6[721] <= 19'd0;
		WeightsStore6[722] <= 19'd0;
		WeightsStore6[723] <= 19'd0;
		WeightsStore6[724] <= 19'd0;
		WeightsStore6[725] <= 19'd0;
		WeightsStore6[726] <= 19'd0;
		WeightsStore6[727] <= 19'd0;
		WeightsStore6[728] <= 19'd0;
		WeightsStore6[729] <= 19'd0;
		WeightsStore6[730] <= 19'd0;
		WeightsStore6[731] <= 19'd0;
		WeightsStore6[732] <= 19'd0;
		WeightsStore6[733] <= 19'd0;
		WeightsStore6[734] <= 19'd0;
		WeightsStore6[735] <= 19'd0;
		WeightsStore6[736] <= 19'd0;
		WeightsStore6[737] <= 19'd0;
		WeightsStore6[738] <= 19'd0;
		WeightsStore6[739] <= 19'd0;
		WeightsStore6[740] <= 19'd0;
		WeightsStore6[741] <= 19'd0;
		WeightsStore6[742] <= 19'd0;
		WeightsStore6[743] <= 19'd0;
		WeightsStore6[744] <= 19'd0;
		WeightsStore6[745] <= 19'd0;
		WeightsStore6[746] <= 19'd0;
		WeightsStore6[747] <= 19'd0;
		WeightsStore6[748] <= 19'd0;
		WeightsStore6[749] <= 19'd0;
		WeightsStore6[750] <= 19'd0;
		WeightsStore6[751] <= 19'd0;
		WeightsStore6[752] <= 19'd0;
		WeightsStore6[753] <= 19'd0;
		WeightsStore6[754] <= 19'd0;
		WeightsStore6[755] <= 19'd0;
		WeightsStore6[756] <= 19'd0;
		WeightsStore6[757] <= 19'd0;
		WeightsStore6[758] <= 19'd0;
		WeightsStore6[759] <= 19'd0;
		WeightsStore6[760] <= 19'd0;
		WeightsStore6[761] <= 19'd0;
		WeightsStore6[762] <= 19'd0;
		WeightsStore6[763] <= 19'd0;
		WeightsStore6[764] <= 19'd0;
		WeightsStore6[765] <= 19'd0;
		WeightsStore6[766] <= 19'd0;
		WeightsStore6[767] <= 19'd0;
		WeightsStore6[768] <= 19'd0;
		WeightsStore6[769] <= 19'd0;
		WeightsStore6[770] <= 19'd0;
		WeightsStore6[771] <= 19'd0;
		WeightsStore6[772] <= 19'd0;
		WeightsStore6[773] <= 19'd0;
		WeightsStore6[774] <= 19'd0;
		WeightsStore6[775] <= 19'd0;
		WeightsStore6[776] <= 19'd0;
		WeightsStore6[777] <= 19'd0;
		WeightsStore6[778] <= 19'd0;
		WeightsStore6[779] <= 19'd0;
		WeightsStore6[780] <= 19'd0;
		WeightsStore6[781] <= 19'd0;
		WeightsStore6[782] <= 19'd0;
		WeightsStore6[783] <= 19'd0;
		WeightsStore6[784] <= 19'd0;
		WeightsStore7[0] <= 19'd0;
		WeightsStore7[1] <= 19'd0;
		WeightsStore7[2] <= 19'd0;
		WeightsStore7[3] <= 19'd0;
		WeightsStore7[4] <= 19'd0;
		WeightsStore7[5] <= 19'd0;
		WeightsStore7[6] <= 19'd0;
		WeightsStore7[7] <= 19'd0;
		WeightsStore7[8] <= 19'd0;
		WeightsStore7[9] <= 19'd0;
		WeightsStore7[10] <= 19'd0;
		WeightsStore7[11] <= 19'd0;
		WeightsStore7[12] <= 19'd0;
		WeightsStore7[13] <= 19'd0;
		WeightsStore7[14] <= 19'd0;
		WeightsStore7[15] <= 19'd0;
		WeightsStore7[16] <= 19'd0;
		WeightsStore7[17] <= 19'd0;
		WeightsStore7[18] <= 19'd0;
		WeightsStore7[19] <= 19'd0;
		WeightsStore7[20] <= 19'd0;
		WeightsStore7[21] <= 19'd0;
		WeightsStore7[22] <= 19'd0;
		WeightsStore7[23] <= 19'd0;
		WeightsStore7[24] <= 19'd0;
		WeightsStore7[25] <= 19'd0;
		WeightsStore7[26] <= 19'd0;
		WeightsStore7[27] <= 19'd0;
		WeightsStore7[28] <= 19'd0;
		WeightsStore7[29] <= 19'd0;
		WeightsStore7[30] <= 19'd0;
		WeightsStore7[31] <= 19'd0;
		WeightsStore7[32] <= 19'd0;
		WeightsStore7[33] <= 19'd0;
		WeightsStore7[34] <= 19'd0;
		WeightsStore7[35] <= 19'd0;
		WeightsStore7[36] <= 19'd0;
		WeightsStore7[37] <= 19'd0;
		WeightsStore7[38] <= 19'd0;
		WeightsStore7[39] <= 19'd0;
		WeightsStore7[40] <= 19'd0;
		WeightsStore7[41] <= 19'd0;
		WeightsStore7[42] <= 19'd0;
		WeightsStore7[43] <= 19'd0;
		WeightsStore7[44] <= 19'd0;
		WeightsStore7[45] <= 19'd0;
		WeightsStore7[46] <= 19'd0;
		WeightsStore7[47] <= 19'd0;
		WeightsStore7[48] <= 19'd0;
		WeightsStore7[49] <= 19'd0;
		WeightsStore7[50] <= 19'd0;
		WeightsStore7[51] <= 19'd0;
		WeightsStore7[52] <= 19'd0;
		WeightsStore7[53] <= 19'd0;
		WeightsStore7[54] <= 19'd0;
		WeightsStore7[55] <= 19'd0;
		WeightsStore7[56] <= 19'd0;
		WeightsStore7[57] <= 19'd0;
		WeightsStore7[58] <= 19'd0;
		WeightsStore7[59] <= 19'd0;
		WeightsStore7[60] <= 19'd0;
		WeightsStore7[61] <= 19'd0;
		WeightsStore7[62] <= 19'd0;
		WeightsStore7[63] <= 19'd0;
		WeightsStore7[64] <= 19'd0;
		WeightsStore7[65] <= 19'd0;
		WeightsStore7[66] <= 19'd0;
		WeightsStore7[67] <= 19'd0;
		WeightsStore7[68] <= 19'd0;
		WeightsStore7[69] <= 19'd0;
		WeightsStore7[70] <= 19'd0;
		WeightsStore7[71] <= 19'd0;
		WeightsStore7[72] <= 19'd0;
		WeightsStore7[73] <= 19'd0;
		WeightsStore7[74] <= 19'd0;
		WeightsStore7[75] <= 19'd0;
		WeightsStore7[76] <= 19'd0;
		WeightsStore7[77] <= 19'd0;
		WeightsStore7[78] <= 19'd0;
		WeightsStore7[79] <= 19'd0;
		WeightsStore7[80] <= 19'd0;
		WeightsStore7[81] <= 19'd0;
		WeightsStore7[82] <= 19'd0;
		WeightsStore7[83] <= 19'd0;
		WeightsStore7[84] <= 19'd0;
		WeightsStore7[85] <= 19'd0;
		WeightsStore7[86] <= 19'd0;
		WeightsStore7[87] <= 19'd0;
		WeightsStore7[88] <= 19'd0;
		WeightsStore7[89] <= 19'd0;
		WeightsStore7[90] <= 19'd0;
		WeightsStore7[91] <= 19'd0;
		WeightsStore7[92] <= 19'd0;
		WeightsStore7[93] <= 19'd0;
		WeightsStore7[94] <= 19'd0;
		WeightsStore7[95] <= 19'd0;
		WeightsStore7[96] <= 19'd0;
		WeightsStore7[97] <= 19'd0;
		WeightsStore7[98] <= 19'd0;
		WeightsStore7[99] <= 19'd0;
		WeightsStore7[100] <= 19'd0;
		WeightsStore7[101] <= 19'd0;
		WeightsStore7[102] <= 19'd0;
		WeightsStore7[103] <= 19'd0;
		WeightsStore7[104] <= 19'd0;
		WeightsStore7[105] <= 19'd0;
		WeightsStore7[106] <= 19'd0;
		WeightsStore7[107] <= 19'd0;
		WeightsStore7[108] <= 19'd0;
		WeightsStore7[109] <= 19'd0;
		WeightsStore7[110] <= 19'd0;
		WeightsStore7[111] <= 19'd0;
		WeightsStore7[112] <= 19'd0;
		WeightsStore7[113] <= 19'd0;
		WeightsStore7[114] <= 19'd0;
		WeightsStore7[115] <= 19'd0;
		WeightsStore7[116] <= 19'd0;
		WeightsStore7[117] <= 19'd0;
		WeightsStore7[118] <= 19'd0;
		WeightsStore7[119] <= 19'd0;
		WeightsStore7[120] <= 19'd0;
		WeightsStore7[121] <= 19'd0;
		WeightsStore7[122] <= 19'd0;
		WeightsStore7[123] <= 19'd0;
		WeightsStore7[124] <= 19'd0;
		WeightsStore7[125] <= 19'd0;
		WeightsStore7[126] <= 19'd0;
		WeightsStore7[127] <= 19'd0;
		WeightsStore7[128] <= 19'd0;
		WeightsStore7[129] <= 19'd0;
		WeightsStore7[130] <= 19'd0;
		WeightsStore7[131] <= 19'd0;
		WeightsStore7[132] <= 19'd0;
		WeightsStore7[133] <= 19'd0;
		WeightsStore7[134] <= 19'd0;
		WeightsStore7[135] <= 19'd0;
		WeightsStore7[136] <= 19'd0;
		WeightsStore7[137] <= 19'd0;
		WeightsStore7[138] <= 19'd0;
		WeightsStore7[139] <= 19'd0;
		WeightsStore7[140] <= 19'd0;
		WeightsStore7[141] <= 19'd0;
		WeightsStore7[142] <= 19'd0;
		WeightsStore7[143] <= 19'd0;
		WeightsStore7[144] <= 19'd0;
		WeightsStore7[145] <= 19'd0;
		WeightsStore7[146] <= 19'd0;
		WeightsStore7[147] <= 19'd0;
		WeightsStore7[148] <= 19'd0;
		WeightsStore7[149] <= 19'd0;
		WeightsStore7[150] <= 19'd0;
		WeightsStore7[151] <= 19'd0;
		WeightsStore7[152] <= 19'd0;
		WeightsStore7[153] <= 19'd0;
		WeightsStore7[154] <= 19'd0;
		WeightsStore7[155] <= 19'd0;
		WeightsStore7[156] <= 19'd0;
		WeightsStore7[157] <= 19'd0;
		WeightsStore7[158] <= 19'd0;
		WeightsStore7[159] <= 19'd0;
		WeightsStore7[160] <= 19'd0;
		WeightsStore7[161] <= 19'd0;
		WeightsStore7[162] <= 19'd0;
		WeightsStore7[163] <= 19'd0;
		WeightsStore7[164] <= 19'd0;
		WeightsStore7[165] <= 19'd0;
		WeightsStore7[166] <= 19'd0;
		WeightsStore7[167] <= 19'd0;
		WeightsStore7[168] <= 19'd0;
		WeightsStore7[169] <= 19'd0;
		WeightsStore7[170] <= 19'd0;
		WeightsStore7[171] <= 19'd0;
		WeightsStore7[172] <= 19'd0;
		WeightsStore7[173] <= 19'd0;
		WeightsStore7[174] <= 19'd0;
		WeightsStore7[175] <= 19'd0;
		WeightsStore7[176] <= 19'd0;
		WeightsStore7[177] <= 19'd0;
		WeightsStore7[178] <= 19'd0;
		WeightsStore7[179] <= 19'd0;
		WeightsStore7[180] <= 19'd0;
		WeightsStore7[181] <= 19'd0;
		WeightsStore7[182] <= 19'd0;
		WeightsStore7[183] <= 19'd0;
		WeightsStore7[184] <= 19'd0;
		WeightsStore7[185] <= 19'd0;
		WeightsStore7[186] <= 19'd0;
		WeightsStore7[187] <= 19'd0;
		WeightsStore7[188] <= 19'd0;
		WeightsStore7[189] <= 19'd0;
		WeightsStore7[190] <= 19'd0;
		WeightsStore7[191] <= 19'd0;
		WeightsStore7[192] <= 19'd0;
		WeightsStore7[193] <= 19'd0;
		WeightsStore7[194] <= 19'd0;
		WeightsStore7[195] <= 19'd0;
		WeightsStore7[196] <= 19'd0;
		WeightsStore7[197] <= 19'd0;
		WeightsStore7[198] <= 19'd0;
		WeightsStore7[199] <= 19'd0;
		WeightsStore7[200] <= 19'd0;
		WeightsStore7[201] <= 19'd0;
		WeightsStore7[202] <= 19'd0;
		WeightsStore7[203] <= 19'd0;
		WeightsStore7[204] <= 19'd0;
		WeightsStore7[205] <= 19'd0;
		WeightsStore7[206] <= 19'd0;
		WeightsStore7[207] <= 19'd0;
		WeightsStore7[208] <= 19'd0;
		WeightsStore7[209] <= 19'd0;
		WeightsStore7[210] <= 19'd0;
		WeightsStore7[211] <= 19'd0;
		WeightsStore7[212] <= 19'd0;
		WeightsStore7[213] <= 19'd0;
		WeightsStore7[214] <= 19'd0;
		WeightsStore7[215] <= 19'd0;
		WeightsStore7[216] <= 19'd0;
		WeightsStore7[217] <= 19'd0;
		WeightsStore7[218] <= 19'd0;
		WeightsStore7[219] <= 19'd0;
		WeightsStore7[220] <= 19'd0;
		WeightsStore7[221] <= 19'd0;
		WeightsStore7[222] <= 19'd0;
		WeightsStore7[223] <= 19'd0;
		WeightsStore7[224] <= 19'd0;
		WeightsStore7[225] <= 19'd0;
		WeightsStore7[226] <= 19'd0;
		WeightsStore7[227] <= 19'd0;
		WeightsStore7[228] <= 19'd0;
		WeightsStore7[229] <= 19'd0;
		WeightsStore7[230] <= 19'd0;
		WeightsStore7[231] <= 19'd0;
		WeightsStore7[232] <= 19'd0;
		WeightsStore7[233] <= 19'd0;
		WeightsStore7[234] <= 19'd0;
		WeightsStore7[235] <= 19'd0;
		WeightsStore7[236] <= 19'd0;
		WeightsStore7[237] <= 19'd0;
		WeightsStore7[238] <= 19'd0;
		WeightsStore7[239] <= 19'd0;
		WeightsStore7[240] <= 19'd0;
		WeightsStore7[241] <= 19'd0;
		WeightsStore7[242] <= 19'd0;
		WeightsStore7[243] <= 19'd0;
		WeightsStore7[244] <= 19'd0;
		WeightsStore7[245] <= 19'd0;
		WeightsStore7[246] <= 19'd0;
		WeightsStore7[247] <= 19'd0;
		WeightsStore7[248] <= 19'd0;
		WeightsStore7[249] <= 19'd0;
		WeightsStore7[250] <= 19'd0;
		WeightsStore7[251] <= 19'd0;
		WeightsStore7[252] <= 19'd0;
		WeightsStore7[253] <= 19'd0;
		WeightsStore7[254] <= 19'd0;
		WeightsStore7[255] <= 19'd0;
		WeightsStore7[256] <= 19'd0;
		WeightsStore7[257] <= 19'd0;
		WeightsStore7[258] <= 19'd0;
		WeightsStore7[259] <= 19'd0;
		WeightsStore7[260] <= 19'd0;
		WeightsStore7[261] <= 19'd0;
		WeightsStore7[262] <= 19'd0;
		WeightsStore7[263] <= 19'd0;
		WeightsStore7[264] <= 19'd0;
		WeightsStore7[265] <= 19'd0;
		WeightsStore7[266] <= 19'd0;
		WeightsStore7[267] <= 19'd0;
		WeightsStore7[268] <= 19'd0;
		WeightsStore7[269] <= 19'd0;
		WeightsStore7[270] <= 19'd0;
		WeightsStore7[271] <= 19'd0;
		WeightsStore7[272] <= 19'd0;
		WeightsStore7[273] <= 19'd0;
		WeightsStore7[274] <= 19'd0;
		WeightsStore7[275] <= 19'd0;
		WeightsStore7[276] <= 19'd0;
		WeightsStore7[277] <= 19'd0;
		WeightsStore7[278] <= 19'd0;
		WeightsStore7[279] <= 19'd0;
		WeightsStore7[280] <= 19'd0;
		WeightsStore7[281] <= 19'd0;
		WeightsStore7[282] <= 19'd0;
		WeightsStore7[283] <= 19'd0;
		WeightsStore7[284] <= 19'd0;
		WeightsStore7[285] <= 19'd0;
		WeightsStore7[286] <= 19'd0;
		WeightsStore7[287] <= 19'd0;
		WeightsStore7[288] <= 19'd0;
		WeightsStore7[289] <= 19'd0;
		WeightsStore7[290] <= 19'd0;
		WeightsStore7[291] <= 19'd0;
		WeightsStore7[292] <= 19'd0;
		WeightsStore7[293] <= 19'd0;
		WeightsStore7[294] <= 19'd0;
		WeightsStore7[295] <= 19'd0;
		WeightsStore7[296] <= 19'd0;
		WeightsStore7[297] <= 19'd0;
		WeightsStore7[298] <= 19'd0;
		WeightsStore7[299] <= 19'd0;
		WeightsStore7[300] <= 19'd0;
		WeightsStore7[301] <= 19'd0;
		WeightsStore7[302] <= 19'd0;
		WeightsStore7[303] <= 19'd0;
		WeightsStore7[304] <= 19'd0;
		WeightsStore7[305] <= 19'd0;
		WeightsStore7[306] <= 19'd0;
		WeightsStore7[307] <= 19'd0;
		WeightsStore7[308] <= 19'd0;
		WeightsStore7[309] <= 19'd0;
		WeightsStore7[310] <= 19'd0;
		WeightsStore7[311] <= 19'd0;
		WeightsStore7[312] <= 19'd0;
		WeightsStore7[313] <= 19'd0;
		WeightsStore7[314] <= 19'd0;
		WeightsStore7[315] <= 19'd0;
		WeightsStore7[316] <= 19'd0;
		WeightsStore7[317] <= 19'd0;
		WeightsStore7[318] <= 19'd0;
		WeightsStore7[319] <= 19'd0;
		WeightsStore7[320] <= 19'd0;
		WeightsStore7[321] <= 19'd0;
		WeightsStore7[322] <= 19'd0;
		WeightsStore7[323] <= 19'd0;
		WeightsStore7[324] <= 19'd0;
		WeightsStore7[325] <= 19'd0;
		WeightsStore7[326] <= 19'd0;
		WeightsStore7[327] <= 19'd0;
		WeightsStore7[328] <= 19'd0;
		WeightsStore7[329] <= 19'd0;
		WeightsStore7[330] <= 19'd0;
		WeightsStore7[331] <= 19'd0;
		WeightsStore7[332] <= 19'd0;
		WeightsStore7[333] <= 19'd0;
		WeightsStore7[334] <= 19'd0;
		WeightsStore7[335] <= 19'd0;
		WeightsStore7[336] <= 19'd0;
		WeightsStore7[337] <= 19'd0;
		WeightsStore7[338] <= 19'd0;
		WeightsStore7[339] <= 19'd0;
		WeightsStore7[340] <= 19'd0;
		WeightsStore7[341] <= 19'd0;
		WeightsStore7[342] <= 19'd0;
		WeightsStore7[343] <= 19'd0;
		WeightsStore7[344] <= 19'd0;
		WeightsStore7[345] <= 19'd0;
		WeightsStore7[346] <= 19'd0;
		WeightsStore7[347] <= 19'd0;
		WeightsStore7[348] <= 19'd0;
		WeightsStore7[349] <= 19'd0;
		WeightsStore7[350] <= 19'd0;
		WeightsStore7[351] <= 19'd0;
		WeightsStore7[352] <= 19'd0;
		WeightsStore7[353] <= 19'd0;
		WeightsStore7[354] <= 19'd0;
		WeightsStore7[355] <= 19'd0;
		WeightsStore7[356] <= 19'd0;
		WeightsStore7[357] <= 19'd0;
		WeightsStore7[358] <= 19'd0;
		WeightsStore7[359] <= 19'd0;
		WeightsStore7[360] <= 19'd0;
		WeightsStore7[361] <= 19'd0;
		WeightsStore7[362] <= 19'd0;
		WeightsStore7[363] <= 19'd0;
		WeightsStore7[364] <= 19'd0;
		WeightsStore7[365] <= 19'd0;
		WeightsStore7[366] <= 19'd0;
		WeightsStore7[367] <= 19'd0;
		WeightsStore7[368] <= 19'd0;
		WeightsStore7[369] <= 19'd0;
		WeightsStore7[370] <= 19'd0;
		WeightsStore7[371] <= 19'd0;
		WeightsStore7[372] <= 19'd0;
		WeightsStore7[373] <= 19'd0;
		WeightsStore7[374] <= 19'd0;
		WeightsStore7[375] <= 19'd0;
		WeightsStore7[376] <= 19'd0;
		WeightsStore7[377] <= 19'd0;
		WeightsStore7[378] <= 19'd0;
		WeightsStore7[379] <= 19'd0;
		WeightsStore7[380] <= 19'd0;
		WeightsStore7[381] <= 19'd0;
		WeightsStore7[382] <= 19'd0;
		WeightsStore7[383] <= 19'd0;
		WeightsStore7[384] <= 19'd0;
		WeightsStore7[385] <= 19'd0;
		WeightsStore7[386] <= 19'd0;
		WeightsStore7[387] <= 19'd0;
		WeightsStore7[388] <= 19'd0;
		WeightsStore7[389] <= 19'd0;
		WeightsStore7[390] <= 19'd0;
		WeightsStore7[391] <= 19'd0;
		WeightsStore7[392] <= 19'd0;
		WeightsStore7[393] <= 19'd0;
		WeightsStore7[394] <= 19'd0;
		WeightsStore7[395] <= 19'd0;
		WeightsStore7[396] <= 19'd0;
		WeightsStore7[397] <= 19'd0;
		WeightsStore7[398] <= 19'd0;
		WeightsStore7[399] <= 19'd0;
		WeightsStore7[400] <= 19'd0;
		WeightsStore7[401] <= 19'd0;
		WeightsStore7[402] <= 19'd0;
		WeightsStore7[403] <= 19'd0;
		WeightsStore7[404] <= 19'd0;
		WeightsStore7[405] <= 19'd0;
		WeightsStore7[406] <= 19'd0;
		WeightsStore7[407] <= 19'd0;
		WeightsStore7[408] <= 19'd0;
		WeightsStore7[409] <= 19'd0;
		WeightsStore7[410] <= 19'd0;
		WeightsStore7[411] <= 19'd0;
		WeightsStore7[412] <= 19'd0;
		WeightsStore7[413] <= 19'd0;
		WeightsStore7[414] <= 19'd0;
		WeightsStore7[415] <= 19'd0;
		WeightsStore7[416] <= 19'd0;
		WeightsStore7[417] <= 19'd0;
		WeightsStore7[418] <= 19'd0;
		WeightsStore7[419] <= 19'd0;
		WeightsStore7[420] <= 19'd0;
		WeightsStore7[421] <= 19'd0;
		WeightsStore7[422] <= 19'd0;
		WeightsStore7[423] <= 19'd0;
		WeightsStore7[424] <= 19'd0;
		WeightsStore7[425] <= 19'd0;
		WeightsStore7[426] <= 19'd0;
		WeightsStore7[427] <= 19'd0;
		WeightsStore7[428] <= 19'd0;
		WeightsStore7[429] <= 19'd0;
		WeightsStore7[430] <= 19'd0;
		WeightsStore7[431] <= 19'd0;
		WeightsStore7[432] <= 19'd0;
		WeightsStore7[433] <= 19'd0;
		WeightsStore7[434] <= 19'd0;
		WeightsStore7[435] <= 19'd0;
		WeightsStore7[436] <= 19'd0;
		WeightsStore7[437] <= 19'd0;
		WeightsStore7[438] <= 19'd0;
		WeightsStore7[439] <= 19'd0;
		WeightsStore7[440] <= 19'd0;
		WeightsStore7[441] <= 19'd0;
		WeightsStore7[442] <= 19'd0;
		WeightsStore7[443] <= 19'd0;
		WeightsStore7[444] <= 19'd0;
		WeightsStore7[445] <= 19'd0;
		WeightsStore7[446] <= 19'd0;
		WeightsStore7[447] <= 19'd0;
		WeightsStore7[448] <= 19'd0;
		WeightsStore7[449] <= 19'd0;
		WeightsStore7[450] <= 19'd0;
		WeightsStore7[451] <= 19'd0;
		WeightsStore7[452] <= 19'd0;
		WeightsStore7[453] <= 19'd0;
		WeightsStore7[454] <= 19'd0;
		WeightsStore7[455] <= 19'd0;
		WeightsStore7[456] <= 19'd0;
		WeightsStore7[457] <= 19'd0;
		WeightsStore7[458] <= 19'd0;
		WeightsStore7[459] <= 19'd0;
		WeightsStore7[460] <= 19'd0;
		WeightsStore7[461] <= 19'd0;
		WeightsStore7[462] <= 19'd0;
		WeightsStore7[463] <= 19'd0;
		WeightsStore7[464] <= 19'd0;
		WeightsStore7[465] <= 19'd0;
		WeightsStore7[466] <= 19'd0;
		WeightsStore7[467] <= 19'd0;
		WeightsStore7[468] <= 19'd0;
		WeightsStore7[469] <= 19'd0;
		WeightsStore7[470] <= 19'd0;
		WeightsStore7[471] <= 19'd0;
		WeightsStore7[472] <= 19'd0;
		WeightsStore7[473] <= 19'd0;
		WeightsStore7[474] <= 19'd0;
		WeightsStore7[475] <= 19'd0;
		WeightsStore7[476] <= 19'd0;
		WeightsStore7[477] <= 19'd0;
		WeightsStore7[478] <= 19'd0;
		WeightsStore7[479] <= 19'd0;
		WeightsStore7[480] <= 19'd0;
		WeightsStore7[481] <= 19'd0;
		WeightsStore7[482] <= 19'd0;
		WeightsStore7[483] <= 19'd0;
		WeightsStore7[484] <= 19'd0;
		WeightsStore7[485] <= 19'd0;
		WeightsStore7[486] <= 19'd0;
		WeightsStore7[487] <= 19'd0;
		WeightsStore7[488] <= 19'd0;
		WeightsStore7[489] <= 19'd0;
		WeightsStore7[490] <= 19'd0;
		WeightsStore7[491] <= 19'd0;
		WeightsStore7[492] <= 19'd0;
		WeightsStore7[493] <= 19'd0;
		WeightsStore7[494] <= 19'd0;
		WeightsStore7[495] <= 19'd0;
		WeightsStore7[496] <= 19'd0;
		WeightsStore7[497] <= 19'd0;
		WeightsStore7[498] <= 19'd0;
		WeightsStore7[499] <= 19'd0;
		WeightsStore7[500] <= 19'd0;
		WeightsStore7[501] <= 19'd0;
		WeightsStore7[502] <= 19'd0;
		WeightsStore7[503] <= 19'd0;
		WeightsStore7[504] <= 19'd0;
		WeightsStore7[505] <= 19'd0;
		WeightsStore7[506] <= 19'd0;
		WeightsStore7[507] <= 19'd0;
		WeightsStore7[508] <= 19'd0;
		WeightsStore7[509] <= 19'd0;
		WeightsStore7[510] <= 19'd0;
		WeightsStore7[511] <= 19'd0;
		WeightsStore7[512] <= 19'd0;
		WeightsStore7[513] <= 19'd0;
		WeightsStore7[514] <= 19'd0;
		WeightsStore7[515] <= 19'd0;
		WeightsStore7[516] <= 19'd0;
		WeightsStore7[517] <= 19'd0;
		WeightsStore7[518] <= 19'd0;
		WeightsStore7[519] <= 19'd0;
		WeightsStore7[520] <= 19'd0;
		WeightsStore7[521] <= 19'd0;
		WeightsStore7[522] <= 19'd0;
		WeightsStore7[523] <= 19'd0;
		WeightsStore7[524] <= 19'd0;
		WeightsStore7[525] <= 19'd0;
		WeightsStore7[526] <= 19'd0;
		WeightsStore7[527] <= 19'd0;
		WeightsStore7[528] <= 19'd0;
		WeightsStore7[529] <= 19'd0;
		WeightsStore7[530] <= 19'd0;
		WeightsStore7[531] <= 19'd0;
		WeightsStore7[532] <= 19'd0;
		WeightsStore7[533] <= 19'd0;
		WeightsStore7[534] <= 19'd0;
		WeightsStore7[535] <= 19'd0;
		WeightsStore7[536] <= 19'd0;
		WeightsStore7[537] <= 19'd0;
		WeightsStore7[538] <= 19'd0;
		WeightsStore7[539] <= 19'd0;
		WeightsStore7[540] <= 19'd0;
		WeightsStore7[541] <= 19'd0;
		WeightsStore7[542] <= 19'd0;
		WeightsStore7[543] <= 19'd0;
		WeightsStore7[544] <= 19'd0;
		WeightsStore7[545] <= 19'd0;
		WeightsStore7[546] <= 19'd0;
		WeightsStore7[547] <= 19'd0;
		WeightsStore7[548] <= 19'd0;
		WeightsStore7[549] <= 19'd0;
		WeightsStore7[550] <= 19'd0;
		WeightsStore7[551] <= 19'd0;
		WeightsStore7[552] <= 19'd0;
		WeightsStore7[553] <= 19'd0;
		WeightsStore7[554] <= 19'd0;
		WeightsStore7[555] <= 19'd0;
		WeightsStore7[556] <= 19'd0;
		WeightsStore7[557] <= 19'd0;
		WeightsStore7[558] <= 19'd0;
		WeightsStore7[559] <= 19'd0;
		WeightsStore7[560] <= 19'd0;
		WeightsStore7[561] <= 19'd0;
		WeightsStore7[562] <= 19'd0;
		WeightsStore7[563] <= 19'd0;
		WeightsStore7[564] <= 19'd0;
		WeightsStore7[565] <= 19'd0;
		WeightsStore7[566] <= 19'd0;
		WeightsStore7[567] <= 19'd0;
		WeightsStore7[568] <= 19'd0;
		WeightsStore7[569] <= 19'd0;
		WeightsStore7[570] <= 19'd0;
		WeightsStore7[571] <= 19'd0;
		WeightsStore7[572] <= 19'd0;
		WeightsStore7[573] <= 19'd0;
		WeightsStore7[574] <= 19'd0;
		WeightsStore7[575] <= 19'd0;
		WeightsStore7[576] <= 19'd0;
		WeightsStore7[577] <= 19'd0;
		WeightsStore7[578] <= 19'd0;
		WeightsStore7[579] <= 19'd0;
		WeightsStore7[580] <= 19'd0;
		WeightsStore7[581] <= 19'd0;
		WeightsStore7[582] <= 19'd0;
		WeightsStore7[583] <= 19'd0;
		WeightsStore7[584] <= 19'd0;
		WeightsStore7[585] <= 19'd0;
		WeightsStore7[586] <= 19'd0;
		WeightsStore7[587] <= 19'd0;
		WeightsStore7[588] <= 19'd0;
		WeightsStore7[589] <= 19'd0;
		WeightsStore7[590] <= 19'd0;
		WeightsStore7[591] <= 19'd0;
		WeightsStore7[592] <= 19'd0;
		WeightsStore7[593] <= 19'd0;
		WeightsStore7[594] <= 19'd0;
		WeightsStore7[595] <= 19'd0;
		WeightsStore7[596] <= 19'd0;
		WeightsStore7[597] <= 19'd0;
		WeightsStore7[598] <= 19'd0;
		WeightsStore7[599] <= 19'd0;
		WeightsStore7[600] <= 19'd0;
		WeightsStore7[601] <= 19'd0;
		WeightsStore7[602] <= 19'd0;
		WeightsStore7[603] <= 19'd0;
		WeightsStore7[604] <= 19'd0;
		WeightsStore7[605] <= 19'd0;
		WeightsStore7[606] <= 19'd0;
		WeightsStore7[607] <= 19'd0;
		WeightsStore7[608] <= 19'd0;
		WeightsStore7[609] <= 19'd0;
		WeightsStore7[610] <= 19'd0;
		WeightsStore7[611] <= 19'd0;
		WeightsStore7[612] <= 19'd0;
		WeightsStore7[613] <= 19'd0;
		WeightsStore7[614] <= 19'd0;
		WeightsStore7[615] <= 19'd0;
		WeightsStore7[616] <= 19'd0;
		WeightsStore7[617] <= 19'd0;
		WeightsStore7[618] <= 19'd0;
		WeightsStore7[619] <= 19'd0;
		WeightsStore7[620] <= 19'd0;
		WeightsStore7[621] <= 19'd0;
		WeightsStore7[622] <= 19'd0;
		WeightsStore7[623] <= 19'd0;
		WeightsStore7[624] <= 19'd0;
		WeightsStore7[625] <= 19'd0;
		WeightsStore7[626] <= 19'd0;
		WeightsStore7[627] <= 19'd0;
		WeightsStore7[628] <= 19'd0;
		WeightsStore7[629] <= 19'd0;
		WeightsStore7[630] <= 19'd0;
		WeightsStore7[631] <= 19'd0;
		WeightsStore7[632] <= 19'd0;
		WeightsStore7[633] <= 19'd0;
		WeightsStore7[634] <= 19'd0;
		WeightsStore7[635] <= 19'd0;
		WeightsStore7[636] <= 19'd0;
		WeightsStore7[637] <= 19'd0;
		WeightsStore7[638] <= 19'd0;
		WeightsStore7[639] <= 19'd0;
		WeightsStore7[640] <= 19'd0;
		WeightsStore7[641] <= 19'd0;
		WeightsStore7[642] <= 19'd0;
		WeightsStore7[643] <= 19'd0;
		WeightsStore7[644] <= 19'd0;
		WeightsStore7[645] <= 19'd0;
		WeightsStore7[646] <= 19'd0;
		WeightsStore7[647] <= 19'd0;
		WeightsStore7[648] <= 19'd0;
		WeightsStore7[649] <= 19'd0;
		WeightsStore7[650] <= 19'd0;
		WeightsStore7[651] <= 19'd0;
		WeightsStore7[652] <= 19'd0;
		WeightsStore7[653] <= 19'd0;
		WeightsStore7[654] <= 19'd0;
		WeightsStore7[655] <= 19'd0;
		WeightsStore7[656] <= 19'd0;
		WeightsStore7[657] <= 19'd0;
		WeightsStore7[658] <= 19'd0;
		WeightsStore7[659] <= 19'd0;
		WeightsStore7[660] <= 19'd0;
		WeightsStore7[661] <= 19'd0;
		WeightsStore7[662] <= 19'd0;
		WeightsStore7[663] <= 19'd0;
		WeightsStore7[664] <= 19'd0;
		WeightsStore7[665] <= 19'd0;
		WeightsStore7[666] <= 19'd0;
		WeightsStore7[667] <= 19'd0;
		WeightsStore7[668] <= 19'd0;
		WeightsStore7[669] <= 19'd0;
		WeightsStore7[670] <= 19'd0;
		WeightsStore7[671] <= 19'd0;
		WeightsStore7[672] <= 19'd0;
		WeightsStore7[673] <= 19'd0;
		WeightsStore7[674] <= 19'd0;
		WeightsStore7[675] <= 19'd0;
		WeightsStore7[676] <= 19'd0;
		WeightsStore7[677] <= 19'd0;
		WeightsStore7[678] <= 19'd0;
		WeightsStore7[679] <= 19'd0;
		WeightsStore7[680] <= 19'd0;
		WeightsStore7[681] <= 19'd0;
		WeightsStore7[682] <= 19'd0;
		WeightsStore7[683] <= 19'd0;
		WeightsStore7[684] <= 19'd0;
		WeightsStore7[685] <= 19'd0;
		WeightsStore7[686] <= 19'd0;
		WeightsStore7[687] <= 19'd0;
		WeightsStore7[688] <= 19'd0;
		WeightsStore7[689] <= 19'd0;
		WeightsStore7[690] <= 19'd0;
		WeightsStore7[691] <= 19'd0;
		WeightsStore7[692] <= 19'd0;
		WeightsStore7[693] <= 19'd0;
		WeightsStore7[694] <= 19'd0;
		WeightsStore7[695] <= 19'd0;
		WeightsStore7[696] <= 19'd0;
		WeightsStore7[697] <= 19'd0;
		WeightsStore7[698] <= 19'd0;
		WeightsStore7[699] <= 19'd0;
		WeightsStore7[700] <= 19'd0;
		WeightsStore7[701] <= 19'd0;
		WeightsStore7[702] <= 19'd0;
		WeightsStore7[703] <= 19'd0;
		WeightsStore7[704] <= 19'd0;
		WeightsStore7[705] <= 19'd0;
		WeightsStore7[706] <= 19'd0;
		WeightsStore7[707] <= 19'd0;
		WeightsStore7[708] <= 19'd0;
		WeightsStore7[709] <= 19'd0;
		WeightsStore7[710] <= 19'd0;
		WeightsStore7[711] <= 19'd0;
		WeightsStore7[712] <= 19'd0;
		WeightsStore7[713] <= 19'd0;
		WeightsStore7[714] <= 19'd0;
		WeightsStore7[715] <= 19'd0;
		WeightsStore7[716] <= 19'd0;
		WeightsStore7[717] <= 19'd0;
		WeightsStore7[718] <= 19'd0;
		WeightsStore7[719] <= 19'd0;
		WeightsStore7[720] <= 19'd0;
		WeightsStore7[721] <= 19'd0;
		WeightsStore7[722] <= 19'd0;
		WeightsStore7[723] <= 19'd0;
		WeightsStore7[724] <= 19'd0;
		WeightsStore7[725] <= 19'd0;
		WeightsStore7[726] <= 19'd0;
		WeightsStore7[727] <= 19'd0;
		WeightsStore7[728] <= 19'd0;
		WeightsStore7[729] <= 19'd0;
		WeightsStore7[730] <= 19'd0;
		WeightsStore7[731] <= 19'd0;
		WeightsStore7[732] <= 19'd0;
		WeightsStore7[733] <= 19'd0;
		WeightsStore7[734] <= 19'd0;
		WeightsStore7[735] <= 19'd0;
		WeightsStore7[736] <= 19'd0;
		WeightsStore7[737] <= 19'd0;
		WeightsStore7[738] <= 19'd0;
		WeightsStore7[739] <= 19'd0;
		WeightsStore7[740] <= 19'd0;
		WeightsStore7[741] <= 19'd0;
		WeightsStore7[742] <= 19'd0;
		WeightsStore7[743] <= 19'd0;
		WeightsStore7[744] <= 19'd0;
		WeightsStore7[745] <= 19'd0;
		WeightsStore7[746] <= 19'd0;
		WeightsStore7[747] <= 19'd0;
		WeightsStore7[748] <= 19'd0;
		WeightsStore7[749] <= 19'd0;
		WeightsStore7[750] <= 19'd0;
		WeightsStore7[751] <= 19'd0;
		WeightsStore7[752] <= 19'd0;
		WeightsStore7[753] <= 19'd0;
		WeightsStore7[754] <= 19'd0;
		WeightsStore7[755] <= 19'd0;
		WeightsStore7[756] <= 19'd0;
		WeightsStore7[757] <= 19'd0;
		WeightsStore7[758] <= 19'd0;
		WeightsStore7[759] <= 19'd0;
		WeightsStore7[760] <= 19'd0;
		WeightsStore7[761] <= 19'd0;
		WeightsStore7[762] <= 19'd0;
		WeightsStore7[763] <= 19'd0;
		WeightsStore7[764] <= 19'd0;
		WeightsStore7[765] <= 19'd0;
		WeightsStore7[766] <= 19'd0;
		WeightsStore7[767] <= 19'd0;
		WeightsStore7[768] <= 19'd0;
		WeightsStore7[769] <= 19'd0;
		WeightsStore7[770] <= 19'd0;
		WeightsStore7[771] <= 19'd0;
		WeightsStore7[772] <= 19'd0;
		WeightsStore7[773] <= 19'd0;
		WeightsStore7[774] <= 19'd0;
		WeightsStore7[775] <= 19'd0;
		WeightsStore7[776] <= 19'd0;
		WeightsStore7[777] <= 19'd0;
		WeightsStore7[778] <= 19'd0;
		WeightsStore7[779] <= 19'd0;
		WeightsStore7[780] <= 19'd0;
		WeightsStore7[781] <= 19'd0;
		WeightsStore7[782] <= 19'd0;
		WeightsStore7[783] <= 19'd0;
		WeightsStore7[784] <= 19'd0;
		WeightsStore8[0] <= 19'd0;
		WeightsStore8[1] <= 19'd0;
		WeightsStore8[2] <= 19'd0;
		WeightsStore8[3] <= 19'd0;
		WeightsStore8[4] <= 19'd0;
		WeightsStore8[5] <= 19'd0;
		WeightsStore8[6] <= 19'd0;
		WeightsStore8[7] <= 19'd0;
		WeightsStore8[8] <= 19'd0;
		WeightsStore8[9] <= 19'd0;
		WeightsStore8[10] <= 19'd0;
		WeightsStore8[11] <= 19'd0;
		WeightsStore8[12] <= 19'd0;
		WeightsStore8[13] <= 19'd0;
		WeightsStore8[14] <= 19'd0;
		WeightsStore8[15] <= 19'd0;
		WeightsStore8[16] <= 19'd0;
		WeightsStore8[17] <= 19'd0;
		WeightsStore8[18] <= 19'd0;
		WeightsStore8[19] <= 19'd0;
		WeightsStore8[20] <= 19'd0;
		WeightsStore8[21] <= 19'd0;
		WeightsStore8[22] <= 19'd0;
		WeightsStore8[23] <= 19'd0;
		WeightsStore8[24] <= 19'd0;
		WeightsStore8[25] <= 19'd0;
		WeightsStore8[26] <= 19'd0;
		WeightsStore8[27] <= 19'd0;
		WeightsStore8[28] <= 19'd0;
		WeightsStore8[29] <= 19'd0;
		WeightsStore8[30] <= 19'd0;
		WeightsStore8[31] <= 19'd0;
		WeightsStore8[32] <= 19'd0;
		WeightsStore8[33] <= 19'd0;
		WeightsStore8[34] <= 19'd0;
		WeightsStore8[35] <= 19'd0;
		WeightsStore8[36] <= 19'd0;
		WeightsStore8[37] <= 19'd0;
		WeightsStore8[38] <= 19'd0;
		WeightsStore8[39] <= 19'd0;
		WeightsStore8[40] <= 19'd0;
		WeightsStore8[41] <= 19'd0;
		WeightsStore8[42] <= 19'd0;
		WeightsStore8[43] <= 19'd0;
		WeightsStore8[44] <= 19'd0;
		WeightsStore8[45] <= 19'd0;
		WeightsStore8[46] <= 19'd0;
		WeightsStore8[47] <= 19'd0;
		WeightsStore8[48] <= 19'd0;
		WeightsStore8[49] <= 19'd0;
		WeightsStore8[50] <= 19'd0;
		WeightsStore8[51] <= 19'd0;
		WeightsStore8[52] <= 19'd0;
		WeightsStore8[53] <= 19'd0;
		WeightsStore8[54] <= 19'd0;
		WeightsStore8[55] <= 19'd0;
		WeightsStore8[56] <= 19'd0;
		WeightsStore8[57] <= 19'd0;
		WeightsStore8[58] <= 19'd0;
		WeightsStore8[59] <= 19'd0;
		WeightsStore8[60] <= 19'd0;
		WeightsStore8[61] <= 19'd0;
		WeightsStore8[62] <= 19'd0;
		WeightsStore8[63] <= 19'd0;
		WeightsStore8[64] <= 19'd0;
		WeightsStore8[65] <= 19'd0;
		WeightsStore8[66] <= 19'd0;
		WeightsStore8[67] <= 19'd0;
		WeightsStore8[68] <= 19'd0;
		WeightsStore8[69] <= 19'd0;
		WeightsStore8[70] <= 19'd0;
		WeightsStore8[71] <= 19'd0;
		WeightsStore8[72] <= 19'd0;
		WeightsStore8[73] <= 19'd0;
		WeightsStore8[74] <= 19'd0;
		WeightsStore8[75] <= 19'd0;
		WeightsStore8[76] <= 19'd0;
		WeightsStore8[77] <= 19'd0;
		WeightsStore8[78] <= 19'd0;
		WeightsStore8[79] <= 19'd0;
		WeightsStore8[80] <= 19'd0;
		WeightsStore8[81] <= 19'd0;
		WeightsStore8[82] <= 19'd0;
		WeightsStore8[83] <= 19'd0;
		WeightsStore8[84] <= 19'd0;
		WeightsStore8[85] <= 19'd0;
		WeightsStore8[86] <= 19'd0;
		WeightsStore8[87] <= 19'd0;
		WeightsStore8[88] <= 19'd0;
		WeightsStore8[89] <= 19'd0;
		WeightsStore8[90] <= 19'd0;
		WeightsStore8[91] <= 19'd0;
		WeightsStore8[92] <= 19'd0;
		WeightsStore8[93] <= 19'd0;
		WeightsStore8[94] <= 19'd0;
		WeightsStore8[95] <= 19'd0;
		WeightsStore8[96] <= 19'd0;
		WeightsStore8[97] <= 19'd0;
		WeightsStore8[98] <= 19'd0;
		WeightsStore8[99] <= 19'd0;
		WeightsStore8[100] <= 19'd0;
		WeightsStore8[101] <= 19'd0;
		WeightsStore8[102] <= 19'd0;
		WeightsStore8[103] <= 19'd0;
		WeightsStore8[104] <= 19'd0;
		WeightsStore8[105] <= 19'd0;
		WeightsStore8[106] <= 19'd0;
		WeightsStore8[107] <= 19'd0;
		WeightsStore8[108] <= 19'd0;
		WeightsStore8[109] <= 19'd0;
		WeightsStore8[110] <= 19'd0;
		WeightsStore8[111] <= 19'd0;
		WeightsStore8[112] <= 19'd0;
		WeightsStore8[113] <= 19'd0;
		WeightsStore8[114] <= 19'd0;
		WeightsStore8[115] <= 19'd0;
		WeightsStore8[116] <= 19'd0;
		WeightsStore8[117] <= 19'd0;
		WeightsStore8[118] <= 19'd0;
		WeightsStore8[119] <= 19'd0;
		WeightsStore8[120] <= 19'd0;
		WeightsStore8[121] <= 19'd0;
		WeightsStore8[122] <= 19'd0;
		WeightsStore8[123] <= 19'd0;
		WeightsStore8[124] <= 19'd0;
		WeightsStore8[125] <= 19'd0;
		WeightsStore8[126] <= 19'd0;
		WeightsStore8[127] <= 19'd0;
		WeightsStore8[128] <= 19'd0;
		WeightsStore8[129] <= 19'd0;
		WeightsStore8[130] <= 19'd0;
		WeightsStore8[131] <= 19'd0;
		WeightsStore8[132] <= 19'd0;
		WeightsStore8[133] <= 19'd0;
		WeightsStore8[134] <= 19'd0;
		WeightsStore8[135] <= 19'd0;
		WeightsStore8[136] <= 19'd0;
		WeightsStore8[137] <= 19'd0;
		WeightsStore8[138] <= 19'd0;
		WeightsStore8[139] <= 19'd0;
		WeightsStore8[140] <= 19'd0;
		WeightsStore8[141] <= 19'd0;
		WeightsStore8[142] <= 19'd0;
		WeightsStore8[143] <= 19'd0;
		WeightsStore8[144] <= 19'd0;
		WeightsStore8[145] <= 19'd0;
		WeightsStore8[146] <= 19'd0;
		WeightsStore8[147] <= 19'd0;
		WeightsStore8[148] <= 19'd0;
		WeightsStore8[149] <= 19'd0;
		WeightsStore8[150] <= 19'd0;
		WeightsStore8[151] <= 19'd0;
		WeightsStore8[152] <= 19'd0;
		WeightsStore8[153] <= 19'd0;
		WeightsStore8[154] <= 19'd0;
		WeightsStore8[155] <= 19'd0;
		WeightsStore8[156] <= 19'd0;
		WeightsStore8[157] <= 19'd0;
		WeightsStore8[158] <= 19'd0;
		WeightsStore8[159] <= 19'd0;
		WeightsStore8[160] <= 19'd0;
		WeightsStore8[161] <= 19'd0;
		WeightsStore8[162] <= 19'd0;
		WeightsStore8[163] <= 19'd0;
		WeightsStore8[164] <= 19'd0;
		WeightsStore8[165] <= 19'd0;
		WeightsStore8[166] <= 19'd0;
		WeightsStore8[167] <= 19'd0;
		WeightsStore8[168] <= 19'd0;
		WeightsStore8[169] <= 19'd0;
		WeightsStore8[170] <= 19'd0;
		WeightsStore8[171] <= 19'd0;
		WeightsStore8[172] <= 19'd0;
		WeightsStore8[173] <= 19'd0;
		WeightsStore8[174] <= 19'd0;
		WeightsStore8[175] <= 19'd0;
		WeightsStore8[176] <= 19'd0;
		WeightsStore8[177] <= 19'd0;
		WeightsStore8[178] <= 19'd0;
		WeightsStore8[179] <= 19'd0;
		WeightsStore8[180] <= 19'd0;
		WeightsStore8[181] <= 19'd0;
		WeightsStore8[182] <= 19'd0;
		WeightsStore8[183] <= 19'd0;
		WeightsStore8[184] <= 19'd0;
		WeightsStore8[185] <= 19'd0;
		WeightsStore8[186] <= 19'd0;
		WeightsStore8[187] <= 19'd0;
		WeightsStore8[188] <= 19'd0;
		WeightsStore8[189] <= 19'd0;
		WeightsStore8[190] <= 19'd0;
		WeightsStore8[191] <= 19'd0;
		WeightsStore8[192] <= 19'd0;
		WeightsStore8[193] <= 19'd0;
		WeightsStore8[194] <= 19'd0;
		WeightsStore8[195] <= 19'd0;
		WeightsStore8[196] <= 19'd0;
		WeightsStore8[197] <= 19'd0;
		WeightsStore8[198] <= 19'd0;
		WeightsStore8[199] <= 19'd0;
		WeightsStore8[200] <= 19'd0;
		WeightsStore8[201] <= 19'd0;
		WeightsStore8[202] <= 19'd0;
		WeightsStore8[203] <= 19'd0;
		WeightsStore8[204] <= 19'd0;
		WeightsStore8[205] <= 19'd0;
		WeightsStore8[206] <= 19'd0;
		WeightsStore8[207] <= 19'd0;
		WeightsStore8[208] <= 19'd0;
		WeightsStore8[209] <= 19'd0;
		WeightsStore8[210] <= 19'd0;
		WeightsStore8[211] <= 19'd0;
		WeightsStore8[212] <= 19'd0;
		WeightsStore8[213] <= 19'd0;
		WeightsStore8[214] <= 19'd0;
		WeightsStore8[215] <= 19'd0;
		WeightsStore8[216] <= 19'd0;
		WeightsStore8[217] <= 19'd0;
		WeightsStore8[218] <= 19'd0;
		WeightsStore8[219] <= 19'd0;
		WeightsStore8[220] <= 19'd0;
		WeightsStore8[221] <= 19'd0;
		WeightsStore8[222] <= 19'd0;
		WeightsStore8[223] <= 19'd0;
		WeightsStore8[224] <= 19'd0;
		WeightsStore8[225] <= 19'd0;
		WeightsStore8[226] <= 19'd0;
		WeightsStore8[227] <= 19'd0;
		WeightsStore8[228] <= 19'd0;
		WeightsStore8[229] <= 19'd0;
		WeightsStore8[230] <= 19'd0;
		WeightsStore8[231] <= 19'd0;
		WeightsStore8[232] <= 19'd0;
		WeightsStore8[233] <= 19'd0;
		WeightsStore8[234] <= 19'd0;
		WeightsStore8[235] <= 19'd0;
		WeightsStore8[236] <= 19'd0;
		WeightsStore8[237] <= 19'd0;
		WeightsStore8[238] <= 19'd0;
		WeightsStore8[239] <= 19'd0;
		WeightsStore8[240] <= 19'd0;
		WeightsStore8[241] <= 19'd0;
		WeightsStore8[242] <= 19'd0;
		WeightsStore8[243] <= 19'd0;
		WeightsStore8[244] <= 19'd0;
		WeightsStore8[245] <= 19'd0;
		WeightsStore8[246] <= 19'd0;
		WeightsStore8[247] <= 19'd0;
		WeightsStore8[248] <= 19'd0;
		WeightsStore8[249] <= 19'd0;
		WeightsStore8[250] <= 19'd0;
		WeightsStore8[251] <= 19'd0;
		WeightsStore8[252] <= 19'd0;
		WeightsStore8[253] <= 19'd0;
		WeightsStore8[254] <= 19'd0;
		WeightsStore8[255] <= 19'd0;
		WeightsStore8[256] <= 19'd0;
		WeightsStore8[257] <= 19'd0;
		WeightsStore8[258] <= 19'd0;
		WeightsStore8[259] <= 19'd0;
		WeightsStore8[260] <= 19'd0;
		WeightsStore8[261] <= 19'd0;
		WeightsStore8[262] <= 19'd0;
		WeightsStore8[263] <= 19'd0;
		WeightsStore8[264] <= 19'd0;
		WeightsStore8[265] <= 19'd0;
		WeightsStore8[266] <= 19'd0;
		WeightsStore8[267] <= 19'd0;
		WeightsStore8[268] <= 19'd0;
		WeightsStore8[269] <= 19'd0;
		WeightsStore8[270] <= 19'd0;
		WeightsStore8[271] <= 19'd0;
		WeightsStore8[272] <= 19'd0;
		WeightsStore8[273] <= 19'd0;
		WeightsStore8[274] <= 19'd0;
		WeightsStore8[275] <= 19'd0;
		WeightsStore8[276] <= 19'd0;
		WeightsStore8[277] <= 19'd0;
		WeightsStore8[278] <= 19'd0;
		WeightsStore8[279] <= 19'd0;
		WeightsStore8[280] <= 19'd0;
		WeightsStore8[281] <= 19'd0;
		WeightsStore8[282] <= 19'd0;
		WeightsStore8[283] <= 19'd0;
		WeightsStore8[284] <= 19'd0;
		WeightsStore8[285] <= 19'd0;
		WeightsStore8[286] <= 19'd0;
		WeightsStore8[287] <= 19'd0;
		WeightsStore8[288] <= 19'd0;
		WeightsStore8[289] <= 19'd0;
		WeightsStore8[290] <= 19'd0;
		WeightsStore8[291] <= 19'd0;
		WeightsStore8[292] <= 19'd0;
		WeightsStore8[293] <= 19'd0;
		WeightsStore8[294] <= 19'd0;
		WeightsStore8[295] <= 19'd0;
		WeightsStore8[296] <= 19'd0;
		WeightsStore8[297] <= 19'd0;
		WeightsStore8[298] <= 19'd0;
		WeightsStore8[299] <= 19'd0;
		WeightsStore8[300] <= 19'd0;
		WeightsStore8[301] <= 19'd0;
		WeightsStore8[302] <= 19'd0;
		WeightsStore8[303] <= 19'd0;
		WeightsStore8[304] <= 19'd0;
		WeightsStore8[305] <= 19'd0;
		WeightsStore8[306] <= 19'd0;
		WeightsStore8[307] <= 19'd0;
		WeightsStore8[308] <= 19'd0;
		WeightsStore8[309] <= 19'd0;
		WeightsStore8[310] <= 19'd0;
		WeightsStore8[311] <= 19'd0;
		WeightsStore8[312] <= 19'd0;
		WeightsStore8[313] <= 19'd0;
		WeightsStore8[314] <= 19'd0;
		WeightsStore8[315] <= 19'd0;
		WeightsStore8[316] <= 19'd0;
		WeightsStore8[317] <= 19'd0;
		WeightsStore8[318] <= 19'd0;
		WeightsStore8[319] <= 19'd0;
		WeightsStore8[320] <= 19'd0;
		WeightsStore8[321] <= 19'd0;
		WeightsStore8[322] <= 19'd0;
		WeightsStore8[323] <= 19'd0;
		WeightsStore8[324] <= 19'd0;
		WeightsStore8[325] <= 19'd0;
		WeightsStore8[326] <= 19'd0;
		WeightsStore8[327] <= 19'd0;
		WeightsStore8[328] <= 19'd0;
		WeightsStore8[329] <= 19'd0;
		WeightsStore8[330] <= 19'd0;
		WeightsStore8[331] <= 19'd0;
		WeightsStore8[332] <= 19'd0;
		WeightsStore8[333] <= 19'd0;
		WeightsStore8[334] <= 19'd0;
		WeightsStore8[335] <= 19'd0;
		WeightsStore8[336] <= 19'd0;
		WeightsStore8[337] <= 19'd0;
		WeightsStore8[338] <= 19'd0;
		WeightsStore8[339] <= 19'd0;
		WeightsStore8[340] <= 19'd0;
		WeightsStore8[341] <= 19'd0;
		WeightsStore8[342] <= 19'd0;
		WeightsStore8[343] <= 19'd0;
		WeightsStore8[344] <= 19'd0;
		WeightsStore8[345] <= 19'd0;
		WeightsStore8[346] <= 19'd0;
		WeightsStore8[347] <= 19'd0;
		WeightsStore8[348] <= 19'd0;
		WeightsStore8[349] <= 19'd0;
		WeightsStore8[350] <= 19'd0;
		WeightsStore8[351] <= 19'd0;
		WeightsStore8[352] <= 19'd0;
		WeightsStore8[353] <= 19'd0;
		WeightsStore8[354] <= 19'd0;
		WeightsStore8[355] <= 19'd0;
		WeightsStore8[356] <= 19'd0;
		WeightsStore8[357] <= 19'd0;
		WeightsStore8[358] <= 19'd0;
		WeightsStore8[359] <= 19'd0;
		WeightsStore8[360] <= 19'd0;
		WeightsStore8[361] <= 19'd0;
		WeightsStore8[362] <= 19'd0;
		WeightsStore8[363] <= 19'd0;
		WeightsStore8[364] <= 19'd0;
		WeightsStore8[365] <= 19'd0;
		WeightsStore8[366] <= 19'd0;
		WeightsStore8[367] <= 19'd0;
		WeightsStore8[368] <= 19'd0;
		WeightsStore8[369] <= 19'd0;
		WeightsStore8[370] <= 19'd0;
		WeightsStore8[371] <= 19'd0;
		WeightsStore8[372] <= 19'd0;
		WeightsStore8[373] <= 19'd0;
		WeightsStore8[374] <= 19'd0;
		WeightsStore8[375] <= 19'd0;
		WeightsStore8[376] <= 19'd0;
		WeightsStore8[377] <= 19'd0;
		WeightsStore8[378] <= 19'd0;
		WeightsStore8[379] <= 19'd0;
		WeightsStore8[380] <= 19'd0;
		WeightsStore8[381] <= 19'd0;
		WeightsStore8[382] <= 19'd0;
		WeightsStore8[383] <= 19'd0;
		WeightsStore8[384] <= 19'd0;
		WeightsStore8[385] <= 19'd0;
		WeightsStore8[386] <= 19'd0;
		WeightsStore8[387] <= 19'd0;
		WeightsStore8[388] <= 19'd0;
		WeightsStore8[389] <= 19'd0;
		WeightsStore8[390] <= 19'd0;
		WeightsStore8[391] <= 19'd0;
		WeightsStore8[392] <= 19'd0;
		WeightsStore8[393] <= 19'd0;
		WeightsStore8[394] <= 19'd0;
		WeightsStore8[395] <= 19'd0;
		WeightsStore8[396] <= 19'd0;
		WeightsStore8[397] <= 19'd0;
		WeightsStore8[398] <= 19'd0;
		WeightsStore8[399] <= 19'd0;
		WeightsStore8[400] <= 19'd0;
		WeightsStore8[401] <= 19'd0;
		WeightsStore8[402] <= 19'd0;
		WeightsStore8[403] <= 19'd0;
		WeightsStore8[404] <= 19'd0;
		WeightsStore8[405] <= 19'd0;
		WeightsStore8[406] <= 19'd0;
		WeightsStore8[407] <= 19'd0;
		WeightsStore8[408] <= 19'd0;
		WeightsStore8[409] <= 19'd0;
		WeightsStore8[410] <= 19'd0;
		WeightsStore8[411] <= 19'd0;
		WeightsStore8[412] <= 19'd0;
		WeightsStore8[413] <= 19'd0;
		WeightsStore8[414] <= 19'd0;
		WeightsStore8[415] <= 19'd0;
		WeightsStore8[416] <= 19'd0;
		WeightsStore8[417] <= 19'd0;
		WeightsStore8[418] <= 19'd0;
		WeightsStore8[419] <= 19'd0;
		WeightsStore8[420] <= 19'd0;
		WeightsStore8[421] <= 19'd0;
		WeightsStore8[422] <= 19'd0;
		WeightsStore8[423] <= 19'd0;
		WeightsStore8[424] <= 19'd0;
		WeightsStore8[425] <= 19'd0;
		WeightsStore8[426] <= 19'd0;
		WeightsStore8[427] <= 19'd0;
		WeightsStore8[428] <= 19'd0;
		WeightsStore8[429] <= 19'd0;
		WeightsStore8[430] <= 19'd0;
		WeightsStore8[431] <= 19'd0;
		WeightsStore8[432] <= 19'd0;
		WeightsStore8[433] <= 19'd0;
		WeightsStore8[434] <= 19'd0;
		WeightsStore8[435] <= 19'd0;
		WeightsStore8[436] <= 19'd0;
		WeightsStore8[437] <= 19'd0;
		WeightsStore8[438] <= 19'd0;
		WeightsStore8[439] <= 19'd0;
		WeightsStore8[440] <= 19'd0;
		WeightsStore8[441] <= 19'd0;
		WeightsStore8[442] <= 19'd0;
		WeightsStore8[443] <= 19'd0;
		WeightsStore8[444] <= 19'd0;
		WeightsStore8[445] <= 19'd0;
		WeightsStore8[446] <= 19'd0;
		WeightsStore8[447] <= 19'd0;
		WeightsStore8[448] <= 19'd0;
		WeightsStore8[449] <= 19'd0;
		WeightsStore8[450] <= 19'd0;
		WeightsStore8[451] <= 19'd0;
		WeightsStore8[452] <= 19'd0;
		WeightsStore8[453] <= 19'd0;
		WeightsStore8[454] <= 19'd0;
		WeightsStore8[455] <= 19'd0;
		WeightsStore8[456] <= 19'd0;
		WeightsStore8[457] <= 19'd0;
		WeightsStore8[458] <= 19'd0;
		WeightsStore8[459] <= 19'd0;
		WeightsStore8[460] <= 19'd0;
		WeightsStore8[461] <= 19'd0;
		WeightsStore8[462] <= 19'd0;
		WeightsStore8[463] <= 19'd0;
		WeightsStore8[464] <= 19'd0;
		WeightsStore8[465] <= 19'd0;
		WeightsStore8[466] <= 19'd0;
		WeightsStore8[467] <= 19'd0;
		WeightsStore8[468] <= 19'd0;
		WeightsStore8[469] <= 19'd0;
		WeightsStore8[470] <= 19'd0;
		WeightsStore8[471] <= 19'd0;
		WeightsStore8[472] <= 19'd0;
		WeightsStore8[473] <= 19'd0;
		WeightsStore8[474] <= 19'd0;
		WeightsStore8[475] <= 19'd0;
		WeightsStore8[476] <= 19'd0;
		WeightsStore8[477] <= 19'd0;
		WeightsStore8[478] <= 19'd0;
		WeightsStore8[479] <= 19'd0;
		WeightsStore8[480] <= 19'd0;
		WeightsStore8[481] <= 19'd0;
		WeightsStore8[482] <= 19'd0;
		WeightsStore8[483] <= 19'd0;
		WeightsStore8[484] <= 19'd0;
		WeightsStore8[485] <= 19'd0;
		WeightsStore8[486] <= 19'd0;
		WeightsStore8[487] <= 19'd0;
		WeightsStore8[488] <= 19'd0;
		WeightsStore8[489] <= 19'd0;
		WeightsStore8[490] <= 19'd0;
		WeightsStore8[491] <= 19'd0;
		WeightsStore8[492] <= 19'd0;
		WeightsStore8[493] <= 19'd0;
		WeightsStore8[494] <= 19'd0;
		WeightsStore8[495] <= 19'd0;
		WeightsStore8[496] <= 19'd0;
		WeightsStore8[497] <= 19'd0;
		WeightsStore8[498] <= 19'd0;
		WeightsStore8[499] <= 19'd0;
		WeightsStore8[500] <= 19'd0;
		WeightsStore8[501] <= 19'd0;
		WeightsStore8[502] <= 19'd0;
		WeightsStore8[503] <= 19'd0;
		WeightsStore8[504] <= 19'd0;
		WeightsStore8[505] <= 19'd0;
		WeightsStore8[506] <= 19'd0;
		WeightsStore8[507] <= 19'd0;
		WeightsStore8[508] <= 19'd0;
		WeightsStore8[509] <= 19'd0;
		WeightsStore8[510] <= 19'd0;
		WeightsStore8[511] <= 19'd0;
		WeightsStore8[512] <= 19'd0;
		WeightsStore8[513] <= 19'd0;
		WeightsStore8[514] <= 19'd0;
		WeightsStore8[515] <= 19'd0;
		WeightsStore8[516] <= 19'd0;
		WeightsStore8[517] <= 19'd0;
		WeightsStore8[518] <= 19'd0;
		WeightsStore8[519] <= 19'd0;
		WeightsStore8[520] <= 19'd0;
		WeightsStore8[521] <= 19'd0;
		WeightsStore8[522] <= 19'd0;
		WeightsStore8[523] <= 19'd0;
		WeightsStore8[524] <= 19'd0;
		WeightsStore8[525] <= 19'd0;
		WeightsStore8[526] <= 19'd0;
		WeightsStore8[527] <= 19'd0;
		WeightsStore8[528] <= 19'd0;
		WeightsStore8[529] <= 19'd0;
		WeightsStore8[530] <= 19'd0;
		WeightsStore8[531] <= 19'd0;
		WeightsStore8[532] <= 19'd0;
		WeightsStore8[533] <= 19'd0;
		WeightsStore8[534] <= 19'd0;
		WeightsStore8[535] <= 19'd0;
		WeightsStore8[536] <= 19'd0;
		WeightsStore8[537] <= 19'd0;
		WeightsStore8[538] <= 19'd0;
		WeightsStore8[539] <= 19'd0;
		WeightsStore8[540] <= 19'd0;
		WeightsStore8[541] <= 19'd0;
		WeightsStore8[542] <= 19'd0;
		WeightsStore8[543] <= 19'd0;
		WeightsStore8[544] <= 19'd0;
		WeightsStore8[545] <= 19'd0;
		WeightsStore8[546] <= 19'd0;
		WeightsStore8[547] <= 19'd0;
		WeightsStore8[548] <= 19'd0;
		WeightsStore8[549] <= 19'd0;
		WeightsStore8[550] <= 19'd0;
		WeightsStore8[551] <= 19'd0;
		WeightsStore8[552] <= 19'd0;
		WeightsStore8[553] <= 19'd0;
		WeightsStore8[554] <= 19'd0;
		WeightsStore8[555] <= 19'd0;
		WeightsStore8[556] <= 19'd0;
		WeightsStore8[557] <= 19'd0;
		WeightsStore8[558] <= 19'd0;
		WeightsStore8[559] <= 19'd0;
		WeightsStore8[560] <= 19'd0;
		WeightsStore8[561] <= 19'd0;
		WeightsStore8[562] <= 19'd0;
		WeightsStore8[563] <= 19'd0;
		WeightsStore8[564] <= 19'd0;
		WeightsStore8[565] <= 19'd0;
		WeightsStore8[566] <= 19'd0;
		WeightsStore8[567] <= 19'd0;
		WeightsStore8[568] <= 19'd0;
		WeightsStore8[569] <= 19'd0;
		WeightsStore8[570] <= 19'd0;
		WeightsStore8[571] <= 19'd0;
		WeightsStore8[572] <= 19'd0;
		WeightsStore8[573] <= 19'd0;
		WeightsStore8[574] <= 19'd0;
		WeightsStore8[575] <= 19'd0;
		WeightsStore8[576] <= 19'd0;
		WeightsStore8[577] <= 19'd0;
		WeightsStore8[578] <= 19'd0;
		WeightsStore8[579] <= 19'd0;
		WeightsStore8[580] <= 19'd0;
		WeightsStore8[581] <= 19'd0;
		WeightsStore8[582] <= 19'd0;
		WeightsStore8[583] <= 19'd0;
		WeightsStore8[584] <= 19'd0;
		WeightsStore8[585] <= 19'd0;
		WeightsStore8[586] <= 19'd0;
		WeightsStore8[587] <= 19'd0;
		WeightsStore8[588] <= 19'd0;
		WeightsStore8[589] <= 19'd0;
		WeightsStore8[590] <= 19'd0;
		WeightsStore8[591] <= 19'd0;
		WeightsStore8[592] <= 19'd0;
		WeightsStore8[593] <= 19'd0;
		WeightsStore8[594] <= 19'd0;
		WeightsStore8[595] <= 19'd0;
		WeightsStore8[596] <= 19'd0;
		WeightsStore8[597] <= 19'd0;
		WeightsStore8[598] <= 19'd0;
		WeightsStore8[599] <= 19'd0;
		WeightsStore8[600] <= 19'd0;
		WeightsStore8[601] <= 19'd0;
		WeightsStore8[602] <= 19'd0;
		WeightsStore8[603] <= 19'd0;
		WeightsStore8[604] <= 19'd0;
		WeightsStore8[605] <= 19'd0;
		WeightsStore8[606] <= 19'd0;
		WeightsStore8[607] <= 19'd0;
		WeightsStore8[608] <= 19'd0;
		WeightsStore8[609] <= 19'd0;
		WeightsStore8[610] <= 19'd0;
		WeightsStore8[611] <= 19'd0;
		WeightsStore8[612] <= 19'd0;
		WeightsStore8[613] <= 19'd0;
		WeightsStore8[614] <= 19'd0;
		WeightsStore8[615] <= 19'd0;
		WeightsStore8[616] <= 19'd0;
		WeightsStore8[617] <= 19'd0;
		WeightsStore8[618] <= 19'd0;
		WeightsStore8[619] <= 19'd0;
		WeightsStore8[620] <= 19'd0;
		WeightsStore8[621] <= 19'd0;
		WeightsStore8[622] <= 19'd0;
		WeightsStore8[623] <= 19'd0;
		WeightsStore8[624] <= 19'd0;
		WeightsStore8[625] <= 19'd0;
		WeightsStore8[626] <= 19'd0;
		WeightsStore8[627] <= 19'd0;
		WeightsStore8[628] <= 19'd0;
		WeightsStore8[629] <= 19'd0;
		WeightsStore8[630] <= 19'd0;
		WeightsStore8[631] <= 19'd0;
		WeightsStore8[632] <= 19'd0;
		WeightsStore8[633] <= 19'd0;
		WeightsStore8[634] <= 19'd0;
		WeightsStore8[635] <= 19'd0;
		WeightsStore8[636] <= 19'd0;
		WeightsStore8[637] <= 19'd0;
		WeightsStore8[638] <= 19'd0;
		WeightsStore8[639] <= 19'd0;
		WeightsStore8[640] <= 19'd0;
		WeightsStore8[641] <= 19'd0;
		WeightsStore8[642] <= 19'd0;
		WeightsStore8[643] <= 19'd0;
		WeightsStore8[644] <= 19'd0;
		WeightsStore8[645] <= 19'd0;
		WeightsStore8[646] <= 19'd0;
		WeightsStore8[647] <= 19'd0;
		WeightsStore8[648] <= 19'd0;
		WeightsStore8[649] <= 19'd0;
		WeightsStore8[650] <= 19'd0;
		WeightsStore8[651] <= 19'd0;
		WeightsStore8[652] <= 19'd0;
		WeightsStore8[653] <= 19'd0;
		WeightsStore8[654] <= 19'd0;
		WeightsStore8[655] <= 19'd0;
		WeightsStore8[656] <= 19'd0;
		WeightsStore8[657] <= 19'd0;
		WeightsStore8[658] <= 19'd0;
		WeightsStore8[659] <= 19'd0;
		WeightsStore8[660] <= 19'd0;
		WeightsStore8[661] <= 19'd0;
		WeightsStore8[662] <= 19'd0;
		WeightsStore8[663] <= 19'd0;
		WeightsStore8[664] <= 19'd0;
		WeightsStore8[665] <= 19'd0;
		WeightsStore8[666] <= 19'd0;
		WeightsStore8[667] <= 19'd0;
		WeightsStore8[668] <= 19'd0;
		WeightsStore8[669] <= 19'd0;
		WeightsStore8[670] <= 19'd0;
		WeightsStore8[671] <= 19'd0;
		WeightsStore8[672] <= 19'd0;
		WeightsStore8[673] <= 19'd0;
		WeightsStore8[674] <= 19'd0;
		WeightsStore8[675] <= 19'd0;
		WeightsStore8[676] <= 19'd0;
		WeightsStore8[677] <= 19'd0;
		WeightsStore8[678] <= 19'd0;
		WeightsStore8[679] <= 19'd0;
		WeightsStore8[680] <= 19'd0;
		WeightsStore8[681] <= 19'd0;
		WeightsStore8[682] <= 19'd0;
		WeightsStore8[683] <= 19'd0;
		WeightsStore8[684] <= 19'd0;
		WeightsStore8[685] <= 19'd0;
		WeightsStore8[686] <= 19'd0;
		WeightsStore8[687] <= 19'd0;
		WeightsStore8[688] <= 19'd0;
		WeightsStore8[689] <= 19'd0;
		WeightsStore8[690] <= 19'd0;
		WeightsStore8[691] <= 19'd0;
		WeightsStore8[692] <= 19'd0;
		WeightsStore8[693] <= 19'd0;
		WeightsStore8[694] <= 19'd0;
		WeightsStore8[695] <= 19'd0;
		WeightsStore8[696] <= 19'd0;
		WeightsStore8[697] <= 19'd0;
		WeightsStore8[698] <= 19'd0;
		WeightsStore8[699] <= 19'd0;
		WeightsStore8[700] <= 19'd0;
		WeightsStore8[701] <= 19'd0;
		WeightsStore8[702] <= 19'd0;
		WeightsStore8[703] <= 19'd0;
		WeightsStore8[704] <= 19'd0;
		WeightsStore8[705] <= 19'd0;
		WeightsStore8[706] <= 19'd0;
		WeightsStore8[707] <= 19'd0;
		WeightsStore8[708] <= 19'd0;
		WeightsStore8[709] <= 19'd0;
		WeightsStore8[710] <= 19'd0;
		WeightsStore8[711] <= 19'd0;
		WeightsStore8[712] <= 19'd0;
		WeightsStore8[713] <= 19'd0;
		WeightsStore8[714] <= 19'd0;
		WeightsStore8[715] <= 19'd0;
		WeightsStore8[716] <= 19'd0;
		WeightsStore8[717] <= 19'd0;
		WeightsStore8[718] <= 19'd0;
		WeightsStore8[719] <= 19'd0;
		WeightsStore8[720] <= 19'd0;
		WeightsStore8[721] <= 19'd0;
		WeightsStore8[722] <= 19'd0;
		WeightsStore8[723] <= 19'd0;
		WeightsStore8[724] <= 19'd0;
		WeightsStore8[725] <= 19'd0;
		WeightsStore8[726] <= 19'd0;
		WeightsStore8[727] <= 19'd0;
		WeightsStore8[728] <= 19'd0;
		WeightsStore8[729] <= 19'd0;
		WeightsStore8[730] <= 19'd0;
		WeightsStore8[731] <= 19'd0;
		WeightsStore8[732] <= 19'd0;
		WeightsStore8[733] <= 19'd0;
		WeightsStore8[734] <= 19'd0;
		WeightsStore8[735] <= 19'd0;
		WeightsStore8[736] <= 19'd0;
		WeightsStore8[737] <= 19'd0;
		WeightsStore8[738] <= 19'd0;
		WeightsStore8[739] <= 19'd0;
		WeightsStore8[740] <= 19'd0;
		WeightsStore8[741] <= 19'd0;
		WeightsStore8[742] <= 19'd0;
		WeightsStore8[743] <= 19'd0;
		WeightsStore8[744] <= 19'd0;
		WeightsStore8[745] <= 19'd0;
		WeightsStore8[746] <= 19'd0;
		WeightsStore8[747] <= 19'd0;
		WeightsStore8[748] <= 19'd0;
		WeightsStore8[749] <= 19'd0;
		WeightsStore8[750] <= 19'd0;
		WeightsStore8[751] <= 19'd0;
		WeightsStore8[752] <= 19'd0;
		WeightsStore8[753] <= 19'd0;
		WeightsStore8[754] <= 19'd0;
		WeightsStore8[755] <= 19'd0;
		WeightsStore8[756] <= 19'd0;
		WeightsStore8[757] <= 19'd0;
		WeightsStore8[758] <= 19'd0;
		WeightsStore8[759] <= 19'd0;
		WeightsStore8[760] <= 19'd0;
		WeightsStore8[761] <= 19'd0;
		WeightsStore8[762] <= 19'd0;
		WeightsStore8[763] <= 19'd0;
		WeightsStore8[764] <= 19'd0;
		WeightsStore8[765] <= 19'd0;
		WeightsStore8[766] <= 19'd0;
		WeightsStore8[767] <= 19'd0;
		WeightsStore8[768] <= 19'd0;
		WeightsStore8[769] <= 19'd0;
		WeightsStore8[770] <= 19'd0;
		WeightsStore8[771] <= 19'd0;
		WeightsStore8[772] <= 19'd0;
		WeightsStore8[773] <= 19'd0;
		WeightsStore8[774] <= 19'd0;
		WeightsStore8[775] <= 19'd0;
		WeightsStore8[776] <= 19'd0;
		WeightsStore8[777] <= 19'd0;
		WeightsStore8[778] <= 19'd0;
		WeightsStore8[779] <= 19'd0;
		WeightsStore8[780] <= 19'd0;
		WeightsStore8[781] <= 19'd0;
		WeightsStore8[782] <= 19'd0;
		WeightsStore8[783] <= 19'd0;
		WeightsStore8[784] <= 19'd0;
		WeightsStore9[0] <= 19'd0;
		WeightsStore9[1] <= 19'd0;
		WeightsStore9[2] <= 19'd0;
		WeightsStore9[3] <= 19'd0;
		WeightsStore9[4] <= 19'd0;
		WeightsStore9[5] <= 19'd0;
		WeightsStore9[6] <= 19'd0;
		WeightsStore9[7] <= 19'd0;
		WeightsStore9[8] <= 19'd0;
		WeightsStore9[9] <= 19'd0;
		WeightsStore9[10] <= 19'd0;
		WeightsStore9[11] <= 19'd0;
		WeightsStore9[12] <= 19'd0;
		WeightsStore9[13] <= 19'd0;
		WeightsStore9[14] <= 19'd0;
		WeightsStore9[15] <= 19'd0;
		WeightsStore9[16] <= 19'd0;
		WeightsStore9[17] <= 19'd0;
		WeightsStore9[18] <= 19'd0;
		WeightsStore9[19] <= 19'd0;
		WeightsStore9[20] <= 19'd0;
		WeightsStore9[21] <= 19'd0;
		WeightsStore9[22] <= 19'd0;
		WeightsStore9[23] <= 19'd0;
		WeightsStore9[24] <= 19'd0;
		WeightsStore9[25] <= 19'd0;
		WeightsStore9[26] <= 19'd0;
		WeightsStore9[27] <= 19'd0;
		WeightsStore9[28] <= 19'd0;
		WeightsStore9[29] <= 19'd0;
		WeightsStore9[30] <= 19'd0;
		WeightsStore9[31] <= 19'd0;
		WeightsStore9[32] <= 19'd0;
		WeightsStore9[33] <= 19'd0;
		WeightsStore9[34] <= 19'd0;
		WeightsStore9[35] <= 19'd0;
		WeightsStore9[36] <= 19'd0;
		WeightsStore9[37] <= 19'd0;
		WeightsStore9[38] <= 19'd0;
		WeightsStore9[39] <= 19'd0;
		WeightsStore9[40] <= 19'd0;
		WeightsStore9[41] <= 19'd0;
		WeightsStore9[42] <= 19'd0;
		WeightsStore9[43] <= 19'd0;
		WeightsStore9[44] <= 19'd0;
		WeightsStore9[45] <= 19'd0;
		WeightsStore9[46] <= 19'd0;
		WeightsStore9[47] <= 19'd0;
		WeightsStore9[48] <= 19'd0;
		WeightsStore9[49] <= 19'd0;
		WeightsStore9[50] <= 19'd0;
		WeightsStore9[51] <= 19'd0;
		WeightsStore9[52] <= 19'd0;
		WeightsStore9[53] <= 19'd0;
		WeightsStore9[54] <= 19'd0;
		WeightsStore9[55] <= 19'd0;
		WeightsStore9[56] <= 19'd0;
		WeightsStore9[57] <= 19'd0;
		WeightsStore9[58] <= 19'd0;
		WeightsStore9[59] <= 19'd0;
		WeightsStore9[60] <= 19'd0;
		WeightsStore9[61] <= 19'd0;
		WeightsStore9[62] <= 19'd0;
		WeightsStore9[63] <= 19'd0;
		WeightsStore9[64] <= 19'd0;
		WeightsStore9[65] <= 19'd0;
		WeightsStore9[66] <= 19'd0;
		WeightsStore9[67] <= 19'd0;
		WeightsStore9[68] <= 19'd0;
		WeightsStore9[69] <= 19'd0;
		WeightsStore9[70] <= 19'd0;
		WeightsStore9[71] <= 19'd0;
		WeightsStore9[72] <= 19'd0;
		WeightsStore9[73] <= 19'd0;
		WeightsStore9[74] <= 19'd0;
		WeightsStore9[75] <= 19'd0;
		WeightsStore9[76] <= 19'd0;
		WeightsStore9[77] <= 19'd0;
		WeightsStore9[78] <= 19'd0;
		WeightsStore9[79] <= 19'd0;
		WeightsStore9[80] <= 19'd0;
		WeightsStore9[81] <= 19'd0;
		WeightsStore9[82] <= 19'd0;
		WeightsStore9[83] <= 19'd0;
		WeightsStore9[84] <= 19'd0;
		WeightsStore9[85] <= 19'd0;
		WeightsStore9[86] <= 19'd0;
		WeightsStore9[87] <= 19'd0;
		WeightsStore9[88] <= 19'd0;
		WeightsStore9[89] <= 19'd0;
		WeightsStore9[90] <= 19'd0;
		WeightsStore9[91] <= 19'd0;
		WeightsStore9[92] <= 19'd0;
		WeightsStore9[93] <= 19'd0;
		WeightsStore9[94] <= 19'd0;
		WeightsStore9[95] <= 19'd0;
		WeightsStore9[96] <= 19'd0;
		WeightsStore9[97] <= 19'd0;
		WeightsStore9[98] <= 19'd0;
		WeightsStore9[99] <= 19'd0;
		WeightsStore9[100] <= 19'd0;
		WeightsStore9[101] <= 19'd0;
		WeightsStore9[102] <= 19'd0;
		WeightsStore9[103] <= 19'd0;
		WeightsStore9[104] <= 19'd0;
		WeightsStore9[105] <= 19'd0;
		WeightsStore9[106] <= 19'd0;
		WeightsStore9[107] <= 19'd0;
		WeightsStore9[108] <= 19'd0;
		WeightsStore9[109] <= 19'd0;
		WeightsStore9[110] <= 19'd0;
		WeightsStore9[111] <= 19'd0;
		WeightsStore9[112] <= 19'd0;
		WeightsStore9[113] <= 19'd0;
		WeightsStore9[114] <= 19'd0;
		WeightsStore9[115] <= 19'd0;
		WeightsStore9[116] <= 19'd0;
		WeightsStore9[117] <= 19'd0;
		WeightsStore9[118] <= 19'd0;
		WeightsStore9[119] <= 19'd0;
		WeightsStore9[120] <= 19'd0;
		WeightsStore9[121] <= 19'd0;
		WeightsStore9[122] <= 19'd0;
		WeightsStore9[123] <= 19'd0;
		WeightsStore9[124] <= 19'd0;
		WeightsStore9[125] <= 19'd0;
		WeightsStore9[126] <= 19'd0;
		WeightsStore9[127] <= 19'd0;
		WeightsStore9[128] <= 19'd0;
		WeightsStore9[129] <= 19'd0;
		WeightsStore9[130] <= 19'd0;
		WeightsStore9[131] <= 19'd0;
		WeightsStore9[132] <= 19'd0;
		WeightsStore9[133] <= 19'd0;
		WeightsStore9[134] <= 19'd0;
		WeightsStore9[135] <= 19'd0;
		WeightsStore9[136] <= 19'd0;
		WeightsStore9[137] <= 19'd0;
		WeightsStore9[138] <= 19'd0;
		WeightsStore9[139] <= 19'd0;
		WeightsStore9[140] <= 19'd0;
		WeightsStore9[141] <= 19'd0;
		WeightsStore9[142] <= 19'd0;
		WeightsStore9[143] <= 19'd0;
		WeightsStore9[144] <= 19'd0;
		WeightsStore9[145] <= 19'd0;
		WeightsStore9[146] <= 19'd0;
		WeightsStore9[147] <= 19'd0;
		WeightsStore9[148] <= 19'd0;
		WeightsStore9[149] <= 19'd0;
		WeightsStore9[150] <= 19'd0;
		WeightsStore9[151] <= 19'd0;
		WeightsStore9[152] <= 19'd0;
		WeightsStore9[153] <= 19'd0;
		WeightsStore9[154] <= 19'd0;
		WeightsStore9[155] <= 19'd0;
		WeightsStore9[156] <= 19'd0;
		WeightsStore9[157] <= 19'd0;
		WeightsStore9[158] <= 19'd0;
		WeightsStore9[159] <= 19'd0;
		WeightsStore9[160] <= 19'd0;
		WeightsStore9[161] <= 19'd0;
		WeightsStore9[162] <= 19'd0;
		WeightsStore9[163] <= 19'd0;
		WeightsStore9[164] <= 19'd0;
		WeightsStore9[165] <= 19'd0;
		WeightsStore9[166] <= 19'd0;
		WeightsStore9[167] <= 19'd0;
		WeightsStore9[168] <= 19'd0;
		WeightsStore9[169] <= 19'd0;
		WeightsStore9[170] <= 19'd0;
		WeightsStore9[171] <= 19'd0;
		WeightsStore9[172] <= 19'd0;
		WeightsStore9[173] <= 19'd0;
		WeightsStore9[174] <= 19'd0;
		WeightsStore9[175] <= 19'd0;
		WeightsStore9[176] <= 19'd0;
		WeightsStore9[177] <= 19'd0;
		WeightsStore9[178] <= 19'd0;
		WeightsStore9[179] <= 19'd0;
		WeightsStore9[180] <= 19'd0;
		WeightsStore9[181] <= 19'd0;
		WeightsStore9[182] <= 19'd0;
		WeightsStore9[183] <= 19'd0;
		WeightsStore9[184] <= 19'd0;
		WeightsStore9[185] <= 19'd0;
		WeightsStore9[186] <= 19'd0;
		WeightsStore9[187] <= 19'd0;
		WeightsStore9[188] <= 19'd0;
		WeightsStore9[189] <= 19'd0;
		WeightsStore9[190] <= 19'd0;
		WeightsStore9[191] <= 19'd0;
		WeightsStore9[192] <= 19'd0;
		WeightsStore9[193] <= 19'd0;
		WeightsStore9[194] <= 19'd0;
		WeightsStore9[195] <= 19'd0;
		WeightsStore9[196] <= 19'd0;
		WeightsStore9[197] <= 19'd0;
		WeightsStore9[198] <= 19'd0;
		WeightsStore9[199] <= 19'd0;
		WeightsStore9[200] <= 19'd0;
		WeightsStore9[201] <= 19'd0;
		WeightsStore9[202] <= 19'd0;
		WeightsStore9[203] <= 19'd0;
		WeightsStore9[204] <= 19'd0;
		WeightsStore9[205] <= 19'd0;
		WeightsStore9[206] <= 19'd0;
		WeightsStore9[207] <= 19'd0;
		WeightsStore9[208] <= 19'd0;
		WeightsStore9[209] <= 19'd0;
		WeightsStore9[210] <= 19'd0;
		WeightsStore9[211] <= 19'd0;
		WeightsStore9[212] <= 19'd0;
		WeightsStore9[213] <= 19'd0;
		WeightsStore9[214] <= 19'd0;
		WeightsStore9[215] <= 19'd0;
		WeightsStore9[216] <= 19'd0;
		WeightsStore9[217] <= 19'd0;
		WeightsStore9[218] <= 19'd0;
		WeightsStore9[219] <= 19'd0;
		WeightsStore9[220] <= 19'd0;
		WeightsStore9[221] <= 19'd0;
		WeightsStore9[222] <= 19'd0;
		WeightsStore9[223] <= 19'd0;
		WeightsStore9[224] <= 19'd0;
		WeightsStore9[225] <= 19'd0;
		WeightsStore9[226] <= 19'd0;
		WeightsStore9[227] <= 19'd0;
		WeightsStore9[228] <= 19'd0;
		WeightsStore9[229] <= 19'd0;
		WeightsStore9[230] <= 19'd0;
		WeightsStore9[231] <= 19'd0;
		WeightsStore9[232] <= 19'd0;
		WeightsStore9[233] <= 19'd0;
		WeightsStore9[234] <= 19'd0;
		WeightsStore9[235] <= 19'd0;
		WeightsStore9[236] <= 19'd0;
		WeightsStore9[237] <= 19'd0;
		WeightsStore9[238] <= 19'd0;
		WeightsStore9[239] <= 19'd0;
		WeightsStore9[240] <= 19'd0;
		WeightsStore9[241] <= 19'd0;
		WeightsStore9[242] <= 19'd0;
		WeightsStore9[243] <= 19'd0;
		WeightsStore9[244] <= 19'd0;
		WeightsStore9[245] <= 19'd0;
		WeightsStore9[246] <= 19'd0;
		WeightsStore9[247] <= 19'd0;
		WeightsStore9[248] <= 19'd0;
		WeightsStore9[249] <= 19'd0;
		WeightsStore9[250] <= 19'd0;
		WeightsStore9[251] <= 19'd0;
		WeightsStore9[252] <= 19'd0;
		WeightsStore9[253] <= 19'd0;
		WeightsStore9[254] <= 19'd0;
		WeightsStore9[255] <= 19'd0;
		WeightsStore9[256] <= 19'd0;
		WeightsStore9[257] <= 19'd0;
		WeightsStore9[258] <= 19'd0;
		WeightsStore9[259] <= 19'd0;
		WeightsStore9[260] <= 19'd0;
		WeightsStore9[261] <= 19'd0;
		WeightsStore9[262] <= 19'd0;
		WeightsStore9[263] <= 19'd0;
		WeightsStore9[264] <= 19'd0;
		WeightsStore9[265] <= 19'd0;
		WeightsStore9[266] <= 19'd0;
		WeightsStore9[267] <= 19'd0;
		WeightsStore9[268] <= 19'd0;
		WeightsStore9[269] <= 19'd0;
		WeightsStore9[270] <= 19'd0;
		WeightsStore9[271] <= 19'd0;
		WeightsStore9[272] <= 19'd0;
		WeightsStore9[273] <= 19'd0;
		WeightsStore9[274] <= 19'd0;
		WeightsStore9[275] <= 19'd0;
		WeightsStore9[276] <= 19'd0;
		WeightsStore9[277] <= 19'd0;
		WeightsStore9[278] <= 19'd0;
		WeightsStore9[279] <= 19'd0;
		WeightsStore9[280] <= 19'd0;
		WeightsStore9[281] <= 19'd0;
		WeightsStore9[282] <= 19'd0;
		WeightsStore9[283] <= 19'd0;
		WeightsStore9[284] <= 19'd0;
		WeightsStore9[285] <= 19'd0;
		WeightsStore9[286] <= 19'd0;
		WeightsStore9[287] <= 19'd0;
		WeightsStore9[288] <= 19'd0;
		WeightsStore9[289] <= 19'd0;
		WeightsStore9[290] <= 19'd0;
		WeightsStore9[291] <= 19'd0;
		WeightsStore9[292] <= 19'd0;
		WeightsStore9[293] <= 19'd0;
		WeightsStore9[294] <= 19'd0;
		WeightsStore9[295] <= 19'd0;
		WeightsStore9[296] <= 19'd0;
		WeightsStore9[297] <= 19'd0;
		WeightsStore9[298] <= 19'd0;
		WeightsStore9[299] <= 19'd0;
		WeightsStore9[300] <= 19'd0;
		WeightsStore9[301] <= 19'd0;
		WeightsStore9[302] <= 19'd0;
		WeightsStore9[303] <= 19'd0;
		WeightsStore9[304] <= 19'd0;
		WeightsStore9[305] <= 19'd0;
		WeightsStore9[306] <= 19'd0;
		WeightsStore9[307] <= 19'd0;
		WeightsStore9[308] <= 19'd0;
		WeightsStore9[309] <= 19'd0;
		WeightsStore9[310] <= 19'd0;
		WeightsStore9[311] <= 19'd0;
		WeightsStore9[312] <= 19'd0;
		WeightsStore9[313] <= 19'd0;
		WeightsStore9[314] <= 19'd0;
		WeightsStore9[315] <= 19'd0;
		WeightsStore9[316] <= 19'd0;
		WeightsStore9[317] <= 19'd0;
		WeightsStore9[318] <= 19'd0;
		WeightsStore9[319] <= 19'd0;
		WeightsStore9[320] <= 19'd0;
		WeightsStore9[321] <= 19'd0;
		WeightsStore9[322] <= 19'd0;
		WeightsStore9[323] <= 19'd0;
		WeightsStore9[324] <= 19'd0;
		WeightsStore9[325] <= 19'd0;
		WeightsStore9[326] <= 19'd0;
		WeightsStore9[327] <= 19'd0;
		WeightsStore9[328] <= 19'd0;
		WeightsStore9[329] <= 19'd0;
		WeightsStore9[330] <= 19'd0;
		WeightsStore9[331] <= 19'd0;
		WeightsStore9[332] <= 19'd0;
		WeightsStore9[333] <= 19'd0;
		WeightsStore9[334] <= 19'd0;
		WeightsStore9[335] <= 19'd0;
		WeightsStore9[336] <= 19'd0;
		WeightsStore9[337] <= 19'd0;
		WeightsStore9[338] <= 19'd0;
		WeightsStore9[339] <= 19'd0;
		WeightsStore9[340] <= 19'd0;
		WeightsStore9[341] <= 19'd0;
		WeightsStore9[342] <= 19'd0;
		WeightsStore9[343] <= 19'd0;
		WeightsStore9[344] <= 19'd0;
		WeightsStore9[345] <= 19'd0;
		WeightsStore9[346] <= 19'd0;
		WeightsStore9[347] <= 19'd0;
		WeightsStore9[348] <= 19'd0;
		WeightsStore9[349] <= 19'd0;
		WeightsStore9[350] <= 19'd0;
		WeightsStore9[351] <= 19'd0;
		WeightsStore9[352] <= 19'd0;
		WeightsStore9[353] <= 19'd0;
		WeightsStore9[354] <= 19'd0;
		WeightsStore9[355] <= 19'd0;
		WeightsStore9[356] <= 19'd0;
		WeightsStore9[357] <= 19'd0;
		WeightsStore9[358] <= 19'd0;
		WeightsStore9[359] <= 19'd0;
		WeightsStore9[360] <= 19'd0;
		WeightsStore9[361] <= 19'd0;
		WeightsStore9[362] <= 19'd0;
		WeightsStore9[363] <= 19'd0;
		WeightsStore9[364] <= 19'd0;
		WeightsStore9[365] <= 19'd0;
		WeightsStore9[366] <= 19'd0;
		WeightsStore9[367] <= 19'd0;
		WeightsStore9[368] <= 19'd0;
		WeightsStore9[369] <= 19'd0;
		WeightsStore9[370] <= 19'd0;
		WeightsStore9[371] <= 19'd0;
		WeightsStore9[372] <= 19'd0;
		WeightsStore9[373] <= 19'd0;
		WeightsStore9[374] <= 19'd0;
		WeightsStore9[375] <= 19'd0;
		WeightsStore9[376] <= 19'd0;
		WeightsStore9[377] <= 19'd0;
		WeightsStore9[378] <= 19'd0;
		WeightsStore9[379] <= 19'd0;
		WeightsStore9[380] <= 19'd0;
		WeightsStore9[381] <= 19'd0;
		WeightsStore9[382] <= 19'd0;
		WeightsStore9[383] <= 19'd0;
		WeightsStore9[384] <= 19'd0;
		WeightsStore9[385] <= 19'd0;
		WeightsStore9[386] <= 19'd0;
		WeightsStore9[387] <= 19'd0;
		WeightsStore9[388] <= 19'd0;
		WeightsStore9[389] <= 19'd0;
		WeightsStore9[390] <= 19'd0;
		WeightsStore9[391] <= 19'd0;
		WeightsStore9[392] <= 19'd0;
		WeightsStore9[393] <= 19'd0;
		WeightsStore9[394] <= 19'd0;
		WeightsStore9[395] <= 19'd0;
		WeightsStore9[396] <= 19'd0;
		WeightsStore9[397] <= 19'd0;
		WeightsStore9[398] <= 19'd0;
		WeightsStore9[399] <= 19'd0;
		WeightsStore9[400] <= 19'd0;
		WeightsStore9[401] <= 19'd0;
		WeightsStore9[402] <= 19'd0;
		WeightsStore9[403] <= 19'd0;
		WeightsStore9[404] <= 19'd0;
		WeightsStore9[405] <= 19'd0;
		WeightsStore9[406] <= 19'd0;
		WeightsStore9[407] <= 19'd0;
		WeightsStore9[408] <= 19'd0;
		WeightsStore9[409] <= 19'd0;
		WeightsStore9[410] <= 19'd0;
		WeightsStore9[411] <= 19'd0;
		WeightsStore9[412] <= 19'd0;
		WeightsStore9[413] <= 19'd0;
		WeightsStore9[414] <= 19'd0;
		WeightsStore9[415] <= 19'd0;
		WeightsStore9[416] <= 19'd0;
		WeightsStore9[417] <= 19'd0;
		WeightsStore9[418] <= 19'd0;
		WeightsStore9[419] <= 19'd0;
		WeightsStore9[420] <= 19'd0;
		WeightsStore9[421] <= 19'd0;
		WeightsStore9[422] <= 19'd0;
		WeightsStore9[423] <= 19'd0;
		WeightsStore9[424] <= 19'd0;
		WeightsStore9[425] <= 19'd0;
		WeightsStore9[426] <= 19'd0;
		WeightsStore9[427] <= 19'd0;
		WeightsStore9[428] <= 19'd0;
		WeightsStore9[429] <= 19'd0;
		WeightsStore9[430] <= 19'd0;
		WeightsStore9[431] <= 19'd0;
		WeightsStore9[432] <= 19'd0;
		WeightsStore9[433] <= 19'd0;
		WeightsStore9[434] <= 19'd0;
		WeightsStore9[435] <= 19'd0;
		WeightsStore9[436] <= 19'd0;
		WeightsStore9[437] <= 19'd0;
		WeightsStore9[438] <= 19'd0;
		WeightsStore9[439] <= 19'd0;
		WeightsStore9[440] <= 19'd0;
		WeightsStore9[441] <= 19'd0;
		WeightsStore9[442] <= 19'd0;
		WeightsStore9[443] <= 19'd0;
		WeightsStore9[444] <= 19'd0;
		WeightsStore9[445] <= 19'd0;
		WeightsStore9[446] <= 19'd0;
		WeightsStore9[447] <= 19'd0;
		WeightsStore9[448] <= 19'd0;
		WeightsStore9[449] <= 19'd0;
		WeightsStore9[450] <= 19'd0;
		WeightsStore9[451] <= 19'd0;
		WeightsStore9[452] <= 19'd0;
		WeightsStore9[453] <= 19'd0;
		WeightsStore9[454] <= 19'd0;
		WeightsStore9[455] <= 19'd0;
		WeightsStore9[456] <= 19'd0;
		WeightsStore9[457] <= 19'd0;
		WeightsStore9[458] <= 19'd0;
		WeightsStore9[459] <= 19'd0;
		WeightsStore9[460] <= 19'd0;
		WeightsStore9[461] <= 19'd0;
		WeightsStore9[462] <= 19'd0;
		WeightsStore9[463] <= 19'd0;
		WeightsStore9[464] <= 19'd0;
		WeightsStore9[465] <= 19'd0;
		WeightsStore9[466] <= 19'd0;
		WeightsStore9[467] <= 19'd0;
		WeightsStore9[468] <= 19'd0;
		WeightsStore9[469] <= 19'd0;
		WeightsStore9[470] <= 19'd0;
		WeightsStore9[471] <= 19'd0;
		WeightsStore9[472] <= 19'd0;
		WeightsStore9[473] <= 19'd0;
		WeightsStore9[474] <= 19'd0;
		WeightsStore9[475] <= 19'd0;
		WeightsStore9[476] <= 19'd0;
		WeightsStore9[477] <= 19'd0;
		WeightsStore9[478] <= 19'd0;
		WeightsStore9[479] <= 19'd0;
		WeightsStore9[480] <= 19'd0;
		WeightsStore9[481] <= 19'd0;
		WeightsStore9[482] <= 19'd0;
		WeightsStore9[483] <= 19'd0;
		WeightsStore9[484] <= 19'd0;
		WeightsStore9[485] <= 19'd0;
		WeightsStore9[486] <= 19'd0;
		WeightsStore9[487] <= 19'd0;
		WeightsStore9[488] <= 19'd0;
		WeightsStore9[489] <= 19'd0;
		WeightsStore9[490] <= 19'd0;
		WeightsStore9[491] <= 19'd0;
		WeightsStore9[492] <= 19'd0;
		WeightsStore9[493] <= 19'd0;
		WeightsStore9[494] <= 19'd0;
		WeightsStore9[495] <= 19'd0;
		WeightsStore9[496] <= 19'd0;
		WeightsStore9[497] <= 19'd0;
		WeightsStore9[498] <= 19'd0;
		WeightsStore9[499] <= 19'd0;
		WeightsStore9[500] <= 19'd0;
		WeightsStore9[501] <= 19'd0;
		WeightsStore9[502] <= 19'd0;
		WeightsStore9[503] <= 19'd0;
		WeightsStore9[504] <= 19'd0;
		WeightsStore9[505] <= 19'd0;
		WeightsStore9[506] <= 19'd0;
		WeightsStore9[507] <= 19'd0;
		WeightsStore9[508] <= 19'd0;
		WeightsStore9[509] <= 19'd0;
		WeightsStore9[510] <= 19'd0;
		WeightsStore9[511] <= 19'd0;
		WeightsStore9[512] <= 19'd0;
		WeightsStore9[513] <= 19'd0;
		WeightsStore9[514] <= 19'd0;
		WeightsStore9[515] <= 19'd0;
		WeightsStore9[516] <= 19'd0;
		WeightsStore9[517] <= 19'd0;
		WeightsStore9[518] <= 19'd0;
		WeightsStore9[519] <= 19'd0;
		WeightsStore9[520] <= 19'd0;
		WeightsStore9[521] <= 19'd0;
		WeightsStore9[522] <= 19'd0;
		WeightsStore9[523] <= 19'd0;
		WeightsStore9[524] <= 19'd0;
		WeightsStore9[525] <= 19'd0;
		WeightsStore9[526] <= 19'd0;
		WeightsStore9[527] <= 19'd0;
		WeightsStore9[528] <= 19'd0;
		WeightsStore9[529] <= 19'd0;
		WeightsStore9[530] <= 19'd0;
		WeightsStore9[531] <= 19'd0;
		WeightsStore9[532] <= 19'd0;
		WeightsStore9[533] <= 19'd0;
		WeightsStore9[534] <= 19'd0;
		WeightsStore9[535] <= 19'd0;
		WeightsStore9[536] <= 19'd0;
		WeightsStore9[537] <= 19'd0;
		WeightsStore9[538] <= 19'd0;
		WeightsStore9[539] <= 19'd0;
		WeightsStore9[540] <= 19'd0;
		WeightsStore9[541] <= 19'd0;
		WeightsStore9[542] <= 19'd0;
		WeightsStore9[543] <= 19'd0;
		WeightsStore9[544] <= 19'd0;
		WeightsStore9[545] <= 19'd0;
		WeightsStore9[546] <= 19'd0;
		WeightsStore9[547] <= 19'd0;
		WeightsStore9[548] <= 19'd0;
		WeightsStore9[549] <= 19'd0;
		WeightsStore9[550] <= 19'd0;
		WeightsStore9[551] <= 19'd0;
		WeightsStore9[552] <= 19'd0;
		WeightsStore9[553] <= 19'd0;
		WeightsStore9[554] <= 19'd0;
		WeightsStore9[555] <= 19'd0;
		WeightsStore9[556] <= 19'd0;
		WeightsStore9[557] <= 19'd0;
		WeightsStore9[558] <= 19'd0;
		WeightsStore9[559] <= 19'd0;
		WeightsStore9[560] <= 19'd0;
		WeightsStore9[561] <= 19'd0;
		WeightsStore9[562] <= 19'd0;
		WeightsStore9[563] <= 19'd0;
		WeightsStore9[564] <= 19'd0;
		WeightsStore9[565] <= 19'd0;
		WeightsStore9[566] <= 19'd0;
		WeightsStore9[567] <= 19'd0;
		WeightsStore9[568] <= 19'd0;
		WeightsStore9[569] <= 19'd0;
		WeightsStore9[570] <= 19'd0;
		WeightsStore9[571] <= 19'd0;
		WeightsStore9[572] <= 19'd0;
		WeightsStore9[573] <= 19'd0;
		WeightsStore9[574] <= 19'd0;
		WeightsStore9[575] <= 19'd0;
		WeightsStore9[576] <= 19'd0;
		WeightsStore9[577] <= 19'd0;
		WeightsStore9[578] <= 19'd0;
		WeightsStore9[579] <= 19'd0;
		WeightsStore9[580] <= 19'd0;
		WeightsStore9[581] <= 19'd0;
		WeightsStore9[582] <= 19'd0;
		WeightsStore9[583] <= 19'd0;
		WeightsStore9[584] <= 19'd0;
		WeightsStore9[585] <= 19'd0;
		WeightsStore9[586] <= 19'd0;
		WeightsStore9[587] <= 19'd0;
		WeightsStore9[588] <= 19'd0;
		WeightsStore9[589] <= 19'd0;
		WeightsStore9[590] <= 19'd0;
		WeightsStore9[591] <= 19'd0;
		WeightsStore9[592] <= 19'd0;
		WeightsStore9[593] <= 19'd0;
		WeightsStore9[594] <= 19'd0;
		WeightsStore9[595] <= 19'd0;
		WeightsStore9[596] <= 19'd0;
		WeightsStore9[597] <= 19'd0;
		WeightsStore9[598] <= 19'd0;
		WeightsStore9[599] <= 19'd0;
		WeightsStore9[600] <= 19'd0;
		WeightsStore9[601] <= 19'd0;
		WeightsStore9[602] <= 19'd0;
		WeightsStore9[603] <= 19'd0;
		WeightsStore9[604] <= 19'd0;
		WeightsStore9[605] <= 19'd0;
		WeightsStore9[606] <= 19'd0;
		WeightsStore9[607] <= 19'd0;
		WeightsStore9[608] <= 19'd0;
		WeightsStore9[609] <= 19'd0;
		WeightsStore9[610] <= 19'd0;
		WeightsStore9[611] <= 19'd0;
		WeightsStore9[612] <= 19'd0;
		WeightsStore9[613] <= 19'd0;
		WeightsStore9[614] <= 19'd0;
		WeightsStore9[615] <= 19'd0;
		WeightsStore9[616] <= 19'd0;
		WeightsStore9[617] <= 19'd0;
		WeightsStore9[618] <= 19'd0;
		WeightsStore9[619] <= 19'd0;
		WeightsStore9[620] <= 19'd0;
		WeightsStore9[621] <= 19'd0;
		WeightsStore9[622] <= 19'd0;
		WeightsStore9[623] <= 19'd0;
		WeightsStore9[624] <= 19'd0;
		WeightsStore9[625] <= 19'd0;
		WeightsStore9[626] <= 19'd0;
		WeightsStore9[627] <= 19'd0;
		WeightsStore9[628] <= 19'd0;
		WeightsStore9[629] <= 19'd0;
		WeightsStore9[630] <= 19'd0;
		WeightsStore9[631] <= 19'd0;
		WeightsStore9[632] <= 19'd0;
		WeightsStore9[633] <= 19'd0;
		WeightsStore9[634] <= 19'd0;
		WeightsStore9[635] <= 19'd0;
		WeightsStore9[636] <= 19'd0;
		WeightsStore9[637] <= 19'd0;
		WeightsStore9[638] <= 19'd0;
		WeightsStore9[639] <= 19'd0;
		WeightsStore9[640] <= 19'd0;
		WeightsStore9[641] <= 19'd0;
		WeightsStore9[642] <= 19'd0;
		WeightsStore9[643] <= 19'd0;
		WeightsStore9[644] <= 19'd0;
		WeightsStore9[645] <= 19'd0;
		WeightsStore9[646] <= 19'd0;
		WeightsStore9[647] <= 19'd0;
		WeightsStore9[648] <= 19'd0;
		WeightsStore9[649] <= 19'd0;
		WeightsStore9[650] <= 19'd0;
		WeightsStore9[651] <= 19'd0;
		WeightsStore9[652] <= 19'd0;
		WeightsStore9[653] <= 19'd0;
		WeightsStore9[654] <= 19'd0;
		WeightsStore9[655] <= 19'd0;
		WeightsStore9[656] <= 19'd0;
		WeightsStore9[657] <= 19'd0;
		WeightsStore9[658] <= 19'd0;
		WeightsStore9[659] <= 19'd0;
		WeightsStore9[660] <= 19'd0;
		WeightsStore9[661] <= 19'd0;
		WeightsStore9[662] <= 19'd0;
		WeightsStore9[663] <= 19'd0;
		WeightsStore9[664] <= 19'd0;
		WeightsStore9[665] <= 19'd0;
		WeightsStore9[666] <= 19'd0;
		WeightsStore9[667] <= 19'd0;
		WeightsStore9[668] <= 19'd0;
		WeightsStore9[669] <= 19'd0;
		WeightsStore9[670] <= 19'd0;
		WeightsStore9[671] <= 19'd0;
		WeightsStore9[672] <= 19'd0;
		WeightsStore9[673] <= 19'd0;
		WeightsStore9[674] <= 19'd0;
		WeightsStore9[675] <= 19'd0;
		WeightsStore9[676] <= 19'd0;
		WeightsStore9[677] <= 19'd0;
		WeightsStore9[678] <= 19'd0;
		WeightsStore9[679] <= 19'd0;
		WeightsStore9[680] <= 19'd0;
		WeightsStore9[681] <= 19'd0;
		WeightsStore9[682] <= 19'd0;
		WeightsStore9[683] <= 19'd0;
		WeightsStore9[684] <= 19'd0;
		WeightsStore9[685] <= 19'd0;
		WeightsStore9[686] <= 19'd0;
		WeightsStore9[687] <= 19'd0;
		WeightsStore9[688] <= 19'd0;
		WeightsStore9[689] <= 19'd0;
		WeightsStore9[690] <= 19'd0;
		WeightsStore9[691] <= 19'd0;
		WeightsStore9[692] <= 19'd0;
		WeightsStore9[693] <= 19'd0;
		WeightsStore9[694] <= 19'd0;
		WeightsStore9[695] <= 19'd0;
		WeightsStore9[696] <= 19'd0;
		WeightsStore9[697] <= 19'd0;
		WeightsStore9[698] <= 19'd0;
		WeightsStore9[699] <= 19'd0;
		WeightsStore9[700] <= 19'd0;
		WeightsStore9[701] <= 19'd0;
		WeightsStore9[702] <= 19'd0;
		WeightsStore9[703] <= 19'd0;
		WeightsStore9[704] <= 19'd0;
		WeightsStore9[705] <= 19'd0;
		WeightsStore9[706] <= 19'd0;
		WeightsStore9[707] <= 19'd0;
		WeightsStore9[708] <= 19'd0;
		WeightsStore9[709] <= 19'd0;
		WeightsStore9[710] <= 19'd0;
		WeightsStore9[711] <= 19'd0;
		WeightsStore9[712] <= 19'd0;
		WeightsStore9[713] <= 19'd0;
		WeightsStore9[714] <= 19'd0;
		WeightsStore9[715] <= 19'd0;
		WeightsStore9[716] <= 19'd0;
		WeightsStore9[717] <= 19'd0;
		WeightsStore9[718] <= 19'd0;
		WeightsStore9[719] <= 19'd0;
		WeightsStore9[720] <= 19'd0;
		WeightsStore9[721] <= 19'd0;
		WeightsStore9[722] <= 19'd0;
		WeightsStore9[723] <= 19'd0;
		WeightsStore9[724] <= 19'd0;
		WeightsStore9[725] <= 19'd0;
		WeightsStore9[726] <= 19'd0;
		WeightsStore9[727] <= 19'd0;
		WeightsStore9[728] <= 19'd0;
		WeightsStore9[729] <= 19'd0;
		WeightsStore9[730] <= 19'd0;
		WeightsStore9[731] <= 19'd0;
		WeightsStore9[732] <= 19'd0;
		WeightsStore9[733] <= 19'd0;
		WeightsStore9[734] <= 19'd0;
		WeightsStore9[735] <= 19'd0;
		WeightsStore9[736] <= 19'd0;
		WeightsStore9[737] <= 19'd0;
		WeightsStore9[738] <= 19'd0;
		WeightsStore9[739] <= 19'd0;
		WeightsStore9[740] <= 19'd0;
		WeightsStore9[741] <= 19'd0;
		WeightsStore9[742] <= 19'd0;
		WeightsStore9[743] <= 19'd0;
		WeightsStore9[744] <= 19'd0;
		WeightsStore9[745] <= 19'd0;
		WeightsStore9[746] <= 19'd0;
		WeightsStore9[747] <= 19'd0;
		WeightsStore9[748] <= 19'd0;
		WeightsStore9[749] <= 19'd0;
		WeightsStore9[750] <= 19'd0;
		WeightsStore9[751] <= 19'd0;
		WeightsStore9[752] <= 19'd0;
		WeightsStore9[753] <= 19'd0;
		WeightsStore9[754] <= 19'd0;
		WeightsStore9[755] <= 19'd0;
		WeightsStore9[756] <= 19'd0;
		WeightsStore9[757] <= 19'd0;
		WeightsStore9[758] <= 19'd0;
		WeightsStore9[759] <= 19'd0;
		WeightsStore9[760] <= 19'd0;
		WeightsStore9[761] <= 19'd0;
		WeightsStore9[762] <= 19'd0;
		WeightsStore9[763] <= 19'd0;
		WeightsStore9[764] <= 19'd0;
		WeightsStore9[765] <= 19'd0;
		WeightsStore9[766] <= 19'd0;
		WeightsStore9[767] <= 19'd0;
		WeightsStore9[768] <= 19'd0;
		WeightsStore9[769] <= 19'd0;
		WeightsStore9[770] <= 19'd0;
		WeightsStore9[771] <= 19'd0;
		WeightsStore9[772] <= 19'd0;
		WeightsStore9[773] <= 19'd0;
		WeightsStore9[774] <= 19'd0;
		WeightsStore9[775] <= 19'd0;
		WeightsStore9[776] <= 19'd0;
		WeightsStore9[777] <= 19'd0;
		WeightsStore9[778] <= 19'd0;
		WeightsStore9[779] <= 19'd0;
		WeightsStore9[780] <= 19'd0;
		WeightsStore9[781] <= 19'd0;
		WeightsStore9[782] <= 19'd0;
		WeightsStore9[783] <= 19'd0;
		WeightsStore9[784] <= 19'd0;
	end
	if(Input_Valid == 1'b1)begin
		switchCounter <= 32'd0;
		ready <= 1'b0;
		internalReset = 1'b0;
		PixelsStore[0] <= Pix_0;
		PixelsStore[1] <= Pix_1;
		PixelsStore[2] <= Pix_2;
		PixelsStore[3] <= Pix_3;
		PixelsStore[4] <= Pix_4;
		PixelsStore[5] <= Pix_5;
		PixelsStore[6] <= Pix_6;
		PixelsStore[7] <= Pix_7;
		PixelsStore[8] <= Pix_8;
		PixelsStore[9] <= Pix_9;
		PixelsStore[10] <= Pix_10;
		PixelsStore[11] <= Pix_11;
		PixelsStore[12] <= Pix_12;
		PixelsStore[13] <= Pix_13;
		PixelsStore[14] <= Pix_14;
		PixelsStore[15] <= Pix_15;
		PixelsStore[16] <= Pix_16;
		PixelsStore[17] <= Pix_17;
		PixelsStore[18] <= Pix_18;
		PixelsStore[19] <= Pix_19;
		PixelsStore[20] <= Pix_20;
		PixelsStore[21] <= Pix_21;
		PixelsStore[22] <= Pix_22;
		PixelsStore[23] <= Pix_23;
		PixelsStore[24] <= Pix_24;
		PixelsStore[25] <= Pix_25;
		PixelsStore[26] <= Pix_26;
		PixelsStore[27] <= Pix_27;
		PixelsStore[28] <= Pix_28;
		PixelsStore[29] <= Pix_29;
		PixelsStore[30] <= Pix_30;
		PixelsStore[31] <= Pix_31;
		PixelsStore[32] <= Pix_32;
		PixelsStore[33] <= Pix_33;
		PixelsStore[34] <= Pix_34;
		PixelsStore[35] <= Pix_35;
		PixelsStore[36] <= Pix_36;
		PixelsStore[37] <= Pix_37;
		PixelsStore[38] <= Pix_38;
		PixelsStore[39] <= Pix_39;
		PixelsStore[40] <= Pix_40;
		PixelsStore[41] <= Pix_41;
		PixelsStore[42] <= Pix_42;
		PixelsStore[43] <= Pix_43;
		PixelsStore[44] <= Pix_44;
		PixelsStore[45] <= Pix_45;
		PixelsStore[46] <= Pix_46;
		PixelsStore[47] <= Pix_47;
		PixelsStore[48] <= Pix_48;
		PixelsStore[49] <= Pix_49;
		PixelsStore[50] <= Pix_50;
		PixelsStore[51] <= Pix_51;
		PixelsStore[52] <= Pix_52;
		PixelsStore[53] <= Pix_53;
		PixelsStore[54] <= Pix_54;
		PixelsStore[55] <= Pix_55;
		PixelsStore[56] <= Pix_56;
		PixelsStore[57] <= Pix_57;
		PixelsStore[58] <= Pix_58;
		PixelsStore[59] <= Pix_59;
		PixelsStore[60] <= Pix_60;
		PixelsStore[61] <= Pix_61;
		PixelsStore[62] <= Pix_62;
		PixelsStore[63] <= Pix_63;
		PixelsStore[64] <= Pix_64;
		PixelsStore[65] <= Pix_65;
		PixelsStore[66] <= Pix_66;
		PixelsStore[67] <= Pix_67;
		PixelsStore[68] <= Pix_68;
		PixelsStore[69] <= Pix_69;
		PixelsStore[70] <= Pix_70;
		PixelsStore[71] <= Pix_71;
		PixelsStore[72] <= Pix_72;
		PixelsStore[73] <= Pix_73;
		PixelsStore[74] <= Pix_74;
		PixelsStore[75] <= Pix_75;
		PixelsStore[76] <= Pix_76;
		PixelsStore[77] <= Pix_77;
		PixelsStore[78] <= Pix_78;
		PixelsStore[79] <= Pix_79;
		PixelsStore[80] <= Pix_80;
		PixelsStore[81] <= Pix_81;
		PixelsStore[82] <= Pix_82;
		PixelsStore[83] <= Pix_83;
		PixelsStore[84] <= Pix_84;
		PixelsStore[85] <= Pix_85;
		PixelsStore[86] <= Pix_86;
		PixelsStore[87] <= Pix_87;
		PixelsStore[88] <= Pix_88;
		PixelsStore[89] <= Pix_89;
		PixelsStore[90] <= Pix_90;
		PixelsStore[91] <= Pix_91;
		PixelsStore[92] <= Pix_92;
		PixelsStore[93] <= Pix_93;
		PixelsStore[94] <= Pix_94;
		PixelsStore[95] <= Pix_95;
		PixelsStore[96] <= Pix_96;
		PixelsStore[97] <= Pix_97;
		PixelsStore[98] <= Pix_98;
		PixelsStore[99] <= Pix_99;
		PixelsStore[100] <= Pix_100;
		PixelsStore[101] <= Pix_101;
		PixelsStore[102] <= Pix_102;
		PixelsStore[103] <= Pix_103;
		PixelsStore[104] <= Pix_104;
		PixelsStore[105] <= Pix_105;
		PixelsStore[106] <= Pix_106;
		PixelsStore[107] <= Pix_107;
		PixelsStore[108] <= Pix_108;
		PixelsStore[109] <= Pix_109;
		PixelsStore[110] <= Pix_110;
		PixelsStore[111] <= Pix_111;
		PixelsStore[112] <= Pix_112;
		PixelsStore[113] <= Pix_113;
		PixelsStore[114] <= Pix_114;
		PixelsStore[115] <= Pix_115;
		PixelsStore[116] <= Pix_116;
		PixelsStore[117] <= Pix_117;
		PixelsStore[118] <= Pix_118;
		PixelsStore[119] <= Pix_119;
		PixelsStore[120] <= Pix_120;
		PixelsStore[121] <= Pix_121;
		PixelsStore[122] <= Pix_122;
		PixelsStore[123] <= Pix_123;
		PixelsStore[124] <= Pix_124;
		PixelsStore[125] <= Pix_125;
		PixelsStore[126] <= Pix_126;
		PixelsStore[127] <= Pix_127;
		PixelsStore[128] <= Pix_128;
		PixelsStore[129] <= Pix_129;
		PixelsStore[130] <= Pix_130;
		PixelsStore[131] <= Pix_131;
		PixelsStore[132] <= Pix_132;
		PixelsStore[133] <= Pix_133;
		PixelsStore[134] <= Pix_134;
		PixelsStore[135] <= Pix_135;
		PixelsStore[136] <= Pix_136;
		PixelsStore[137] <= Pix_137;
		PixelsStore[138] <= Pix_138;
		PixelsStore[139] <= Pix_139;
		PixelsStore[140] <= Pix_140;
		PixelsStore[141] <= Pix_141;
		PixelsStore[142] <= Pix_142;
		PixelsStore[143] <= Pix_143;
		PixelsStore[144] <= Pix_144;
		PixelsStore[145] <= Pix_145;
		PixelsStore[146] <= Pix_146;
		PixelsStore[147] <= Pix_147;
		PixelsStore[148] <= Pix_148;
		PixelsStore[149] <= Pix_149;
		PixelsStore[150] <= Pix_150;
		PixelsStore[151] <= Pix_151;
		PixelsStore[152] <= Pix_152;
		PixelsStore[153] <= Pix_153;
		PixelsStore[154] <= Pix_154;
		PixelsStore[155] <= Pix_155;
		PixelsStore[156] <= Pix_156;
		PixelsStore[157] <= Pix_157;
		PixelsStore[158] <= Pix_158;
		PixelsStore[159] <= Pix_159;
		PixelsStore[160] <= Pix_160;
		PixelsStore[161] <= Pix_161;
		PixelsStore[162] <= Pix_162;
		PixelsStore[163] <= Pix_163;
		PixelsStore[164] <= Pix_164;
		PixelsStore[165] <= Pix_165;
		PixelsStore[166] <= Pix_166;
		PixelsStore[167] <= Pix_167;
		PixelsStore[168] <= Pix_168;
		PixelsStore[169] <= Pix_169;
		PixelsStore[170] <= Pix_170;
		PixelsStore[171] <= Pix_171;
		PixelsStore[172] <= Pix_172;
		PixelsStore[173] <= Pix_173;
		PixelsStore[174] <= Pix_174;
		PixelsStore[175] <= Pix_175;
		PixelsStore[176] <= Pix_176;
		PixelsStore[177] <= Pix_177;
		PixelsStore[178] <= Pix_178;
		PixelsStore[179] <= Pix_179;
		PixelsStore[180] <= Pix_180;
		PixelsStore[181] <= Pix_181;
		PixelsStore[182] <= Pix_182;
		PixelsStore[183] <= Pix_183;
		PixelsStore[184] <= Pix_184;
		PixelsStore[185] <= Pix_185;
		PixelsStore[186] <= Pix_186;
		PixelsStore[187] <= Pix_187;
		PixelsStore[188] <= Pix_188;
		PixelsStore[189] <= Pix_189;
		PixelsStore[190] <= Pix_190;
		PixelsStore[191] <= Pix_191;
		PixelsStore[192] <= Pix_192;
		PixelsStore[193] <= Pix_193;
		PixelsStore[194] <= Pix_194;
		PixelsStore[195] <= Pix_195;
		PixelsStore[196] <= Pix_196;
		PixelsStore[197] <= Pix_197;
		PixelsStore[198] <= Pix_198;
		PixelsStore[199] <= Pix_199;
		PixelsStore[200] <= Pix_200;
		PixelsStore[201] <= Pix_201;
		PixelsStore[202] <= Pix_202;
		PixelsStore[203] <= Pix_203;
		PixelsStore[204] <= Pix_204;
		PixelsStore[205] <= Pix_205;
		PixelsStore[206] <= Pix_206;
		PixelsStore[207] <= Pix_207;
		PixelsStore[208] <= Pix_208;
		PixelsStore[209] <= Pix_209;
		PixelsStore[210] <= Pix_210;
		PixelsStore[211] <= Pix_211;
		PixelsStore[212] <= Pix_212;
		PixelsStore[213] <= Pix_213;
		PixelsStore[214] <= Pix_214;
		PixelsStore[215] <= Pix_215;
		PixelsStore[216] <= Pix_216;
		PixelsStore[217] <= Pix_217;
		PixelsStore[218] <= Pix_218;
		PixelsStore[219] <= Pix_219;
		PixelsStore[220] <= Pix_220;
		PixelsStore[221] <= Pix_221;
		PixelsStore[222] <= Pix_222;
		PixelsStore[223] <= Pix_223;
		PixelsStore[224] <= Pix_224;
		PixelsStore[225] <= Pix_225;
		PixelsStore[226] <= Pix_226;
		PixelsStore[227] <= Pix_227;
		PixelsStore[228] <= Pix_228;
		PixelsStore[229] <= Pix_229;
		PixelsStore[230] <= Pix_230;
		PixelsStore[231] <= Pix_231;
		PixelsStore[232] <= Pix_232;
		PixelsStore[233] <= Pix_233;
		PixelsStore[234] <= Pix_234;
		PixelsStore[235] <= Pix_235;
		PixelsStore[236] <= Pix_236;
		PixelsStore[237] <= Pix_237;
		PixelsStore[238] <= Pix_238;
		PixelsStore[239] <= Pix_239;
		PixelsStore[240] <= Pix_240;
		PixelsStore[241] <= Pix_241;
		PixelsStore[242] <= Pix_242;
		PixelsStore[243] <= Pix_243;
		PixelsStore[244] <= Pix_244;
		PixelsStore[245] <= Pix_245;
		PixelsStore[246] <= Pix_246;
		PixelsStore[247] <= Pix_247;
		PixelsStore[248] <= Pix_248;
		PixelsStore[249] <= Pix_249;
		PixelsStore[250] <= Pix_250;
		PixelsStore[251] <= Pix_251;
		PixelsStore[252] <= Pix_252;
		PixelsStore[253] <= Pix_253;
		PixelsStore[254] <= Pix_254;
		PixelsStore[255] <= Pix_255;
		PixelsStore[256] <= Pix_256;
		PixelsStore[257] <= Pix_257;
		PixelsStore[258] <= Pix_258;
		PixelsStore[259] <= Pix_259;
		PixelsStore[260] <= Pix_260;
		PixelsStore[261] <= Pix_261;
		PixelsStore[262] <= Pix_262;
		PixelsStore[263] <= Pix_263;
		PixelsStore[264] <= Pix_264;
		PixelsStore[265] <= Pix_265;
		PixelsStore[266] <= Pix_266;
		PixelsStore[267] <= Pix_267;
		PixelsStore[268] <= Pix_268;
		PixelsStore[269] <= Pix_269;
		PixelsStore[270] <= Pix_270;
		PixelsStore[271] <= Pix_271;
		PixelsStore[272] <= Pix_272;
		PixelsStore[273] <= Pix_273;
		PixelsStore[274] <= Pix_274;
		PixelsStore[275] <= Pix_275;
		PixelsStore[276] <= Pix_276;
		PixelsStore[277] <= Pix_277;
		PixelsStore[278] <= Pix_278;
		PixelsStore[279] <= Pix_279;
		PixelsStore[280] <= Pix_280;
		PixelsStore[281] <= Pix_281;
		PixelsStore[282] <= Pix_282;
		PixelsStore[283] <= Pix_283;
		PixelsStore[284] <= Pix_284;
		PixelsStore[285] <= Pix_285;
		PixelsStore[286] <= Pix_286;
		PixelsStore[287] <= Pix_287;
		PixelsStore[288] <= Pix_288;
		PixelsStore[289] <= Pix_289;
		PixelsStore[290] <= Pix_290;
		PixelsStore[291] <= Pix_291;
		PixelsStore[292] <= Pix_292;
		PixelsStore[293] <= Pix_293;
		PixelsStore[294] <= Pix_294;
		PixelsStore[295] <= Pix_295;
		PixelsStore[296] <= Pix_296;
		PixelsStore[297] <= Pix_297;
		PixelsStore[298] <= Pix_298;
		PixelsStore[299] <= Pix_299;
		PixelsStore[300] <= Pix_300;
		PixelsStore[301] <= Pix_301;
		PixelsStore[302] <= Pix_302;
		PixelsStore[303] <= Pix_303;
		PixelsStore[304] <= Pix_304;
		PixelsStore[305] <= Pix_305;
		PixelsStore[306] <= Pix_306;
		PixelsStore[307] <= Pix_307;
		PixelsStore[308] <= Pix_308;
		PixelsStore[309] <= Pix_309;
		PixelsStore[310] <= Pix_310;
		PixelsStore[311] <= Pix_311;
		PixelsStore[312] <= Pix_312;
		PixelsStore[313] <= Pix_313;
		PixelsStore[314] <= Pix_314;
		PixelsStore[315] <= Pix_315;
		PixelsStore[316] <= Pix_316;
		PixelsStore[317] <= Pix_317;
		PixelsStore[318] <= Pix_318;
		PixelsStore[319] <= Pix_319;
		PixelsStore[320] <= Pix_320;
		PixelsStore[321] <= Pix_321;
		PixelsStore[322] <= Pix_322;
		PixelsStore[323] <= Pix_323;
		PixelsStore[324] <= Pix_324;
		PixelsStore[325] <= Pix_325;
		PixelsStore[326] <= Pix_326;
		PixelsStore[327] <= Pix_327;
		PixelsStore[328] <= Pix_328;
		PixelsStore[329] <= Pix_329;
		PixelsStore[330] <= Pix_330;
		PixelsStore[331] <= Pix_331;
		PixelsStore[332] <= Pix_332;
		PixelsStore[333] <= Pix_333;
		PixelsStore[334] <= Pix_334;
		PixelsStore[335] <= Pix_335;
		PixelsStore[336] <= Pix_336;
		PixelsStore[337] <= Pix_337;
		PixelsStore[338] <= Pix_338;
		PixelsStore[339] <= Pix_339;
		PixelsStore[340] <= Pix_340;
		PixelsStore[341] <= Pix_341;
		PixelsStore[342] <= Pix_342;
		PixelsStore[343] <= Pix_343;
		PixelsStore[344] <= Pix_344;
		PixelsStore[345] <= Pix_345;
		PixelsStore[346] <= Pix_346;
		PixelsStore[347] <= Pix_347;
		PixelsStore[348] <= Pix_348;
		PixelsStore[349] <= Pix_349;
		PixelsStore[350] <= Pix_350;
		PixelsStore[351] <= Pix_351;
		PixelsStore[352] <= Pix_352;
		PixelsStore[353] <= Pix_353;
		PixelsStore[354] <= Pix_354;
		PixelsStore[355] <= Pix_355;
		PixelsStore[356] <= Pix_356;
		PixelsStore[357] <= Pix_357;
		PixelsStore[358] <= Pix_358;
		PixelsStore[359] <= Pix_359;
		PixelsStore[360] <= Pix_360;
		PixelsStore[361] <= Pix_361;
		PixelsStore[362] <= Pix_362;
		PixelsStore[363] <= Pix_363;
		PixelsStore[364] <= Pix_364;
		PixelsStore[365] <= Pix_365;
		PixelsStore[366] <= Pix_366;
		PixelsStore[367] <= Pix_367;
		PixelsStore[368] <= Pix_368;
		PixelsStore[369] <= Pix_369;
		PixelsStore[370] <= Pix_370;
		PixelsStore[371] <= Pix_371;
		PixelsStore[372] <= Pix_372;
		PixelsStore[373] <= Pix_373;
		PixelsStore[374] <= Pix_374;
		PixelsStore[375] <= Pix_375;
		PixelsStore[376] <= Pix_376;
		PixelsStore[377] <= Pix_377;
		PixelsStore[378] <= Pix_378;
		PixelsStore[379] <= Pix_379;
		PixelsStore[380] <= Pix_380;
		PixelsStore[381] <= Pix_381;
		PixelsStore[382] <= Pix_382;
		PixelsStore[383] <= Pix_383;
		PixelsStore[384] <= Pix_384;
		PixelsStore[385] <= Pix_385;
		PixelsStore[386] <= Pix_386;
		PixelsStore[387] <= Pix_387;
		PixelsStore[388] <= Pix_388;
		PixelsStore[389] <= Pix_389;
		PixelsStore[390] <= Pix_390;
		PixelsStore[391] <= Pix_391;
		PixelsStore[392] <= Pix_392;
		PixelsStore[393] <= Pix_393;
		PixelsStore[394] <= Pix_394;
		PixelsStore[395] <= Pix_395;
		PixelsStore[396] <= Pix_396;
		PixelsStore[397] <= Pix_397;
		PixelsStore[398] <= Pix_398;
		PixelsStore[399] <= Pix_399;
		PixelsStore[400] <= Pix_400;
		PixelsStore[401] <= Pix_401;
		PixelsStore[402] <= Pix_402;
		PixelsStore[403] <= Pix_403;
		PixelsStore[404] <= Pix_404;
		PixelsStore[405] <= Pix_405;
		PixelsStore[406] <= Pix_406;
		PixelsStore[407] <= Pix_407;
		PixelsStore[408] <= Pix_408;
		PixelsStore[409] <= Pix_409;
		PixelsStore[410] <= Pix_410;
		PixelsStore[411] <= Pix_411;
		PixelsStore[412] <= Pix_412;
		PixelsStore[413] <= Pix_413;
		PixelsStore[414] <= Pix_414;
		PixelsStore[415] <= Pix_415;
		PixelsStore[416] <= Pix_416;
		PixelsStore[417] <= Pix_417;
		PixelsStore[418] <= Pix_418;
		PixelsStore[419] <= Pix_419;
		PixelsStore[420] <= Pix_420;
		PixelsStore[421] <= Pix_421;
		PixelsStore[422] <= Pix_422;
		PixelsStore[423] <= Pix_423;
		PixelsStore[424] <= Pix_424;
		PixelsStore[425] <= Pix_425;
		PixelsStore[426] <= Pix_426;
		PixelsStore[427] <= Pix_427;
		PixelsStore[428] <= Pix_428;
		PixelsStore[429] <= Pix_429;
		PixelsStore[430] <= Pix_430;
		PixelsStore[431] <= Pix_431;
		PixelsStore[432] <= Pix_432;
		PixelsStore[433] <= Pix_433;
		PixelsStore[434] <= Pix_434;
		PixelsStore[435] <= Pix_435;
		PixelsStore[436] <= Pix_436;
		PixelsStore[437] <= Pix_437;
		PixelsStore[438] <= Pix_438;
		PixelsStore[439] <= Pix_439;
		PixelsStore[440] <= Pix_440;
		PixelsStore[441] <= Pix_441;
		PixelsStore[442] <= Pix_442;
		PixelsStore[443] <= Pix_443;
		PixelsStore[444] <= Pix_444;
		PixelsStore[445] <= Pix_445;
		PixelsStore[446] <= Pix_446;
		PixelsStore[447] <= Pix_447;
		PixelsStore[448] <= Pix_448;
		PixelsStore[449] <= Pix_449;
		PixelsStore[450] <= Pix_450;
		PixelsStore[451] <= Pix_451;
		PixelsStore[452] <= Pix_452;
		PixelsStore[453] <= Pix_453;
		PixelsStore[454] <= Pix_454;
		PixelsStore[455] <= Pix_455;
		PixelsStore[456] <= Pix_456;
		PixelsStore[457] <= Pix_457;
		PixelsStore[458] <= Pix_458;
		PixelsStore[459] <= Pix_459;
		PixelsStore[460] <= Pix_460;
		PixelsStore[461] <= Pix_461;
		PixelsStore[462] <= Pix_462;
		PixelsStore[463] <= Pix_463;
		PixelsStore[464] <= Pix_464;
		PixelsStore[465] <= Pix_465;
		PixelsStore[466] <= Pix_466;
		PixelsStore[467] <= Pix_467;
		PixelsStore[468] <= Pix_468;
		PixelsStore[469] <= Pix_469;
		PixelsStore[470] <= Pix_470;
		PixelsStore[471] <= Pix_471;
		PixelsStore[472] <= Pix_472;
		PixelsStore[473] <= Pix_473;
		PixelsStore[474] <= Pix_474;
		PixelsStore[475] <= Pix_475;
		PixelsStore[476] <= Pix_476;
		PixelsStore[477] <= Pix_477;
		PixelsStore[478] <= Pix_478;
		PixelsStore[479] <= Pix_479;
		PixelsStore[480] <= Pix_480;
		PixelsStore[481] <= Pix_481;
		PixelsStore[482] <= Pix_482;
		PixelsStore[483] <= Pix_483;
		PixelsStore[484] <= Pix_484;
		PixelsStore[485] <= Pix_485;
		PixelsStore[486] <= Pix_486;
		PixelsStore[487] <= Pix_487;
		PixelsStore[488] <= Pix_488;
		PixelsStore[489] <= Pix_489;
		PixelsStore[490] <= Pix_490;
		PixelsStore[491] <= Pix_491;
		PixelsStore[492] <= Pix_492;
		PixelsStore[493] <= Pix_493;
		PixelsStore[494] <= Pix_494;
		PixelsStore[495] <= Pix_495;
		PixelsStore[496] <= Pix_496;
		PixelsStore[497] <= Pix_497;
		PixelsStore[498] <= Pix_498;
		PixelsStore[499] <= Pix_499;
		PixelsStore[500] <= Pix_500;
		PixelsStore[501] <= Pix_501;
		PixelsStore[502] <= Pix_502;
		PixelsStore[503] <= Pix_503;
		PixelsStore[504] <= Pix_504;
		PixelsStore[505] <= Pix_505;
		PixelsStore[506] <= Pix_506;
		PixelsStore[507] <= Pix_507;
		PixelsStore[508] <= Pix_508;
		PixelsStore[509] <= Pix_509;
		PixelsStore[510] <= Pix_510;
		PixelsStore[511] <= Pix_511;
		PixelsStore[512] <= Pix_512;
		PixelsStore[513] <= Pix_513;
		PixelsStore[514] <= Pix_514;
		PixelsStore[515] <= Pix_515;
		PixelsStore[516] <= Pix_516;
		PixelsStore[517] <= Pix_517;
		PixelsStore[518] <= Pix_518;
		PixelsStore[519] <= Pix_519;
		PixelsStore[520] <= Pix_520;
		PixelsStore[521] <= Pix_521;
		PixelsStore[522] <= Pix_522;
		PixelsStore[523] <= Pix_523;
		PixelsStore[524] <= Pix_524;
		PixelsStore[525] <= Pix_525;
		PixelsStore[526] <= Pix_526;
		PixelsStore[527] <= Pix_527;
		PixelsStore[528] <= Pix_528;
		PixelsStore[529] <= Pix_529;
		PixelsStore[530] <= Pix_530;
		PixelsStore[531] <= Pix_531;
		PixelsStore[532] <= Pix_532;
		PixelsStore[533] <= Pix_533;
		PixelsStore[534] <= Pix_534;
		PixelsStore[535] <= Pix_535;
		PixelsStore[536] <= Pix_536;
		PixelsStore[537] <= Pix_537;
		PixelsStore[538] <= Pix_538;
		PixelsStore[539] <= Pix_539;
		PixelsStore[540] <= Pix_540;
		PixelsStore[541] <= Pix_541;
		PixelsStore[542] <= Pix_542;
		PixelsStore[543] <= Pix_543;
		PixelsStore[544] <= Pix_544;
		PixelsStore[545] <= Pix_545;
		PixelsStore[546] <= Pix_546;
		PixelsStore[547] <= Pix_547;
		PixelsStore[548] <= Pix_548;
		PixelsStore[549] <= Pix_549;
		PixelsStore[550] <= Pix_550;
		PixelsStore[551] <= Pix_551;
		PixelsStore[552] <= Pix_552;
		PixelsStore[553] <= Pix_553;
		PixelsStore[554] <= Pix_554;
		PixelsStore[555] <= Pix_555;
		PixelsStore[556] <= Pix_556;
		PixelsStore[557] <= Pix_557;
		PixelsStore[558] <= Pix_558;
		PixelsStore[559] <= Pix_559;
		PixelsStore[560] <= Pix_560;
		PixelsStore[561] <= Pix_561;
		PixelsStore[562] <= Pix_562;
		PixelsStore[563] <= Pix_563;
		PixelsStore[564] <= Pix_564;
		PixelsStore[565] <= Pix_565;
		PixelsStore[566] <= Pix_566;
		PixelsStore[567] <= Pix_567;
		PixelsStore[568] <= Pix_568;
		PixelsStore[569] <= Pix_569;
		PixelsStore[570] <= Pix_570;
		PixelsStore[571] <= Pix_571;
		PixelsStore[572] <= Pix_572;
		PixelsStore[573] <= Pix_573;
		PixelsStore[574] <= Pix_574;
		PixelsStore[575] <= Pix_575;
		PixelsStore[576] <= Pix_576;
		PixelsStore[577] <= Pix_577;
		PixelsStore[578] <= Pix_578;
		PixelsStore[579] <= Pix_579;
		PixelsStore[580] <= Pix_580;
		PixelsStore[581] <= Pix_581;
		PixelsStore[582] <= Pix_582;
		PixelsStore[583] <= Pix_583;
		PixelsStore[584] <= Pix_584;
		PixelsStore[585] <= Pix_585;
		PixelsStore[586] <= Pix_586;
		PixelsStore[587] <= Pix_587;
		PixelsStore[588] <= Pix_588;
		PixelsStore[589] <= Pix_589;
		PixelsStore[590] <= Pix_590;
		PixelsStore[591] <= Pix_591;
		PixelsStore[592] <= Pix_592;
		PixelsStore[593] <= Pix_593;
		PixelsStore[594] <= Pix_594;
		PixelsStore[595] <= Pix_595;
		PixelsStore[596] <= Pix_596;
		PixelsStore[597] <= Pix_597;
		PixelsStore[598] <= Pix_598;
		PixelsStore[599] <= Pix_599;
		PixelsStore[600] <= Pix_600;
		PixelsStore[601] <= Pix_601;
		PixelsStore[602] <= Pix_602;
		PixelsStore[603] <= Pix_603;
		PixelsStore[604] <= Pix_604;
		PixelsStore[605] <= Pix_605;
		PixelsStore[606] <= Pix_606;
		PixelsStore[607] <= Pix_607;
		PixelsStore[608] <= Pix_608;
		PixelsStore[609] <= Pix_609;
		PixelsStore[610] <= Pix_610;
		PixelsStore[611] <= Pix_611;
		PixelsStore[612] <= Pix_612;
		PixelsStore[613] <= Pix_613;
		PixelsStore[614] <= Pix_614;
		PixelsStore[615] <= Pix_615;
		PixelsStore[616] <= Pix_616;
		PixelsStore[617] <= Pix_617;
		PixelsStore[618] <= Pix_618;
		PixelsStore[619] <= Pix_619;
		PixelsStore[620] <= Pix_620;
		PixelsStore[621] <= Pix_621;
		PixelsStore[622] <= Pix_622;
		PixelsStore[623] <= Pix_623;
		PixelsStore[624] <= Pix_624;
		PixelsStore[625] <= Pix_625;
		PixelsStore[626] <= Pix_626;
		PixelsStore[627] <= Pix_627;
		PixelsStore[628] <= Pix_628;
		PixelsStore[629] <= Pix_629;
		PixelsStore[630] <= Pix_630;
		PixelsStore[631] <= Pix_631;
		PixelsStore[632] <= Pix_632;
		PixelsStore[633] <= Pix_633;
		PixelsStore[634] <= Pix_634;
		PixelsStore[635] <= Pix_635;
		PixelsStore[636] <= Pix_636;
		PixelsStore[637] <= Pix_637;
		PixelsStore[638] <= Pix_638;
		PixelsStore[639] <= Pix_639;
		PixelsStore[640] <= Pix_640;
		PixelsStore[641] <= Pix_641;
		PixelsStore[642] <= Pix_642;
		PixelsStore[643] <= Pix_643;
		PixelsStore[644] <= Pix_644;
		PixelsStore[645] <= Pix_645;
		PixelsStore[646] <= Pix_646;
		PixelsStore[647] <= Pix_647;
		PixelsStore[648] <= Pix_648;
		PixelsStore[649] <= Pix_649;
		PixelsStore[650] <= Pix_650;
		PixelsStore[651] <= Pix_651;
		PixelsStore[652] <= Pix_652;
		PixelsStore[653] <= Pix_653;
		PixelsStore[654] <= Pix_654;
		PixelsStore[655] <= Pix_655;
		PixelsStore[656] <= Pix_656;
		PixelsStore[657] <= Pix_657;
		PixelsStore[658] <= Pix_658;
		PixelsStore[659] <= Pix_659;
		PixelsStore[660] <= Pix_660;
		PixelsStore[661] <= Pix_661;
		PixelsStore[662] <= Pix_662;
		PixelsStore[663] <= Pix_663;
		PixelsStore[664] <= Pix_664;
		PixelsStore[665] <= Pix_665;
		PixelsStore[666] <= Pix_666;
		PixelsStore[667] <= Pix_667;
		PixelsStore[668] <= Pix_668;
		PixelsStore[669] <= Pix_669;
		PixelsStore[670] <= Pix_670;
		PixelsStore[671] <= Pix_671;
		PixelsStore[672] <= Pix_672;
		PixelsStore[673] <= Pix_673;
		PixelsStore[674] <= Pix_674;
		PixelsStore[675] <= Pix_675;
		PixelsStore[676] <= Pix_676;
		PixelsStore[677] <= Pix_677;
		PixelsStore[678] <= Pix_678;
		PixelsStore[679] <= Pix_679;
		PixelsStore[680] <= Pix_680;
		PixelsStore[681] <= Pix_681;
		PixelsStore[682] <= Pix_682;
		PixelsStore[683] <= Pix_683;
		PixelsStore[684] <= Pix_684;
		PixelsStore[685] <= Pix_685;
		PixelsStore[686] <= Pix_686;
		PixelsStore[687] <= Pix_687;
		PixelsStore[688] <= Pix_688;
		PixelsStore[689] <= Pix_689;
		PixelsStore[690] <= Pix_690;
		PixelsStore[691] <= Pix_691;
		PixelsStore[692] <= Pix_692;
		PixelsStore[693] <= Pix_693;
		PixelsStore[694] <= Pix_694;
		PixelsStore[695] <= Pix_695;
		PixelsStore[696] <= Pix_696;
		PixelsStore[697] <= Pix_697;
		PixelsStore[698] <= Pix_698;
		PixelsStore[699] <= Pix_699;
		PixelsStore[700] <= Pix_700;
		PixelsStore[701] <= Pix_701;
		PixelsStore[702] <= Pix_702;
		PixelsStore[703] <= Pix_703;
		PixelsStore[704] <= Pix_704;
		PixelsStore[705] <= Pix_705;
		PixelsStore[706] <= Pix_706;
		PixelsStore[707] <= Pix_707;
		PixelsStore[708] <= Pix_708;
		PixelsStore[709] <= Pix_709;
		PixelsStore[710] <= Pix_710;
		PixelsStore[711] <= Pix_711;
		PixelsStore[712] <= Pix_712;
		PixelsStore[713] <= Pix_713;
		PixelsStore[714] <= Pix_714;
		PixelsStore[715] <= Pix_715;
		PixelsStore[716] <= Pix_716;
		PixelsStore[717] <= Pix_717;
		PixelsStore[718] <= Pix_718;
		PixelsStore[719] <= Pix_719;
		PixelsStore[720] <= Pix_720;
		PixelsStore[721] <= Pix_721;
		PixelsStore[722] <= Pix_722;
		PixelsStore[723] <= Pix_723;
		PixelsStore[724] <= Pix_724;
		PixelsStore[725] <= Pix_725;
		PixelsStore[726] <= Pix_726;
		PixelsStore[727] <= Pix_727;
		PixelsStore[728] <= Pix_728;
		PixelsStore[729] <= Pix_729;
		PixelsStore[730] <= Pix_730;
		PixelsStore[731] <= Pix_731;
		PixelsStore[732] <= Pix_732;
		PixelsStore[733] <= Pix_733;
		PixelsStore[734] <= Pix_734;
		PixelsStore[735] <= Pix_735;
		PixelsStore[736] <= Pix_736;
		PixelsStore[737] <= Pix_737;
		PixelsStore[738] <= Pix_738;
		PixelsStore[739] <= Pix_739;
		PixelsStore[740] <= Pix_740;
		PixelsStore[741] <= Pix_741;
		PixelsStore[742] <= Pix_742;
		PixelsStore[743] <= Pix_743;
		PixelsStore[744] <= Pix_744;
		PixelsStore[745] <= Pix_745;
		PixelsStore[746] <= Pix_746;
		PixelsStore[747] <= Pix_747;
		PixelsStore[748] <= Pix_748;
		PixelsStore[749] <= Pix_749;
		PixelsStore[750] <= Pix_750;
		PixelsStore[751] <= Pix_751;
		PixelsStore[752] <= Pix_752;
		PixelsStore[753] <= Pix_753;
		PixelsStore[754] <= Pix_754;
		PixelsStore[755] <= Pix_755;
		PixelsStore[756] <= Pix_756;
		PixelsStore[757] <= Pix_757;
		PixelsStore[758] <= Pix_758;
		PixelsStore[759] <= Pix_759;
		PixelsStore[760] <= Pix_760;
		PixelsStore[761] <= Pix_761;
		PixelsStore[762] <= Pix_762;
		PixelsStore[763] <= Pix_763;
		PixelsStore[764] <= Pix_764;
		PixelsStore[765] <= Pix_765;
		PixelsStore[766] <= Pix_766;
		PixelsStore[767] <= Pix_767;
		PixelsStore[768] <= Pix_768;
		PixelsStore[769] <= Pix_769;
		PixelsStore[770] <= Pix_770;
		PixelsStore[771] <= Pix_771;
		PixelsStore[772] <= Pix_772;
		PixelsStore[773] <= Pix_773;
		PixelsStore[774] <= Pix_774;
		PixelsStore[775] <= Pix_775;
		PixelsStore[776] <= Pix_776;
		PixelsStore[777] <= Pix_777;
		PixelsStore[778] <= Pix_778;
		PixelsStore[779] <= Pix_779;
		PixelsStore[780] <= Pix_780;
		PixelsStore[781] <= Pix_781;
		PixelsStore[782] <= Pix_782;
		PixelsStore[783] <= Pix_783;
		PixelsStore[784] <= Pix_784;
		WeightsStore0[0] <= Wgt_0_0;
		WeightsStore0[1] <= Wgt_0_1;
		WeightsStore0[2] <= Wgt_0_2;
		WeightsStore0[3] <= Wgt_0_3;
		WeightsStore0[4] <= Wgt_0_4;
		WeightsStore0[5] <= Wgt_0_5;
		WeightsStore0[6] <= Wgt_0_6;
		WeightsStore0[7] <= Wgt_0_7;
		WeightsStore0[8] <= Wgt_0_8;
		WeightsStore0[9] <= Wgt_0_9;
		WeightsStore0[10] <= Wgt_0_10;
		WeightsStore0[11] <= Wgt_0_11;
		WeightsStore0[12] <= Wgt_0_12;
		WeightsStore0[13] <= Wgt_0_13;
		WeightsStore0[14] <= Wgt_0_14;
		WeightsStore0[15] <= Wgt_0_15;
		WeightsStore0[16] <= Wgt_0_16;
		WeightsStore0[17] <= Wgt_0_17;
		WeightsStore0[18] <= Wgt_0_18;
		WeightsStore0[19] <= Wgt_0_19;
		WeightsStore0[20] <= Wgt_0_20;
		WeightsStore0[21] <= Wgt_0_21;
		WeightsStore0[22] <= Wgt_0_22;
		WeightsStore0[23] <= Wgt_0_23;
		WeightsStore0[24] <= Wgt_0_24;
		WeightsStore0[25] <= Wgt_0_25;
		WeightsStore0[26] <= Wgt_0_26;
		WeightsStore0[27] <= Wgt_0_27;
		WeightsStore0[28] <= Wgt_0_28;
		WeightsStore0[29] <= Wgt_0_29;
		WeightsStore0[30] <= Wgt_0_30;
		WeightsStore0[31] <= Wgt_0_31;
		WeightsStore0[32] <= Wgt_0_32;
		WeightsStore0[33] <= Wgt_0_33;
		WeightsStore0[34] <= Wgt_0_34;
		WeightsStore0[35] <= Wgt_0_35;
		WeightsStore0[36] <= Wgt_0_36;
		WeightsStore0[37] <= Wgt_0_37;
		WeightsStore0[38] <= Wgt_0_38;
		WeightsStore0[39] <= Wgt_0_39;
		WeightsStore0[40] <= Wgt_0_40;
		WeightsStore0[41] <= Wgt_0_41;
		WeightsStore0[42] <= Wgt_0_42;
		WeightsStore0[43] <= Wgt_0_43;
		WeightsStore0[44] <= Wgt_0_44;
		WeightsStore0[45] <= Wgt_0_45;
		WeightsStore0[46] <= Wgt_0_46;
		WeightsStore0[47] <= Wgt_0_47;
		WeightsStore0[48] <= Wgt_0_48;
		WeightsStore0[49] <= Wgt_0_49;
		WeightsStore0[50] <= Wgt_0_50;
		WeightsStore0[51] <= Wgt_0_51;
		WeightsStore0[52] <= Wgt_0_52;
		WeightsStore0[53] <= Wgt_0_53;
		WeightsStore0[54] <= Wgt_0_54;
		WeightsStore0[55] <= Wgt_0_55;
		WeightsStore0[56] <= Wgt_0_56;
		WeightsStore0[57] <= Wgt_0_57;
		WeightsStore0[58] <= Wgt_0_58;
		WeightsStore0[59] <= Wgt_0_59;
		WeightsStore0[60] <= Wgt_0_60;
		WeightsStore0[61] <= Wgt_0_61;
		WeightsStore0[62] <= Wgt_0_62;
		WeightsStore0[63] <= Wgt_0_63;
		WeightsStore0[64] <= Wgt_0_64;
		WeightsStore0[65] <= Wgt_0_65;
		WeightsStore0[66] <= Wgt_0_66;
		WeightsStore0[67] <= Wgt_0_67;
		WeightsStore0[68] <= Wgt_0_68;
		WeightsStore0[69] <= Wgt_0_69;
		WeightsStore0[70] <= Wgt_0_70;
		WeightsStore0[71] <= Wgt_0_71;
		WeightsStore0[72] <= Wgt_0_72;
		WeightsStore0[73] <= Wgt_0_73;
		WeightsStore0[74] <= Wgt_0_74;
		WeightsStore0[75] <= Wgt_0_75;
		WeightsStore0[76] <= Wgt_0_76;
		WeightsStore0[77] <= Wgt_0_77;
		WeightsStore0[78] <= Wgt_0_78;
		WeightsStore0[79] <= Wgt_0_79;
		WeightsStore0[80] <= Wgt_0_80;
		WeightsStore0[81] <= Wgt_0_81;
		WeightsStore0[82] <= Wgt_0_82;
		WeightsStore0[83] <= Wgt_0_83;
		WeightsStore0[84] <= Wgt_0_84;
		WeightsStore0[85] <= Wgt_0_85;
		WeightsStore0[86] <= Wgt_0_86;
		WeightsStore0[87] <= Wgt_0_87;
		WeightsStore0[88] <= Wgt_0_88;
		WeightsStore0[89] <= Wgt_0_89;
		WeightsStore0[90] <= Wgt_0_90;
		WeightsStore0[91] <= Wgt_0_91;
		WeightsStore0[92] <= Wgt_0_92;
		WeightsStore0[93] <= Wgt_0_93;
		WeightsStore0[94] <= Wgt_0_94;
		WeightsStore0[95] <= Wgt_0_95;
		WeightsStore0[96] <= Wgt_0_96;
		WeightsStore0[97] <= Wgt_0_97;
		WeightsStore0[98] <= Wgt_0_98;
		WeightsStore0[99] <= Wgt_0_99;
		WeightsStore0[100] <= Wgt_0_100;
		WeightsStore0[101] <= Wgt_0_101;
		WeightsStore0[102] <= Wgt_0_102;
		WeightsStore0[103] <= Wgt_0_103;
		WeightsStore0[104] <= Wgt_0_104;
		WeightsStore0[105] <= Wgt_0_105;
		WeightsStore0[106] <= Wgt_0_106;
		WeightsStore0[107] <= Wgt_0_107;
		WeightsStore0[108] <= Wgt_0_108;
		WeightsStore0[109] <= Wgt_0_109;
		WeightsStore0[110] <= Wgt_0_110;
		WeightsStore0[111] <= Wgt_0_111;
		WeightsStore0[112] <= Wgt_0_112;
		WeightsStore0[113] <= Wgt_0_113;
		WeightsStore0[114] <= Wgt_0_114;
		WeightsStore0[115] <= Wgt_0_115;
		WeightsStore0[116] <= Wgt_0_116;
		WeightsStore0[117] <= Wgt_0_117;
		WeightsStore0[118] <= Wgt_0_118;
		WeightsStore0[119] <= Wgt_0_119;
		WeightsStore0[120] <= Wgt_0_120;
		WeightsStore0[121] <= Wgt_0_121;
		WeightsStore0[122] <= Wgt_0_122;
		WeightsStore0[123] <= Wgt_0_123;
		WeightsStore0[124] <= Wgt_0_124;
		WeightsStore0[125] <= Wgt_0_125;
		WeightsStore0[126] <= Wgt_0_126;
		WeightsStore0[127] <= Wgt_0_127;
		WeightsStore0[128] <= Wgt_0_128;
		WeightsStore0[129] <= Wgt_0_129;
		WeightsStore0[130] <= Wgt_0_130;
		WeightsStore0[131] <= Wgt_0_131;
		WeightsStore0[132] <= Wgt_0_132;
		WeightsStore0[133] <= Wgt_0_133;
		WeightsStore0[134] <= Wgt_0_134;
		WeightsStore0[135] <= Wgt_0_135;
		WeightsStore0[136] <= Wgt_0_136;
		WeightsStore0[137] <= Wgt_0_137;
		WeightsStore0[138] <= Wgt_0_138;
		WeightsStore0[139] <= Wgt_0_139;
		WeightsStore0[140] <= Wgt_0_140;
		WeightsStore0[141] <= Wgt_0_141;
		WeightsStore0[142] <= Wgt_0_142;
		WeightsStore0[143] <= Wgt_0_143;
		WeightsStore0[144] <= Wgt_0_144;
		WeightsStore0[145] <= Wgt_0_145;
		WeightsStore0[146] <= Wgt_0_146;
		WeightsStore0[147] <= Wgt_0_147;
		WeightsStore0[148] <= Wgt_0_148;
		WeightsStore0[149] <= Wgt_0_149;
		WeightsStore0[150] <= Wgt_0_150;
		WeightsStore0[151] <= Wgt_0_151;
		WeightsStore0[152] <= Wgt_0_152;
		WeightsStore0[153] <= Wgt_0_153;
		WeightsStore0[154] <= Wgt_0_154;
		WeightsStore0[155] <= Wgt_0_155;
		WeightsStore0[156] <= Wgt_0_156;
		WeightsStore0[157] <= Wgt_0_157;
		WeightsStore0[158] <= Wgt_0_158;
		WeightsStore0[159] <= Wgt_0_159;
		WeightsStore0[160] <= Wgt_0_160;
		WeightsStore0[161] <= Wgt_0_161;
		WeightsStore0[162] <= Wgt_0_162;
		WeightsStore0[163] <= Wgt_0_163;
		WeightsStore0[164] <= Wgt_0_164;
		WeightsStore0[165] <= Wgt_0_165;
		WeightsStore0[166] <= Wgt_0_166;
		WeightsStore0[167] <= Wgt_0_167;
		WeightsStore0[168] <= Wgt_0_168;
		WeightsStore0[169] <= Wgt_0_169;
		WeightsStore0[170] <= Wgt_0_170;
		WeightsStore0[171] <= Wgt_0_171;
		WeightsStore0[172] <= Wgt_0_172;
		WeightsStore0[173] <= Wgt_0_173;
		WeightsStore0[174] <= Wgt_0_174;
		WeightsStore0[175] <= Wgt_0_175;
		WeightsStore0[176] <= Wgt_0_176;
		WeightsStore0[177] <= Wgt_0_177;
		WeightsStore0[178] <= Wgt_0_178;
		WeightsStore0[179] <= Wgt_0_179;
		WeightsStore0[180] <= Wgt_0_180;
		WeightsStore0[181] <= Wgt_0_181;
		WeightsStore0[182] <= Wgt_0_182;
		WeightsStore0[183] <= Wgt_0_183;
		WeightsStore0[184] <= Wgt_0_184;
		WeightsStore0[185] <= Wgt_0_185;
		WeightsStore0[186] <= Wgt_0_186;
		WeightsStore0[187] <= Wgt_0_187;
		WeightsStore0[188] <= Wgt_0_188;
		WeightsStore0[189] <= Wgt_0_189;
		WeightsStore0[190] <= Wgt_0_190;
		WeightsStore0[191] <= Wgt_0_191;
		WeightsStore0[192] <= Wgt_0_192;
		WeightsStore0[193] <= Wgt_0_193;
		WeightsStore0[194] <= Wgt_0_194;
		WeightsStore0[195] <= Wgt_0_195;
		WeightsStore0[196] <= Wgt_0_196;
		WeightsStore0[197] <= Wgt_0_197;
		WeightsStore0[198] <= Wgt_0_198;
		WeightsStore0[199] <= Wgt_0_199;
		WeightsStore0[200] <= Wgt_0_200;
		WeightsStore0[201] <= Wgt_0_201;
		WeightsStore0[202] <= Wgt_0_202;
		WeightsStore0[203] <= Wgt_0_203;
		WeightsStore0[204] <= Wgt_0_204;
		WeightsStore0[205] <= Wgt_0_205;
		WeightsStore0[206] <= Wgt_0_206;
		WeightsStore0[207] <= Wgt_0_207;
		WeightsStore0[208] <= Wgt_0_208;
		WeightsStore0[209] <= Wgt_0_209;
		WeightsStore0[210] <= Wgt_0_210;
		WeightsStore0[211] <= Wgt_0_211;
		WeightsStore0[212] <= Wgt_0_212;
		WeightsStore0[213] <= Wgt_0_213;
		WeightsStore0[214] <= Wgt_0_214;
		WeightsStore0[215] <= Wgt_0_215;
		WeightsStore0[216] <= Wgt_0_216;
		WeightsStore0[217] <= Wgt_0_217;
		WeightsStore0[218] <= Wgt_0_218;
		WeightsStore0[219] <= Wgt_0_219;
		WeightsStore0[220] <= Wgt_0_220;
		WeightsStore0[221] <= Wgt_0_221;
		WeightsStore0[222] <= Wgt_0_222;
		WeightsStore0[223] <= Wgt_0_223;
		WeightsStore0[224] <= Wgt_0_224;
		WeightsStore0[225] <= Wgt_0_225;
		WeightsStore0[226] <= Wgt_0_226;
		WeightsStore0[227] <= Wgt_0_227;
		WeightsStore0[228] <= Wgt_0_228;
		WeightsStore0[229] <= Wgt_0_229;
		WeightsStore0[230] <= Wgt_0_230;
		WeightsStore0[231] <= Wgt_0_231;
		WeightsStore0[232] <= Wgt_0_232;
		WeightsStore0[233] <= Wgt_0_233;
		WeightsStore0[234] <= Wgt_0_234;
		WeightsStore0[235] <= Wgt_0_235;
		WeightsStore0[236] <= Wgt_0_236;
		WeightsStore0[237] <= Wgt_0_237;
		WeightsStore0[238] <= Wgt_0_238;
		WeightsStore0[239] <= Wgt_0_239;
		WeightsStore0[240] <= Wgt_0_240;
		WeightsStore0[241] <= Wgt_0_241;
		WeightsStore0[242] <= Wgt_0_242;
		WeightsStore0[243] <= Wgt_0_243;
		WeightsStore0[244] <= Wgt_0_244;
		WeightsStore0[245] <= Wgt_0_245;
		WeightsStore0[246] <= Wgt_0_246;
		WeightsStore0[247] <= Wgt_0_247;
		WeightsStore0[248] <= Wgt_0_248;
		WeightsStore0[249] <= Wgt_0_249;
		WeightsStore0[250] <= Wgt_0_250;
		WeightsStore0[251] <= Wgt_0_251;
		WeightsStore0[252] <= Wgt_0_252;
		WeightsStore0[253] <= Wgt_0_253;
		WeightsStore0[254] <= Wgt_0_254;
		WeightsStore0[255] <= Wgt_0_255;
		WeightsStore0[256] <= Wgt_0_256;
		WeightsStore0[257] <= Wgt_0_257;
		WeightsStore0[258] <= Wgt_0_258;
		WeightsStore0[259] <= Wgt_0_259;
		WeightsStore0[260] <= Wgt_0_260;
		WeightsStore0[261] <= Wgt_0_261;
		WeightsStore0[262] <= Wgt_0_262;
		WeightsStore0[263] <= Wgt_0_263;
		WeightsStore0[264] <= Wgt_0_264;
		WeightsStore0[265] <= Wgt_0_265;
		WeightsStore0[266] <= Wgt_0_266;
		WeightsStore0[267] <= Wgt_0_267;
		WeightsStore0[268] <= Wgt_0_268;
		WeightsStore0[269] <= Wgt_0_269;
		WeightsStore0[270] <= Wgt_0_270;
		WeightsStore0[271] <= Wgt_0_271;
		WeightsStore0[272] <= Wgt_0_272;
		WeightsStore0[273] <= Wgt_0_273;
		WeightsStore0[274] <= Wgt_0_274;
		WeightsStore0[275] <= Wgt_0_275;
		WeightsStore0[276] <= Wgt_0_276;
		WeightsStore0[277] <= Wgt_0_277;
		WeightsStore0[278] <= Wgt_0_278;
		WeightsStore0[279] <= Wgt_0_279;
		WeightsStore0[280] <= Wgt_0_280;
		WeightsStore0[281] <= Wgt_0_281;
		WeightsStore0[282] <= Wgt_0_282;
		WeightsStore0[283] <= Wgt_0_283;
		WeightsStore0[284] <= Wgt_0_284;
		WeightsStore0[285] <= Wgt_0_285;
		WeightsStore0[286] <= Wgt_0_286;
		WeightsStore0[287] <= Wgt_0_287;
		WeightsStore0[288] <= Wgt_0_288;
		WeightsStore0[289] <= Wgt_0_289;
		WeightsStore0[290] <= Wgt_0_290;
		WeightsStore0[291] <= Wgt_0_291;
		WeightsStore0[292] <= Wgt_0_292;
		WeightsStore0[293] <= Wgt_0_293;
		WeightsStore0[294] <= Wgt_0_294;
		WeightsStore0[295] <= Wgt_0_295;
		WeightsStore0[296] <= Wgt_0_296;
		WeightsStore0[297] <= Wgt_0_297;
		WeightsStore0[298] <= Wgt_0_298;
		WeightsStore0[299] <= Wgt_0_299;
		WeightsStore0[300] <= Wgt_0_300;
		WeightsStore0[301] <= Wgt_0_301;
		WeightsStore0[302] <= Wgt_0_302;
		WeightsStore0[303] <= Wgt_0_303;
		WeightsStore0[304] <= Wgt_0_304;
		WeightsStore0[305] <= Wgt_0_305;
		WeightsStore0[306] <= Wgt_0_306;
		WeightsStore0[307] <= Wgt_0_307;
		WeightsStore0[308] <= Wgt_0_308;
		WeightsStore0[309] <= Wgt_0_309;
		WeightsStore0[310] <= Wgt_0_310;
		WeightsStore0[311] <= Wgt_0_311;
		WeightsStore0[312] <= Wgt_0_312;
		WeightsStore0[313] <= Wgt_0_313;
		WeightsStore0[314] <= Wgt_0_314;
		WeightsStore0[315] <= Wgt_0_315;
		WeightsStore0[316] <= Wgt_0_316;
		WeightsStore0[317] <= Wgt_0_317;
		WeightsStore0[318] <= Wgt_0_318;
		WeightsStore0[319] <= Wgt_0_319;
		WeightsStore0[320] <= Wgt_0_320;
		WeightsStore0[321] <= Wgt_0_321;
		WeightsStore0[322] <= Wgt_0_322;
		WeightsStore0[323] <= Wgt_0_323;
		WeightsStore0[324] <= Wgt_0_324;
		WeightsStore0[325] <= Wgt_0_325;
		WeightsStore0[326] <= Wgt_0_326;
		WeightsStore0[327] <= Wgt_0_327;
		WeightsStore0[328] <= Wgt_0_328;
		WeightsStore0[329] <= Wgt_0_329;
		WeightsStore0[330] <= Wgt_0_330;
		WeightsStore0[331] <= Wgt_0_331;
		WeightsStore0[332] <= Wgt_0_332;
		WeightsStore0[333] <= Wgt_0_333;
		WeightsStore0[334] <= Wgt_0_334;
		WeightsStore0[335] <= Wgt_0_335;
		WeightsStore0[336] <= Wgt_0_336;
		WeightsStore0[337] <= Wgt_0_337;
		WeightsStore0[338] <= Wgt_0_338;
		WeightsStore0[339] <= Wgt_0_339;
		WeightsStore0[340] <= Wgt_0_340;
		WeightsStore0[341] <= Wgt_0_341;
		WeightsStore0[342] <= Wgt_0_342;
		WeightsStore0[343] <= Wgt_0_343;
		WeightsStore0[344] <= Wgt_0_344;
		WeightsStore0[345] <= Wgt_0_345;
		WeightsStore0[346] <= Wgt_0_346;
		WeightsStore0[347] <= Wgt_0_347;
		WeightsStore0[348] <= Wgt_0_348;
		WeightsStore0[349] <= Wgt_0_349;
		WeightsStore0[350] <= Wgt_0_350;
		WeightsStore0[351] <= Wgt_0_351;
		WeightsStore0[352] <= Wgt_0_352;
		WeightsStore0[353] <= Wgt_0_353;
		WeightsStore0[354] <= Wgt_0_354;
		WeightsStore0[355] <= Wgt_0_355;
		WeightsStore0[356] <= Wgt_0_356;
		WeightsStore0[357] <= Wgt_0_357;
		WeightsStore0[358] <= Wgt_0_358;
		WeightsStore0[359] <= Wgt_0_359;
		WeightsStore0[360] <= Wgt_0_360;
		WeightsStore0[361] <= Wgt_0_361;
		WeightsStore0[362] <= Wgt_0_362;
		WeightsStore0[363] <= Wgt_0_363;
		WeightsStore0[364] <= Wgt_0_364;
		WeightsStore0[365] <= Wgt_0_365;
		WeightsStore0[366] <= Wgt_0_366;
		WeightsStore0[367] <= Wgt_0_367;
		WeightsStore0[368] <= Wgt_0_368;
		WeightsStore0[369] <= Wgt_0_369;
		WeightsStore0[370] <= Wgt_0_370;
		WeightsStore0[371] <= Wgt_0_371;
		WeightsStore0[372] <= Wgt_0_372;
		WeightsStore0[373] <= Wgt_0_373;
		WeightsStore0[374] <= Wgt_0_374;
		WeightsStore0[375] <= Wgt_0_375;
		WeightsStore0[376] <= Wgt_0_376;
		WeightsStore0[377] <= Wgt_0_377;
		WeightsStore0[378] <= Wgt_0_378;
		WeightsStore0[379] <= Wgt_0_379;
		WeightsStore0[380] <= Wgt_0_380;
		WeightsStore0[381] <= Wgt_0_381;
		WeightsStore0[382] <= Wgt_0_382;
		WeightsStore0[383] <= Wgt_0_383;
		WeightsStore0[384] <= Wgt_0_384;
		WeightsStore0[385] <= Wgt_0_385;
		WeightsStore0[386] <= Wgt_0_386;
		WeightsStore0[387] <= Wgt_0_387;
		WeightsStore0[388] <= Wgt_0_388;
		WeightsStore0[389] <= Wgt_0_389;
		WeightsStore0[390] <= Wgt_0_390;
		WeightsStore0[391] <= Wgt_0_391;
		WeightsStore0[392] <= Wgt_0_392;
		WeightsStore0[393] <= Wgt_0_393;
		WeightsStore0[394] <= Wgt_0_394;
		WeightsStore0[395] <= Wgt_0_395;
		WeightsStore0[396] <= Wgt_0_396;
		WeightsStore0[397] <= Wgt_0_397;
		WeightsStore0[398] <= Wgt_0_398;
		WeightsStore0[399] <= Wgt_0_399;
		WeightsStore0[400] <= Wgt_0_400;
		WeightsStore0[401] <= Wgt_0_401;
		WeightsStore0[402] <= Wgt_0_402;
		WeightsStore0[403] <= Wgt_0_403;
		WeightsStore0[404] <= Wgt_0_404;
		WeightsStore0[405] <= Wgt_0_405;
		WeightsStore0[406] <= Wgt_0_406;
		WeightsStore0[407] <= Wgt_0_407;
		WeightsStore0[408] <= Wgt_0_408;
		WeightsStore0[409] <= Wgt_0_409;
		WeightsStore0[410] <= Wgt_0_410;
		WeightsStore0[411] <= Wgt_0_411;
		WeightsStore0[412] <= Wgt_0_412;
		WeightsStore0[413] <= Wgt_0_413;
		WeightsStore0[414] <= Wgt_0_414;
		WeightsStore0[415] <= Wgt_0_415;
		WeightsStore0[416] <= Wgt_0_416;
		WeightsStore0[417] <= Wgt_0_417;
		WeightsStore0[418] <= Wgt_0_418;
		WeightsStore0[419] <= Wgt_0_419;
		WeightsStore0[420] <= Wgt_0_420;
		WeightsStore0[421] <= Wgt_0_421;
		WeightsStore0[422] <= Wgt_0_422;
		WeightsStore0[423] <= Wgt_0_423;
		WeightsStore0[424] <= Wgt_0_424;
		WeightsStore0[425] <= Wgt_0_425;
		WeightsStore0[426] <= Wgt_0_426;
		WeightsStore0[427] <= Wgt_0_427;
		WeightsStore0[428] <= Wgt_0_428;
		WeightsStore0[429] <= Wgt_0_429;
		WeightsStore0[430] <= Wgt_0_430;
		WeightsStore0[431] <= Wgt_0_431;
		WeightsStore0[432] <= Wgt_0_432;
		WeightsStore0[433] <= Wgt_0_433;
		WeightsStore0[434] <= Wgt_0_434;
		WeightsStore0[435] <= Wgt_0_435;
		WeightsStore0[436] <= Wgt_0_436;
		WeightsStore0[437] <= Wgt_0_437;
		WeightsStore0[438] <= Wgt_0_438;
		WeightsStore0[439] <= Wgt_0_439;
		WeightsStore0[440] <= Wgt_0_440;
		WeightsStore0[441] <= Wgt_0_441;
		WeightsStore0[442] <= Wgt_0_442;
		WeightsStore0[443] <= Wgt_0_443;
		WeightsStore0[444] <= Wgt_0_444;
		WeightsStore0[445] <= Wgt_0_445;
		WeightsStore0[446] <= Wgt_0_446;
		WeightsStore0[447] <= Wgt_0_447;
		WeightsStore0[448] <= Wgt_0_448;
		WeightsStore0[449] <= Wgt_0_449;
		WeightsStore0[450] <= Wgt_0_450;
		WeightsStore0[451] <= Wgt_0_451;
		WeightsStore0[452] <= Wgt_0_452;
		WeightsStore0[453] <= Wgt_0_453;
		WeightsStore0[454] <= Wgt_0_454;
		WeightsStore0[455] <= Wgt_0_455;
		WeightsStore0[456] <= Wgt_0_456;
		WeightsStore0[457] <= Wgt_0_457;
		WeightsStore0[458] <= Wgt_0_458;
		WeightsStore0[459] <= Wgt_0_459;
		WeightsStore0[460] <= Wgt_0_460;
		WeightsStore0[461] <= Wgt_0_461;
		WeightsStore0[462] <= Wgt_0_462;
		WeightsStore0[463] <= Wgt_0_463;
		WeightsStore0[464] <= Wgt_0_464;
		WeightsStore0[465] <= Wgt_0_465;
		WeightsStore0[466] <= Wgt_0_466;
		WeightsStore0[467] <= Wgt_0_467;
		WeightsStore0[468] <= Wgt_0_468;
		WeightsStore0[469] <= Wgt_0_469;
		WeightsStore0[470] <= Wgt_0_470;
		WeightsStore0[471] <= Wgt_0_471;
		WeightsStore0[472] <= Wgt_0_472;
		WeightsStore0[473] <= Wgt_0_473;
		WeightsStore0[474] <= Wgt_0_474;
		WeightsStore0[475] <= Wgt_0_475;
		WeightsStore0[476] <= Wgt_0_476;
		WeightsStore0[477] <= Wgt_0_477;
		WeightsStore0[478] <= Wgt_0_478;
		WeightsStore0[479] <= Wgt_0_479;
		WeightsStore0[480] <= Wgt_0_480;
		WeightsStore0[481] <= Wgt_0_481;
		WeightsStore0[482] <= Wgt_0_482;
		WeightsStore0[483] <= Wgt_0_483;
		WeightsStore0[484] <= Wgt_0_484;
		WeightsStore0[485] <= Wgt_0_485;
		WeightsStore0[486] <= Wgt_0_486;
		WeightsStore0[487] <= Wgt_0_487;
		WeightsStore0[488] <= Wgt_0_488;
		WeightsStore0[489] <= Wgt_0_489;
		WeightsStore0[490] <= Wgt_0_490;
		WeightsStore0[491] <= Wgt_0_491;
		WeightsStore0[492] <= Wgt_0_492;
		WeightsStore0[493] <= Wgt_0_493;
		WeightsStore0[494] <= Wgt_0_494;
		WeightsStore0[495] <= Wgt_0_495;
		WeightsStore0[496] <= Wgt_0_496;
		WeightsStore0[497] <= Wgt_0_497;
		WeightsStore0[498] <= Wgt_0_498;
		WeightsStore0[499] <= Wgt_0_499;
		WeightsStore0[500] <= Wgt_0_500;
		WeightsStore0[501] <= Wgt_0_501;
		WeightsStore0[502] <= Wgt_0_502;
		WeightsStore0[503] <= Wgt_0_503;
		WeightsStore0[504] <= Wgt_0_504;
		WeightsStore0[505] <= Wgt_0_505;
		WeightsStore0[506] <= Wgt_0_506;
		WeightsStore0[507] <= Wgt_0_507;
		WeightsStore0[508] <= Wgt_0_508;
		WeightsStore0[509] <= Wgt_0_509;
		WeightsStore0[510] <= Wgt_0_510;
		WeightsStore0[511] <= Wgt_0_511;
		WeightsStore0[512] <= Wgt_0_512;
		WeightsStore0[513] <= Wgt_0_513;
		WeightsStore0[514] <= Wgt_0_514;
		WeightsStore0[515] <= Wgt_0_515;
		WeightsStore0[516] <= Wgt_0_516;
		WeightsStore0[517] <= Wgt_0_517;
		WeightsStore0[518] <= Wgt_0_518;
		WeightsStore0[519] <= Wgt_0_519;
		WeightsStore0[520] <= Wgt_0_520;
		WeightsStore0[521] <= Wgt_0_521;
		WeightsStore0[522] <= Wgt_0_522;
		WeightsStore0[523] <= Wgt_0_523;
		WeightsStore0[524] <= Wgt_0_524;
		WeightsStore0[525] <= Wgt_0_525;
		WeightsStore0[526] <= Wgt_0_526;
		WeightsStore0[527] <= Wgt_0_527;
		WeightsStore0[528] <= Wgt_0_528;
		WeightsStore0[529] <= Wgt_0_529;
		WeightsStore0[530] <= Wgt_0_530;
		WeightsStore0[531] <= Wgt_0_531;
		WeightsStore0[532] <= Wgt_0_532;
		WeightsStore0[533] <= Wgt_0_533;
		WeightsStore0[534] <= Wgt_0_534;
		WeightsStore0[535] <= Wgt_0_535;
		WeightsStore0[536] <= Wgt_0_536;
		WeightsStore0[537] <= Wgt_0_537;
		WeightsStore0[538] <= Wgt_0_538;
		WeightsStore0[539] <= Wgt_0_539;
		WeightsStore0[540] <= Wgt_0_540;
		WeightsStore0[541] <= Wgt_0_541;
		WeightsStore0[542] <= Wgt_0_542;
		WeightsStore0[543] <= Wgt_0_543;
		WeightsStore0[544] <= Wgt_0_544;
		WeightsStore0[545] <= Wgt_0_545;
		WeightsStore0[546] <= Wgt_0_546;
		WeightsStore0[547] <= Wgt_0_547;
		WeightsStore0[548] <= Wgt_0_548;
		WeightsStore0[549] <= Wgt_0_549;
		WeightsStore0[550] <= Wgt_0_550;
		WeightsStore0[551] <= Wgt_0_551;
		WeightsStore0[552] <= Wgt_0_552;
		WeightsStore0[553] <= Wgt_0_553;
		WeightsStore0[554] <= Wgt_0_554;
		WeightsStore0[555] <= Wgt_0_555;
		WeightsStore0[556] <= Wgt_0_556;
		WeightsStore0[557] <= Wgt_0_557;
		WeightsStore0[558] <= Wgt_0_558;
		WeightsStore0[559] <= Wgt_0_559;
		WeightsStore0[560] <= Wgt_0_560;
		WeightsStore0[561] <= Wgt_0_561;
		WeightsStore0[562] <= Wgt_0_562;
		WeightsStore0[563] <= Wgt_0_563;
		WeightsStore0[564] <= Wgt_0_564;
		WeightsStore0[565] <= Wgt_0_565;
		WeightsStore0[566] <= Wgt_0_566;
		WeightsStore0[567] <= Wgt_0_567;
		WeightsStore0[568] <= Wgt_0_568;
		WeightsStore0[569] <= Wgt_0_569;
		WeightsStore0[570] <= Wgt_0_570;
		WeightsStore0[571] <= Wgt_0_571;
		WeightsStore0[572] <= Wgt_0_572;
		WeightsStore0[573] <= Wgt_0_573;
		WeightsStore0[574] <= Wgt_0_574;
		WeightsStore0[575] <= Wgt_0_575;
		WeightsStore0[576] <= Wgt_0_576;
		WeightsStore0[577] <= Wgt_0_577;
		WeightsStore0[578] <= Wgt_0_578;
		WeightsStore0[579] <= Wgt_0_579;
		WeightsStore0[580] <= Wgt_0_580;
		WeightsStore0[581] <= Wgt_0_581;
		WeightsStore0[582] <= Wgt_0_582;
		WeightsStore0[583] <= Wgt_0_583;
		WeightsStore0[584] <= Wgt_0_584;
		WeightsStore0[585] <= Wgt_0_585;
		WeightsStore0[586] <= Wgt_0_586;
		WeightsStore0[587] <= Wgt_0_587;
		WeightsStore0[588] <= Wgt_0_588;
		WeightsStore0[589] <= Wgt_0_589;
		WeightsStore0[590] <= Wgt_0_590;
		WeightsStore0[591] <= Wgt_0_591;
		WeightsStore0[592] <= Wgt_0_592;
		WeightsStore0[593] <= Wgt_0_593;
		WeightsStore0[594] <= Wgt_0_594;
		WeightsStore0[595] <= Wgt_0_595;
		WeightsStore0[596] <= Wgt_0_596;
		WeightsStore0[597] <= Wgt_0_597;
		WeightsStore0[598] <= Wgt_0_598;
		WeightsStore0[599] <= Wgt_0_599;
		WeightsStore0[600] <= Wgt_0_600;
		WeightsStore0[601] <= Wgt_0_601;
		WeightsStore0[602] <= Wgt_0_602;
		WeightsStore0[603] <= Wgt_0_603;
		WeightsStore0[604] <= Wgt_0_604;
		WeightsStore0[605] <= Wgt_0_605;
		WeightsStore0[606] <= Wgt_0_606;
		WeightsStore0[607] <= Wgt_0_607;
		WeightsStore0[608] <= Wgt_0_608;
		WeightsStore0[609] <= Wgt_0_609;
		WeightsStore0[610] <= Wgt_0_610;
		WeightsStore0[611] <= Wgt_0_611;
		WeightsStore0[612] <= Wgt_0_612;
		WeightsStore0[613] <= Wgt_0_613;
		WeightsStore0[614] <= Wgt_0_614;
		WeightsStore0[615] <= Wgt_0_615;
		WeightsStore0[616] <= Wgt_0_616;
		WeightsStore0[617] <= Wgt_0_617;
		WeightsStore0[618] <= Wgt_0_618;
		WeightsStore0[619] <= Wgt_0_619;
		WeightsStore0[620] <= Wgt_0_620;
		WeightsStore0[621] <= Wgt_0_621;
		WeightsStore0[622] <= Wgt_0_622;
		WeightsStore0[623] <= Wgt_0_623;
		WeightsStore0[624] <= Wgt_0_624;
		WeightsStore0[625] <= Wgt_0_625;
		WeightsStore0[626] <= Wgt_0_626;
		WeightsStore0[627] <= Wgt_0_627;
		WeightsStore0[628] <= Wgt_0_628;
		WeightsStore0[629] <= Wgt_0_629;
		WeightsStore0[630] <= Wgt_0_630;
		WeightsStore0[631] <= Wgt_0_631;
		WeightsStore0[632] <= Wgt_0_632;
		WeightsStore0[633] <= Wgt_0_633;
		WeightsStore0[634] <= Wgt_0_634;
		WeightsStore0[635] <= Wgt_0_635;
		WeightsStore0[636] <= Wgt_0_636;
		WeightsStore0[637] <= Wgt_0_637;
		WeightsStore0[638] <= Wgt_0_638;
		WeightsStore0[639] <= Wgt_0_639;
		WeightsStore0[640] <= Wgt_0_640;
		WeightsStore0[641] <= Wgt_0_641;
		WeightsStore0[642] <= Wgt_0_642;
		WeightsStore0[643] <= Wgt_0_643;
		WeightsStore0[644] <= Wgt_0_644;
		WeightsStore0[645] <= Wgt_0_645;
		WeightsStore0[646] <= Wgt_0_646;
		WeightsStore0[647] <= Wgt_0_647;
		WeightsStore0[648] <= Wgt_0_648;
		WeightsStore0[649] <= Wgt_0_649;
		WeightsStore0[650] <= Wgt_0_650;
		WeightsStore0[651] <= Wgt_0_651;
		WeightsStore0[652] <= Wgt_0_652;
		WeightsStore0[653] <= Wgt_0_653;
		WeightsStore0[654] <= Wgt_0_654;
		WeightsStore0[655] <= Wgt_0_655;
		WeightsStore0[656] <= Wgt_0_656;
		WeightsStore0[657] <= Wgt_0_657;
		WeightsStore0[658] <= Wgt_0_658;
		WeightsStore0[659] <= Wgt_0_659;
		WeightsStore0[660] <= Wgt_0_660;
		WeightsStore0[661] <= Wgt_0_661;
		WeightsStore0[662] <= Wgt_0_662;
		WeightsStore0[663] <= Wgt_0_663;
		WeightsStore0[664] <= Wgt_0_664;
		WeightsStore0[665] <= Wgt_0_665;
		WeightsStore0[666] <= Wgt_0_666;
		WeightsStore0[667] <= Wgt_0_667;
		WeightsStore0[668] <= Wgt_0_668;
		WeightsStore0[669] <= Wgt_0_669;
		WeightsStore0[670] <= Wgt_0_670;
		WeightsStore0[671] <= Wgt_0_671;
		WeightsStore0[672] <= Wgt_0_672;
		WeightsStore0[673] <= Wgt_0_673;
		WeightsStore0[674] <= Wgt_0_674;
		WeightsStore0[675] <= Wgt_0_675;
		WeightsStore0[676] <= Wgt_0_676;
		WeightsStore0[677] <= Wgt_0_677;
		WeightsStore0[678] <= Wgt_0_678;
		WeightsStore0[679] <= Wgt_0_679;
		WeightsStore0[680] <= Wgt_0_680;
		WeightsStore0[681] <= Wgt_0_681;
		WeightsStore0[682] <= Wgt_0_682;
		WeightsStore0[683] <= Wgt_0_683;
		WeightsStore0[684] <= Wgt_0_684;
		WeightsStore0[685] <= Wgt_0_685;
		WeightsStore0[686] <= Wgt_0_686;
		WeightsStore0[687] <= Wgt_0_687;
		WeightsStore0[688] <= Wgt_0_688;
		WeightsStore0[689] <= Wgt_0_689;
		WeightsStore0[690] <= Wgt_0_690;
		WeightsStore0[691] <= Wgt_0_691;
		WeightsStore0[692] <= Wgt_0_692;
		WeightsStore0[693] <= Wgt_0_693;
		WeightsStore0[694] <= Wgt_0_694;
		WeightsStore0[695] <= Wgt_0_695;
		WeightsStore0[696] <= Wgt_0_696;
		WeightsStore0[697] <= Wgt_0_697;
		WeightsStore0[698] <= Wgt_0_698;
		WeightsStore0[699] <= Wgt_0_699;
		WeightsStore0[700] <= Wgt_0_700;
		WeightsStore0[701] <= Wgt_0_701;
		WeightsStore0[702] <= Wgt_0_702;
		WeightsStore0[703] <= Wgt_0_703;
		WeightsStore0[704] <= Wgt_0_704;
		WeightsStore0[705] <= Wgt_0_705;
		WeightsStore0[706] <= Wgt_0_706;
		WeightsStore0[707] <= Wgt_0_707;
		WeightsStore0[708] <= Wgt_0_708;
		WeightsStore0[709] <= Wgt_0_709;
		WeightsStore0[710] <= Wgt_0_710;
		WeightsStore0[711] <= Wgt_0_711;
		WeightsStore0[712] <= Wgt_0_712;
		WeightsStore0[713] <= Wgt_0_713;
		WeightsStore0[714] <= Wgt_0_714;
		WeightsStore0[715] <= Wgt_0_715;
		WeightsStore0[716] <= Wgt_0_716;
		WeightsStore0[717] <= Wgt_0_717;
		WeightsStore0[718] <= Wgt_0_718;
		WeightsStore0[719] <= Wgt_0_719;
		WeightsStore0[720] <= Wgt_0_720;
		WeightsStore0[721] <= Wgt_0_721;
		WeightsStore0[722] <= Wgt_0_722;
		WeightsStore0[723] <= Wgt_0_723;
		WeightsStore0[724] <= Wgt_0_724;
		WeightsStore0[725] <= Wgt_0_725;
		WeightsStore0[726] <= Wgt_0_726;
		WeightsStore0[727] <= Wgt_0_727;
		WeightsStore0[728] <= Wgt_0_728;
		WeightsStore0[729] <= Wgt_0_729;
		WeightsStore0[730] <= Wgt_0_730;
		WeightsStore0[731] <= Wgt_0_731;
		WeightsStore0[732] <= Wgt_0_732;
		WeightsStore0[733] <= Wgt_0_733;
		WeightsStore0[734] <= Wgt_0_734;
		WeightsStore0[735] <= Wgt_0_735;
		WeightsStore0[736] <= Wgt_0_736;
		WeightsStore0[737] <= Wgt_0_737;
		WeightsStore0[738] <= Wgt_0_738;
		WeightsStore0[739] <= Wgt_0_739;
		WeightsStore0[740] <= Wgt_0_740;
		WeightsStore0[741] <= Wgt_0_741;
		WeightsStore0[742] <= Wgt_0_742;
		WeightsStore0[743] <= Wgt_0_743;
		WeightsStore0[744] <= Wgt_0_744;
		WeightsStore0[745] <= Wgt_0_745;
		WeightsStore0[746] <= Wgt_0_746;
		WeightsStore0[747] <= Wgt_0_747;
		WeightsStore0[748] <= Wgt_0_748;
		WeightsStore0[749] <= Wgt_0_749;
		WeightsStore0[750] <= Wgt_0_750;
		WeightsStore0[751] <= Wgt_0_751;
		WeightsStore0[752] <= Wgt_0_752;
		WeightsStore0[753] <= Wgt_0_753;
		WeightsStore0[754] <= Wgt_0_754;
		WeightsStore0[755] <= Wgt_0_755;
		WeightsStore0[756] <= Wgt_0_756;
		WeightsStore0[757] <= Wgt_0_757;
		WeightsStore0[758] <= Wgt_0_758;
		WeightsStore0[759] <= Wgt_0_759;
		WeightsStore0[760] <= Wgt_0_760;
		WeightsStore0[761] <= Wgt_0_761;
		WeightsStore0[762] <= Wgt_0_762;
		WeightsStore0[763] <= Wgt_0_763;
		WeightsStore0[764] <= Wgt_0_764;
		WeightsStore0[765] <= Wgt_0_765;
		WeightsStore0[766] <= Wgt_0_766;
		WeightsStore0[767] <= Wgt_0_767;
		WeightsStore0[768] <= Wgt_0_768;
		WeightsStore0[769] <= Wgt_0_769;
		WeightsStore0[770] <= Wgt_0_770;
		WeightsStore0[771] <= Wgt_0_771;
		WeightsStore0[772] <= Wgt_0_772;
		WeightsStore0[773] <= Wgt_0_773;
		WeightsStore0[774] <= Wgt_0_774;
		WeightsStore0[775] <= Wgt_0_775;
		WeightsStore0[776] <= Wgt_0_776;
		WeightsStore0[777] <= Wgt_0_777;
		WeightsStore0[778] <= Wgt_0_778;
		WeightsStore0[779] <= Wgt_0_779;
		WeightsStore0[780] <= Wgt_0_780;
		WeightsStore0[781] <= Wgt_0_781;
		WeightsStore0[782] <= Wgt_0_782;
		WeightsStore0[783] <= Wgt_0_783;
		WeightsStore0[784] <= Wgt_0_784;
		WeightsStore1[0] <= Wgt_1_0;
		WeightsStore1[1] <= Wgt_1_1;
		WeightsStore1[2] <= Wgt_1_2;
		WeightsStore1[3] <= Wgt_1_3;
		WeightsStore1[4] <= Wgt_1_4;
		WeightsStore1[5] <= Wgt_1_5;
		WeightsStore1[6] <= Wgt_1_6;
		WeightsStore1[7] <= Wgt_1_7;
		WeightsStore1[8] <= Wgt_1_8;
		WeightsStore1[9] <= Wgt_1_9;
		WeightsStore1[10] <= Wgt_1_10;
		WeightsStore1[11] <= Wgt_1_11;
		WeightsStore1[12] <= Wgt_1_12;
		WeightsStore1[13] <= Wgt_1_13;
		WeightsStore1[14] <= Wgt_1_14;
		WeightsStore1[15] <= Wgt_1_15;
		WeightsStore1[16] <= Wgt_1_16;
		WeightsStore1[17] <= Wgt_1_17;
		WeightsStore1[18] <= Wgt_1_18;
		WeightsStore1[19] <= Wgt_1_19;
		WeightsStore1[20] <= Wgt_1_20;
		WeightsStore1[21] <= Wgt_1_21;
		WeightsStore1[22] <= Wgt_1_22;
		WeightsStore1[23] <= Wgt_1_23;
		WeightsStore1[24] <= Wgt_1_24;
		WeightsStore1[25] <= Wgt_1_25;
		WeightsStore1[26] <= Wgt_1_26;
		WeightsStore1[27] <= Wgt_1_27;
		WeightsStore1[28] <= Wgt_1_28;
		WeightsStore1[29] <= Wgt_1_29;
		WeightsStore1[30] <= Wgt_1_30;
		WeightsStore1[31] <= Wgt_1_31;
		WeightsStore1[32] <= Wgt_1_32;
		WeightsStore1[33] <= Wgt_1_33;
		WeightsStore1[34] <= Wgt_1_34;
		WeightsStore1[35] <= Wgt_1_35;
		WeightsStore1[36] <= Wgt_1_36;
		WeightsStore1[37] <= Wgt_1_37;
		WeightsStore1[38] <= Wgt_1_38;
		WeightsStore1[39] <= Wgt_1_39;
		WeightsStore1[40] <= Wgt_1_40;
		WeightsStore1[41] <= Wgt_1_41;
		WeightsStore1[42] <= Wgt_1_42;
		WeightsStore1[43] <= Wgt_1_43;
		WeightsStore1[44] <= Wgt_1_44;
		WeightsStore1[45] <= Wgt_1_45;
		WeightsStore1[46] <= Wgt_1_46;
		WeightsStore1[47] <= Wgt_1_47;
		WeightsStore1[48] <= Wgt_1_48;
		WeightsStore1[49] <= Wgt_1_49;
		WeightsStore1[50] <= Wgt_1_50;
		WeightsStore1[51] <= Wgt_1_51;
		WeightsStore1[52] <= Wgt_1_52;
		WeightsStore1[53] <= Wgt_1_53;
		WeightsStore1[54] <= Wgt_1_54;
		WeightsStore1[55] <= Wgt_1_55;
		WeightsStore1[56] <= Wgt_1_56;
		WeightsStore1[57] <= Wgt_1_57;
		WeightsStore1[58] <= Wgt_1_58;
		WeightsStore1[59] <= Wgt_1_59;
		WeightsStore1[60] <= Wgt_1_60;
		WeightsStore1[61] <= Wgt_1_61;
		WeightsStore1[62] <= Wgt_1_62;
		WeightsStore1[63] <= Wgt_1_63;
		WeightsStore1[64] <= Wgt_1_64;
		WeightsStore1[65] <= Wgt_1_65;
		WeightsStore1[66] <= Wgt_1_66;
		WeightsStore1[67] <= Wgt_1_67;
		WeightsStore1[68] <= Wgt_1_68;
		WeightsStore1[69] <= Wgt_1_69;
		WeightsStore1[70] <= Wgt_1_70;
		WeightsStore1[71] <= Wgt_1_71;
		WeightsStore1[72] <= Wgt_1_72;
		WeightsStore1[73] <= Wgt_1_73;
		WeightsStore1[74] <= Wgt_1_74;
		WeightsStore1[75] <= Wgt_1_75;
		WeightsStore1[76] <= Wgt_1_76;
		WeightsStore1[77] <= Wgt_1_77;
		WeightsStore1[78] <= Wgt_1_78;
		WeightsStore1[79] <= Wgt_1_79;
		WeightsStore1[80] <= Wgt_1_80;
		WeightsStore1[81] <= Wgt_1_81;
		WeightsStore1[82] <= Wgt_1_82;
		WeightsStore1[83] <= Wgt_1_83;
		WeightsStore1[84] <= Wgt_1_84;
		WeightsStore1[85] <= Wgt_1_85;
		WeightsStore1[86] <= Wgt_1_86;
		WeightsStore1[87] <= Wgt_1_87;
		WeightsStore1[88] <= Wgt_1_88;
		WeightsStore1[89] <= Wgt_1_89;
		WeightsStore1[90] <= Wgt_1_90;
		WeightsStore1[91] <= Wgt_1_91;
		WeightsStore1[92] <= Wgt_1_92;
		WeightsStore1[93] <= Wgt_1_93;
		WeightsStore1[94] <= Wgt_1_94;
		WeightsStore1[95] <= Wgt_1_95;
		WeightsStore1[96] <= Wgt_1_96;
		WeightsStore1[97] <= Wgt_1_97;
		WeightsStore1[98] <= Wgt_1_98;
		WeightsStore1[99] <= Wgt_1_99;
		WeightsStore1[100] <= Wgt_1_100;
		WeightsStore1[101] <= Wgt_1_101;
		WeightsStore1[102] <= Wgt_1_102;
		WeightsStore1[103] <= Wgt_1_103;
		WeightsStore1[104] <= Wgt_1_104;
		WeightsStore1[105] <= Wgt_1_105;
		WeightsStore1[106] <= Wgt_1_106;
		WeightsStore1[107] <= Wgt_1_107;
		WeightsStore1[108] <= Wgt_1_108;
		WeightsStore1[109] <= Wgt_1_109;
		WeightsStore1[110] <= Wgt_1_110;
		WeightsStore1[111] <= Wgt_1_111;
		WeightsStore1[112] <= Wgt_1_112;
		WeightsStore1[113] <= Wgt_1_113;
		WeightsStore1[114] <= Wgt_1_114;
		WeightsStore1[115] <= Wgt_1_115;
		WeightsStore1[116] <= Wgt_1_116;
		WeightsStore1[117] <= Wgt_1_117;
		WeightsStore1[118] <= Wgt_1_118;
		WeightsStore1[119] <= Wgt_1_119;
		WeightsStore1[120] <= Wgt_1_120;
		WeightsStore1[121] <= Wgt_1_121;
		WeightsStore1[122] <= Wgt_1_122;
		WeightsStore1[123] <= Wgt_1_123;
		WeightsStore1[124] <= Wgt_1_124;
		WeightsStore1[125] <= Wgt_1_125;
		WeightsStore1[126] <= Wgt_1_126;
		WeightsStore1[127] <= Wgt_1_127;
		WeightsStore1[128] <= Wgt_1_128;
		WeightsStore1[129] <= Wgt_1_129;
		WeightsStore1[130] <= Wgt_1_130;
		WeightsStore1[131] <= Wgt_1_131;
		WeightsStore1[132] <= Wgt_1_132;
		WeightsStore1[133] <= Wgt_1_133;
		WeightsStore1[134] <= Wgt_1_134;
		WeightsStore1[135] <= Wgt_1_135;
		WeightsStore1[136] <= Wgt_1_136;
		WeightsStore1[137] <= Wgt_1_137;
		WeightsStore1[138] <= Wgt_1_138;
		WeightsStore1[139] <= Wgt_1_139;
		WeightsStore1[140] <= Wgt_1_140;
		WeightsStore1[141] <= Wgt_1_141;
		WeightsStore1[142] <= Wgt_1_142;
		WeightsStore1[143] <= Wgt_1_143;
		WeightsStore1[144] <= Wgt_1_144;
		WeightsStore1[145] <= Wgt_1_145;
		WeightsStore1[146] <= Wgt_1_146;
		WeightsStore1[147] <= Wgt_1_147;
		WeightsStore1[148] <= Wgt_1_148;
		WeightsStore1[149] <= Wgt_1_149;
		WeightsStore1[150] <= Wgt_1_150;
		WeightsStore1[151] <= Wgt_1_151;
		WeightsStore1[152] <= Wgt_1_152;
		WeightsStore1[153] <= Wgt_1_153;
		WeightsStore1[154] <= Wgt_1_154;
		WeightsStore1[155] <= Wgt_1_155;
		WeightsStore1[156] <= Wgt_1_156;
		WeightsStore1[157] <= Wgt_1_157;
		WeightsStore1[158] <= Wgt_1_158;
		WeightsStore1[159] <= Wgt_1_159;
		WeightsStore1[160] <= Wgt_1_160;
		WeightsStore1[161] <= Wgt_1_161;
		WeightsStore1[162] <= Wgt_1_162;
		WeightsStore1[163] <= Wgt_1_163;
		WeightsStore1[164] <= Wgt_1_164;
		WeightsStore1[165] <= Wgt_1_165;
		WeightsStore1[166] <= Wgt_1_166;
		WeightsStore1[167] <= Wgt_1_167;
		WeightsStore1[168] <= Wgt_1_168;
		WeightsStore1[169] <= Wgt_1_169;
		WeightsStore1[170] <= Wgt_1_170;
		WeightsStore1[171] <= Wgt_1_171;
		WeightsStore1[172] <= Wgt_1_172;
		WeightsStore1[173] <= Wgt_1_173;
		WeightsStore1[174] <= Wgt_1_174;
		WeightsStore1[175] <= Wgt_1_175;
		WeightsStore1[176] <= Wgt_1_176;
		WeightsStore1[177] <= Wgt_1_177;
		WeightsStore1[178] <= Wgt_1_178;
		WeightsStore1[179] <= Wgt_1_179;
		WeightsStore1[180] <= Wgt_1_180;
		WeightsStore1[181] <= Wgt_1_181;
		WeightsStore1[182] <= Wgt_1_182;
		WeightsStore1[183] <= Wgt_1_183;
		WeightsStore1[184] <= Wgt_1_184;
		WeightsStore1[185] <= Wgt_1_185;
		WeightsStore1[186] <= Wgt_1_186;
		WeightsStore1[187] <= Wgt_1_187;
		WeightsStore1[188] <= Wgt_1_188;
		WeightsStore1[189] <= Wgt_1_189;
		WeightsStore1[190] <= Wgt_1_190;
		WeightsStore1[191] <= Wgt_1_191;
		WeightsStore1[192] <= Wgt_1_192;
		WeightsStore1[193] <= Wgt_1_193;
		WeightsStore1[194] <= Wgt_1_194;
		WeightsStore1[195] <= Wgt_1_195;
		WeightsStore1[196] <= Wgt_1_196;
		WeightsStore1[197] <= Wgt_1_197;
		WeightsStore1[198] <= Wgt_1_198;
		WeightsStore1[199] <= Wgt_1_199;
		WeightsStore1[200] <= Wgt_1_200;
		WeightsStore1[201] <= Wgt_1_201;
		WeightsStore1[202] <= Wgt_1_202;
		WeightsStore1[203] <= Wgt_1_203;
		WeightsStore1[204] <= Wgt_1_204;
		WeightsStore1[205] <= Wgt_1_205;
		WeightsStore1[206] <= Wgt_1_206;
		WeightsStore1[207] <= Wgt_1_207;
		WeightsStore1[208] <= Wgt_1_208;
		WeightsStore1[209] <= Wgt_1_209;
		WeightsStore1[210] <= Wgt_1_210;
		WeightsStore1[211] <= Wgt_1_211;
		WeightsStore1[212] <= Wgt_1_212;
		WeightsStore1[213] <= Wgt_1_213;
		WeightsStore1[214] <= Wgt_1_214;
		WeightsStore1[215] <= Wgt_1_215;
		WeightsStore1[216] <= Wgt_1_216;
		WeightsStore1[217] <= Wgt_1_217;
		WeightsStore1[218] <= Wgt_1_218;
		WeightsStore1[219] <= Wgt_1_219;
		WeightsStore1[220] <= Wgt_1_220;
		WeightsStore1[221] <= Wgt_1_221;
		WeightsStore1[222] <= Wgt_1_222;
		WeightsStore1[223] <= Wgt_1_223;
		WeightsStore1[224] <= Wgt_1_224;
		WeightsStore1[225] <= Wgt_1_225;
		WeightsStore1[226] <= Wgt_1_226;
		WeightsStore1[227] <= Wgt_1_227;
		WeightsStore1[228] <= Wgt_1_228;
		WeightsStore1[229] <= Wgt_1_229;
		WeightsStore1[230] <= Wgt_1_230;
		WeightsStore1[231] <= Wgt_1_231;
		WeightsStore1[232] <= Wgt_1_232;
		WeightsStore1[233] <= Wgt_1_233;
		WeightsStore1[234] <= Wgt_1_234;
		WeightsStore1[235] <= Wgt_1_235;
		WeightsStore1[236] <= Wgt_1_236;
		WeightsStore1[237] <= Wgt_1_237;
		WeightsStore1[238] <= Wgt_1_238;
		WeightsStore1[239] <= Wgt_1_239;
		WeightsStore1[240] <= Wgt_1_240;
		WeightsStore1[241] <= Wgt_1_241;
		WeightsStore1[242] <= Wgt_1_242;
		WeightsStore1[243] <= Wgt_1_243;
		WeightsStore1[244] <= Wgt_1_244;
		WeightsStore1[245] <= Wgt_1_245;
		WeightsStore1[246] <= Wgt_1_246;
		WeightsStore1[247] <= Wgt_1_247;
		WeightsStore1[248] <= Wgt_1_248;
		WeightsStore1[249] <= Wgt_1_249;
		WeightsStore1[250] <= Wgt_1_250;
		WeightsStore1[251] <= Wgt_1_251;
		WeightsStore1[252] <= Wgt_1_252;
		WeightsStore1[253] <= Wgt_1_253;
		WeightsStore1[254] <= Wgt_1_254;
		WeightsStore1[255] <= Wgt_1_255;
		WeightsStore1[256] <= Wgt_1_256;
		WeightsStore1[257] <= Wgt_1_257;
		WeightsStore1[258] <= Wgt_1_258;
		WeightsStore1[259] <= Wgt_1_259;
		WeightsStore1[260] <= Wgt_1_260;
		WeightsStore1[261] <= Wgt_1_261;
		WeightsStore1[262] <= Wgt_1_262;
		WeightsStore1[263] <= Wgt_1_263;
		WeightsStore1[264] <= Wgt_1_264;
		WeightsStore1[265] <= Wgt_1_265;
		WeightsStore1[266] <= Wgt_1_266;
		WeightsStore1[267] <= Wgt_1_267;
		WeightsStore1[268] <= Wgt_1_268;
		WeightsStore1[269] <= Wgt_1_269;
		WeightsStore1[270] <= Wgt_1_270;
		WeightsStore1[271] <= Wgt_1_271;
		WeightsStore1[272] <= Wgt_1_272;
		WeightsStore1[273] <= Wgt_1_273;
		WeightsStore1[274] <= Wgt_1_274;
		WeightsStore1[275] <= Wgt_1_275;
		WeightsStore1[276] <= Wgt_1_276;
		WeightsStore1[277] <= Wgt_1_277;
		WeightsStore1[278] <= Wgt_1_278;
		WeightsStore1[279] <= Wgt_1_279;
		WeightsStore1[280] <= Wgt_1_280;
		WeightsStore1[281] <= Wgt_1_281;
		WeightsStore1[282] <= Wgt_1_282;
		WeightsStore1[283] <= Wgt_1_283;
		WeightsStore1[284] <= Wgt_1_284;
		WeightsStore1[285] <= Wgt_1_285;
		WeightsStore1[286] <= Wgt_1_286;
		WeightsStore1[287] <= Wgt_1_287;
		WeightsStore1[288] <= Wgt_1_288;
		WeightsStore1[289] <= Wgt_1_289;
		WeightsStore1[290] <= Wgt_1_290;
		WeightsStore1[291] <= Wgt_1_291;
		WeightsStore1[292] <= Wgt_1_292;
		WeightsStore1[293] <= Wgt_1_293;
		WeightsStore1[294] <= Wgt_1_294;
		WeightsStore1[295] <= Wgt_1_295;
		WeightsStore1[296] <= Wgt_1_296;
		WeightsStore1[297] <= Wgt_1_297;
		WeightsStore1[298] <= Wgt_1_298;
		WeightsStore1[299] <= Wgt_1_299;
		WeightsStore1[300] <= Wgt_1_300;
		WeightsStore1[301] <= Wgt_1_301;
		WeightsStore1[302] <= Wgt_1_302;
		WeightsStore1[303] <= Wgt_1_303;
		WeightsStore1[304] <= Wgt_1_304;
		WeightsStore1[305] <= Wgt_1_305;
		WeightsStore1[306] <= Wgt_1_306;
		WeightsStore1[307] <= Wgt_1_307;
		WeightsStore1[308] <= Wgt_1_308;
		WeightsStore1[309] <= Wgt_1_309;
		WeightsStore1[310] <= Wgt_1_310;
		WeightsStore1[311] <= Wgt_1_311;
		WeightsStore1[312] <= Wgt_1_312;
		WeightsStore1[313] <= Wgt_1_313;
		WeightsStore1[314] <= Wgt_1_314;
		WeightsStore1[315] <= Wgt_1_315;
		WeightsStore1[316] <= Wgt_1_316;
		WeightsStore1[317] <= Wgt_1_317;
		WeightsStore1[318] <= Wgt_1_318;
		WeightsStore1[319] <= Wgt_1_319;
		WeightsStore1[320] <= Wgt_1_320;
		WeightsStore1[321] <= Wgt_1_321;
		WeightsStore1[322] <= Wgt_1_322;
		WeightsStore1[323] <= Wgt_1_323;
		WeightsStore1[324] <= Wgt_1_324;
		WeightsStore1[325] <= Wgt_1_325;
		WeightsStore1[326] <= Wgt_1_326;
		WeightsStore1[327] <= Wgt_1_327;
		WeightsStore1[328] <= Wgt_1_328;
		WeightsStore1[329] <= Wgt_1_329;
		WeightsStore1[330] <= Wgt_1_330;
		WeightsStore1[331] <= Wgt_1_331;
		WeightsStore1[332] <= Wgt_1_332;
		WeightsStore1[333] <= Wgt_1_333;
		WeightsStore1[334] <= Wgt_1_334;
		WeightsStore1[335] <= Wgt_1_335;
		WeightsStore1[336] <= Wgt_1_336;
		WeightsStore1[337] <= Wgt_1_337;
		WeightsStore1[338] <= Wgt_1_338;
		WeightsStore1[339] <= Wgt_1_339;
		WeightsStore1[340] <= Wgt_1_340;
		WeightsStore1[341] <= Wgt_1_341;
		WeightsStore1[342] <= Wgt_1_342;
		WeightsStore1[343] <= Wgt_1_343;
		WeightsStore1[344] <= Wgt_1_344;
		WeightsStore1[345] <= Wgt_1_345;
		WeightsStore1[346] <= Wgt_1_346;
		WeightsStore1[347] <= Wgt_1_347;
		WeightsStore1[348] <= Wgt_1_348;
		WeightsStore1[349] <= Wgt_1_349;
		WeightsStore1[350] <= Wgt_1_350;
		WeightsStore1[351] <= Wgt_1_351;
		WeightsStore1[352] <= Wgt_1_352;
		WeightsStore1[353] <= Wgt_1_353;
		WeightsStore1[354] <= Wgt_1_354;
		WeightsStore1[355] <= Wgt_1_355;
		WeightsStore1[356] <= Wgt_1_356;
		WeightsStore1[357] <= Wgt_1_357;
		WeightsStore1[358] <= Wgt_1_358;
		WeightsStore1[359] <= Wgt_1_359;
		WeightsStore1[360] <= Wgt_1_360;
		WeightsStore1[361] <= Wgt_1_361;
		WeightsStore1[362] <= Wgt_1_362;
		WeightsStore1[363] <= Wgt_1_363;
		WeightsStore1[364] <= Wgt_1_364;
		WeightsStore1[365] <= Wgt_1_365;
		WeightsStore1[366] <= Wgt_1_366;
		WeightsStore1[367] <= Wgt_1_367;
		WeightsStore1[368] <= Wgt_1_368;
		WeightsStore1[369] <= Wgt_1_369;
		WeightsStore1[370] <= Wgt_1_370;
		WeightsStore1[371] <= Wgt_1_371;
		WeightsStore1[372] <= Wgt_1_372;
		WeightsStore1[373] <= Wgt_1_373;
		WeightsStore1[374] <= Wgt_1_374;
		WeightsStore1[375] <= Wgt_1_375;
		WeightsStore1[376] <= Wgt_1_376;
		WeightsStore1[377] <= Wgt_1_377;
		WeightsStore1[378] <= Wgt_1_378;
		WeightsStore1[379] <= Wgt_1_379;
		WeightsStore1[380] <= Wgt_1_380;
		WeightsStore1[381] <= Wgt_1_381;
		WeightsStore1[382] <= Wgt_1_382;
		WeightsStore1[383] <= Wgt_1_383;
		WeightsStore1[384] <= Wgt_1_384;
		WeightsStore1[385] <= Wgt_1_385;
		WeightsStore1[386] <= Wgt_1_386;
		WeightsStore1[387] <= Wgt_1_387;
		WeightsStore1[388] <= Wgt_1_388;
		WeightsStore1[389] <= Wgt_1_389;
		WeightsStore1[390] <= Wgt_1_390;
		WeightsStore1[391] <= Wgt_1_391;
		WeightsStore1[392] <= Wgt_1_392;
		WeightsStore1[393] <= Wgt_1_393;
		WeightsStore1[394] <= Wgt_1_394;
		WeightsStore1[395] <= Wgt_1_395;
		WeightsStore1[396] <= Wgt_1_396;
		WeightsStore1[397] <= Wgt_1_397;
		WeightsStore1[398] <= Wgt_1_398;
		WeightsStore1[399] <= Wgt_1_399;
		WeightsStore1[400] <= Wgt_1_400;
		WeightsStore1[401] <= Wgt_1_401;
		WeightsStore1[402] <= Wgt_1_402;
		WeightsStore1[403] <= Wgt_1_403;
		WeightsStore1[404] <= Wgt_1_404;
		WeightsStore1[405] <= Wgt_1_405;
		WeightsStore1[406] <= Wgt_1_406;
		WeightsStore1[407] <= Wgt_1_407;
		WeightsStore1[408] <= Wgt_1_408;
		WeightsStore1[409] <= Wgt_1_409;
		WeightsStore1[410] <= Wgt_1_410;
		WeightsStore1[411] <= Wgt_1_411;
		WeightsStore1[412] <= Wgt_1_412;
		WeightsStore1[413] <= Wgt_1_413;
		WeightsStore1[414] <= Wgt_1_414;
		WeightsStore1[415] <= Wgt_1_415;
		WeightsStore1[416] <= Wgt_1_416;
		WeightsStore1[417] <= Wgt_1_417;
		WeightsStore1[418] <= Wgt_1_418;
		WeightsStore1[419] <= Wgt_1_419;
		WeightsStore1[420] <= Wgt_1_420;
		WeightsStore1[421] <= Wgt_1_421;
		WeightsStore1[422] <= Wgt_1_422;
		WeightsStore1[423] <= Wgt_1_423;
		WeightsStore1[424] <= Wgt_1_424;
		WeightsStore1[425] <= Wgt_1_425;
		WeightsStore1[426] <= Wgt_1_426;
		WeightsStore1[427] <= Wgt_1_427;
		WeightsStore1[428] <= Wgt_1_428;
		WeightsStore1[429] <= Wgt_1_429;
		WeightsStore1[430] <= Wgt_1_430;
		WeightsStore1[431] <= Wgt_1_431;
		WeightsStore1[432] <= Wgt_1_432;
		WeightsStore1[433] <= Wgt_1_433;
		WeightsStore1[434] <= Wgt_1_434;
		WeightsStore1[435] <= Wgt_1_435;
		WeightsStore1[436] <= Wgt_1_436;
		WeightsStore1[437] <= Wgt_1_437;
		WeightsStore1[438] <= Wgt_1_438;
		WeightsStore1[439] <= Wgt_1_439;
		WeightsStore1[440] <= Wgt_1_440;
		WeightsStore1[441] <= Wgt_1_441;
		WeightsStore1[442] <= Wgt_1_442;
		WeightsStore1[443] <= Wgt_1_443;
		WeightsStore1[444] <= Wgt_1_444;
		WeightsStore1[445] <= Wgt_1_445;
		WeightsStore1[446] <= Wgt_1_446;
		WeightsStore1[447] <= Wgt_1_447;
		WeightsStore1[448] <= Wgt_1_448;
		WeightsStore1[449] <= Wgt_1_449;
		WeightsStore1[450] <= Wgt_1_450;
		WeightsStore1[451] <= Wgt_1_451;
		WeightsStore1[452] <= Wgt_1_452;
		WeightsStore1[453] <= Wgt_1_453;
		WeightsStore1[454] <= Wgt_1_454;
		WeightsStore1[455] <= Wgt_1_455;
		WeightsStore1[456] <= Wgt_1_456;
		WeightsStore1[457] <= Wgt_1_457;
		WeightsStore1[458] <= Wgt_1_458;
		WeightsStore1[459] <= Wgt_1_459;
		WeightsStore1[460] <= Wgt_1_460;
		WeightsStore1[461] <= Wgt_1_461;
		WeightsStore1[462] <= Wgt_1_462;
		WeightsStore1[463] <= Wgt_1_463;
		WeightsStore1[464] <= Wgt_1_464;
		WeightsStore1[465] <= Wgt_1_465;
		WeightsStore1[466] <= Wgt_1_466;
		WeightsStore1[467] <= Wgt_1_467;
		WeightsStore1[468] <= Wgt_1_468;
		WeightsStore1[469] <= Wgt_1_469;
		WeightsStore1[470] <= Wgt_1_470;
		WeightsStore1[471] <= Wgt_1_471;
		WeightsStore1[472] <= Wgt_1_472;
		WeightsStore1[473] <= Wgt_1_473;
		WeightsStore1[474] <= Wgt_1_474;
		WeightsStore1[475] <= Wgt_1_475;
		WeightsStore1[476] <= Wgt_1_476;
		WeightsStore1[477] <= Wgt_1_477;
		WeightsStore1[478] <= Wgt_1_478;
		WeightsStore1[479] <= Wgt_1_479;
		WeightsStore1[480] <= Wgt_1_480;
		WeightsStore1[481] <= Wgt_1_481;
		WeightsStore1[482] <= Wgt_1_482;
		WeightsStore1[483] <= Wgt_1_483;
		WeightsStore1[484] <= Wgt_1_484;
		WeightsStore1[485] <= Wgt_1_485;
		WeightsStore1[486] <= Wgt_1_486;
		WeightsStore1[487] <= Wgt_1_487;
		WeightsStore1[488] <= Wgt_1_488;
		WeightsStore1[489] <= Wgt_1_489;
		WeightsStore1[490] <= Wgt_1_490;
		WeightsStore1[491] <= Wgt_1_491;
		WeightsStore1[492] <= Wgt_1_492;
		WeightsStore1[493] <= Wgt_1_493;
		WeightsStore1[494] <= Wgt_1_494;
		WeightsStore1[495] <= Wgt_1_495;
		WeightsStore1[496] <= Wgt_1_496;
		WeightsStore1[497] <= Wgt_1_497;
		WeightsStore1[498] <= Wgt_1_498;
		WeightsStore1[499] <= Wgt_1_499;
		WeightsStore1[500] <= Wgt_1_500;
		WeightsStore1[501] <= Wgt_1_501;
		WeightsStore1[502] <= Wgt_1_502;
		WeightsStore1[503] <= Wgt_1_503;
		WeightsStore1[504] <= Wgt_1_504;
		WeightsStore1[505] <= Wgt_1_505;
		WeightsStore1[506] <= Wgt_1_506;
		WeightsStore1[507] <= Wgt_1_507;
		WeightsStore1[508] <= Wgt_1_508;
		WeightsStore1[509] <= Wgt_1_509;
		WeightsStore1[510] <= Wgt_1_510;
		WeightsStore1[511] <= Wgt_1_511;
		WeightsStore1[512] <= Wgt_1_512;
		WeightsStore1[513] <= Wgt_1_513;
		WeightsStore1[514] <= Wgt_1_514;
		WeightsStore1[515] <= Wgt_1_515;
		WeightsStore1[516] <= Wgt_1_516;
		WeightsStore1[517] <= Wgt_1_517;
		WeightsStore1[518] <= Wgt_1_518;
		WeightsStore1[519] <= Wgt_1_519;
		WeightsStore1[520] <= Wgt_1_520;
		WeightsStore1[521] <= Wgt_1_521;
		WeightsStore1[522] <= Wgt_1_522;
		WeightsStore1[523] <= Wgt_1_523;
		WeightsStore1[524] <= Wgt_1_524;
		WeightsStore1[525] <= Wgt_1_525;
		WeightsStore1[526] <= Wgt_1_526;
		WeightsStore1[527] <= Wgt_1_527;
		WeightsStore1[528] <= Wgt_1_528;
		WeightsStore1[529] <= Wgt_1_529;
		WeightsStore1[530] <= Wgt_1_530;
		WeightsStore1[531] <= Wgt_1_531;
		WeightsStore1[532] <= Wgt_1_532;
		WeightsStore1[533] <= Wgt_1_533;
		WeightsStore1[534] <= Wgt_1_534;
		WeightsStore1[535] <= Wgt_1_535;
		WeightsStore1[536] <= Wgt_1_536;
		WeightsStore1[537] <= Wgt_1_537;
		WeightsStore1[538] <= Wgt_1_538;
		WeightsStore1[539] <= Wgt_1_539;
		WeightsStore1[540] <= Wgt_1_540;
		WeightsStore1[541] <= Wgt_1_541;
		WeightsStore1[542] <= Wgt_1_542;
		WeightsStore1[543] <= Wgt_1_543;
		WeightsStore1[544] <= Wgt_1_544;
		WeightsStore1[545] <= Wgt_1_545;
		WeightsStore1[546] <= Wgt_1_546;
		WeightsStore1[547] <= Wgt_1_547;
		WeightsStore1[548] <= Wgt_1_548;
		WeightsStore1[549] <= Wgt_1_549;
		WeightsStore1[550] <= Wgt_1_550;
		WeightsStore1[551] <= Wgt_1_551;
		WeightsStore1[552] <= Wgt_1_552;
		WeightsStore1[553] <= Wgt_1_553;
		WeightsStore1[554] <= Wgt_1_554;
		WeightsStore1[555] <= Wgt_1_555;
		WeightsStore1[556] <= Wgt_1_556;
		WeightsStore1[557] <= Wgt_1_557;
		WeightsStore1[558] <= Wgt_1_558;
		WeightsStore1[559] <= Wgt_1_559;
		WeightsStore1[560] <= Wgt_1_560;
		WeightsStore1[561] <= Wgt_1_561;
		WeightsStore1[562] <= Wgt_1_562;
		WeightsStore1[563] <= Wgt_1_563;
		WeightsStore1[564] <= Wgt_1_564;
		WeightsStore1[565] <= Wgt_1_565;
		WeightsStore1[566] <= Wgt_1_566;
		WeightsStore1[567] <= Wgt_1_567;
		WeightsStore1[568] <= Wgt_1_568;
		WeightsStore1[569] <= Wgt_1_569;
		WeightsStore1[570] <= Wgt_1_570;
		WeightsStore1[571] <= Wgt_1_571;
		WeightsStore1[572] <= Wgt_1_572;
		WeightsStore1[573] <= Wgt_1_573;
		WeightsStore1[574] <= Wgt_1_574;
		WeightsStore1[575] <= Wgt_1_575;
		WeightsStore1[576] <= Wgt_1_576;
		WeightsStore1[577] <= Wgt_1_577;
		WeightsStore1[578] <= Wgt_1_578;
		WeightsStore1[579] <= Wgt_1_579;
		WeightsStore1[580] <= Wgt_1_580;
		WeightsStore1[581] <= Wgt_1_581;
		WeightsStore1[582] <= Wgt_1_582;
		WeightsStore1[583] <= Wgt_1_583;
		WeightsStore1[584] <= Wgt_1_584;
		WeightsStore1[585] <= Wgt_1_585;
		WeightsStore1[586] <= Wgt_1_586;
		WeightsStore1[587] <= Wgt_1_587;
		WeightsStore1[588] <= Wgt_1_588;
		WeightsStore1[589] <= Wgt_1_589;
		WeightsStore1[590] <= Wgt_1_590;
		WeightsStore1[591] <= Wgt_1_591;
		WeightsStore1[592] <= Wgt_1_592;
		WeightsStore1[593] <= Wgt_1_593;
		WeightsStore1[594] <= Wgt_1_594;
		WeightsStore1[595] <= Wgt_1_595;
		WeightsStore1[596] <= Wgt_1_596;
		WeightsStore1[597] <= Wgt_1_597;
		WeightsStore1[598] <= Wgt_1_598;
		WeightsStore1[599] <= Wgt_1_599;
		WeightsStore1[600] <= Wgt_1_600;
		WeightsStore1[601] <= Wgt_1_601;
		WeightsStore1[602] <= Wgt_1_602;
		WeightsStore1[603] <= Wgt_1_603;
		WeightsStore1[604] <= Wgt_1_604;
		WeightsStore1[605] <= Wgt_1_605;
		WeightsStore1[606] <= Wgt_1_606;
		WeightsStore1[607] <= Wgt_1_607;
		WeightsStore1[608] <= Wgt_1_608;
		WeightsStore1[609] <= Wgt_1_609;
		WeightsStore1[610] <= Wgt_1_610;
		WeightsStore1[611] <= Wgt_1_611;
		WeightsStore1[612] <= Wgt_1_612;
		WeightsStore1[613] <= Wgt_1_613;
		WeightsStore1[614] <= Wgt_1_614;
		WeightsStore1[615] <= Wgt_1_615;
		WeightsStore1[616] <= Wgt_1_616;
		WeightsStore1[617] <= Wgt_1_617;
		WeightsStore1[618] <= Wgt_1_618;
		WeightsStore1[619] <= Wgt_1_619;
		WeightsStore1[620] <= Wgt_1_620;
		WeightsStore1[621] <= Wgt_1_621;
		WeightsStore1[622] <= Wgt_1_622;
		WeightsStore1[623] <= Wgt_1_623;
		WeightsStore1[624] <= Wgt_1_624;
		WeightsStore1[625] <= Wgt_1_625;
		WeightsStore1[626] <= Wgt_1_626;
		WeightsStore1[627] <= Wgt_1_627;
		WeightsStore1[628] <= Wgt_1_628;
		WeightsStore1[629] <= Wgt_1_629;
		WeightsStore1[630] <= Wgt_1_630;
		WeightsStore1[631] <= Wgt_1_631;
		WeightsStore1[632] <= Wgt_1_632;
		WeightsStore1[633] <= Wgt_1_633;
		WeightsStore1[634] <= Wgt_1_634;
		WeightsStore1[635] <= Wgt_1_635;
		WeightsStore1[636] <= Wgt_1_636;
		WeightsStore1[637] <= Wgt_1_637;
		WeightsStore1[638] <= Wgt_1_638;
		WeightsStore1[639] <= Wgt_1_639;
		WeightsStore1[640] <= Wgt_1_640;
		WeightsStore1[641] <= Wgt_1_641;
		WeightsStore1[642] <= Wgt_1_642;
		WeightsStore1[643] <= Wgt_1_643;
		WeightsStore1[644] <= Wgt_1_644;
		WeightsStore1[645] <= Wgt_1_645;
		WeightsStore1[646] <= Wgt_1_646;
		WeightsStore1[647] <= Wgt_1_647;
		WeightsStore1[648] <= Wgt_1_648;
		WeightsStore1[649] <= Wgt_1_649;
		WeightsStore1[650] <= Wgt_1_650;
		WeightsStore1[651] <= Wgt_1_651;
		WeightsStore1[652] <= Wgt_1_652;
		WeightsStore1[653] <= Wgt_1_653;
		WeightsStore1[654] <= Wgt_1_654;
		WeightsStore1[655] <= Wgt_1_655;
		WeightsStore1[656] <= Wgt_1_656;
		WeightsStore1[657] <= Wgt_1_657;
		WeightsStore1[658] <= Wgt_1_658;
		WeightsStore1[659] <= Wgt_1_659;
		WeightsStore1[660] <= Wgt_1_660;
		WeightsStore1[661] <= Wgt_1_661;
		WeightsStore1[662] <= Wgt_1_662;
		WeightsStore1[663] <= Wgt_1_663;
		WeightsStore1[664] <= Wgt_1_664;
		WeightsStore1[665] <= Wgt_1_665;
		WeightsStore1[666] <= Wgt_1_666;
		WeightsStore1[667] <= Wgt_1_667;
		WeightsStore1[668] <= Wgt_1_668;
		WeightsStore1[669] <= Wgt_1_669;
		WeightsStore1[670] <= Wgt_1_670;
		WeightsStore1[671] <= Wgt_1_671;
		WeightsStore1[672] <= Wgt_1_672;
		WeightsStore1[673] <= Wgt_1_673;
		WeightsStore1[674] <= Wgt_1_674;
		WeightsStore1[675] <= Wgt_1_675;
		WeightsStore1[676] <= Wgt_1_676;
		WeightsStore1[677] <= Wgt_1_677;
		WeightsStore1[678] <= Wgt_1_678;
		WeightsStore1[679] <= Wgt_1_679;
		WeightsStore1[680] <= Wgt_1_680;
		WeightsStore1[681] <= Wgt_1_681;
		WeightsStore1[682] <= Wgt_1_682;
		WeightsStore1[683] <= Wgt_1_683;
		WeightsStore1[684] <= Wgt_1_684;
		WeightsStore1[685] <= Wgt_1_685;
		WeightsStore1[686] <= Wgt_1_686;
		WeightsStore1[687] <= Wgt_1_687;
		WeightsStore1[688] <= Wgt_1_688;
		WeightsStore1[689] <= Wgt_1_689;
		WeightsStore1[690] <= Wgt_1_690;
		WeightsStore1[691] <= Wgt_1_691;
		WeightsStore1[692] <= Wgt_1_692;
		WeightsStore1[693] <= Wgt_1_693;
		WeightsStore1[694] <= Wgt_1_694;
		WeightsStore1[695] <= Wgt_1_695;
		WeightsStore1[696] <= Wgt_1_696;
		WeightsStore1[697] <= Wgt_1_697;
		WeightsStore1[698] <= Wgt_1_698;
		WeightsStore1[699] <= Wgt_1_699;
		WeightsStore1[700] <= Wgt_1_700;
		WeightsStore1[701] <= Wgt_1_701;
		WeightsStore1[702] <= Wgt_1_702;
		WeightsStore1[703] <= Wgt_1_703;
		WeightsStore1[704] <= Wgt_1_704;
		WeightsStore1[705] <= Wgt_1_705;
		WeightsStore1[706] <= Wgt_1_706;
		WeightsStore1[707] <= Wgt_1_707;
		WeightsStore1[708] <= Wgt_1_708;
		WeightsStore1[709] <= Wgt_1_709;
		WeightsStore1[710] <= Wgt_1_710;
		WeightsStore1[711] <= Wgt_1_711;
		WeightsStore1[712] <= Wgt_1_712;
		WeightsStore1[713] <= Wgt_1_713;
		WeightsStore1[714] <= Wgt_1_714;
		WeightsStore1[715] <= Wgt_1_715;
		WeightsStore1[716] <= Wgt_1_716;
		WeightsStore1[717] <= Wgt_1_717;
		WeightsStore1[718] <= Wgt_1_718;
		WeightsStore1[719] <= Wgt_1_719;
		WeightsStore1[720] <= Wgt_1_720;
		WeightsStore1[721] <= Wgt_1_721;
		WeightsStore1[722] <= Wgt_1_722;
		WeightsStore1[723] <= Wgt_1_723;
		WeightsStore1[724] <= Wgt_1_724;
		WeightsStore1[725] <= Wgt_1_725;
		WeightsStore1[726] <= Wgt_1_726;
		WeightsStore1[727] <= Wgt_1_727;
		WeightsStore1[728] <= Wgt_1_728;
		WeightsStore1[729] <= Wgt_1_729;
		WeightsStore1[730] <= Wgt_1_730;
		WeightsStore1[731] <= Wgt_1_731;
		WeightsStore1[732] <= Wgt_1_732;
		WeightsStore1[733] <= Wgt_1_733;
		WeightsStore1[734] <= Wgt_1_734;
		WeightsStore1[735] <= Wgt_1_735;
		WeightsStore1[736] <= Wgt_1_736;
		WeightsStore1[737] <= Wgt_1_737;
		WeightsStore1[738] <= Wgt_1_738;
		WeightsStore1[739] <= Wgt_1_739;
		WeightsStore1[740] <= Wgt_1_740;
		WeightsStore1[741] <= Wgt_1_741;
		WeightsStore1[742] <= Wgt_1_742;
		WeightsStore1[743] <= Wgt_1_743;
		WeightsStore1[744] <= Wgt_1_744;
		WeightsStore1[745] <= Wgt_1_745;
		WeightsStore1[746] <= Wgt_1_746;
		WeightsStore1[747] <= Wgt_1_747;
		WeightsStore1[748] <= Wgt_1_748;
		WeightsStore1[749] <= Wgt_1_749;
		WeightsStore1[750] <= Wgt_1_750;
		WeightsStore1[751] <= Wgt_1_751;
		WeightsStore1[752] <= Wgt_1_752;
		WeightsStore1[753] <= Wgt_1_753;
		WeightsStore1[754] <= Wgt_1_754;
		WeightsStore1[755] <= Wgt_1_755;
		WeightsStore1[756] <= Wgt_1_756;
		WeightsStore1[757] <= Wgt_1_757;
		WeightsStore1[758] <= Wgt_1_758;
		WeightsStore1[759] <= Wgt_1_759;
		WeightsStore1[760] <= Wgt_1_760;
		WeightsStore1[761] <= Wgt_1_761;
		WeightsStore1[762] <= Wgt_1_762;
		WeightsStore1[763] <= Wgt_1_763;
		WeightsStore1[764] <= Wgt_1_764;
		WeightsStore1[765] <= Wgt_1_765;
		WeightsStore1[766] <= Wgt_1_766;
		WeightsStore1[767] <= Wgt_1_767;
		WeightsStore1[768] <= Wgt_1_768;
		WeightsStore1[769] <= Wgt_1_769;
		WeightsStore1[770] <= Wgt_1_770;
		WeightsStore1[771] <= Wgt_1_771;
		WeightsStore1[772] <= Wgt_1_772;
		WeightsStore1[773] <= Wgt_1_773;
		WeightsStore1[774] <= Wgt_1_774;
		WeightsStore1[775] <= Wgt_1_775;
		WeightsStore1[776] <= Wgt_1_776;
		WeightsStore1[777] <= Wgt_1_777;
		WeightsStore1[778] <= Wgt_1_778;
		WeightsStore1[779] <= Wgt_1_779;
		WeightsStore1[780] <= Wgt_1_780;
		WeightsStore1[781] <= Wgt_1_781;
		WeightsStore1[782] <= Wgt_1_782;
		WeightsStore1[783] <= Wgt_1_783;
		WeightsStore1[784] <= Wgt_1_784;
		WeightsStore2[0] <= Wgt_2_0;
		WeightsStore2[1] <= Wgt_2_1;
		WeightsStore2[2] <= Wgt_2_2;
		WeightsStore2[3] <= Wgt_2_3;
		WeightsStore2[4] <= Wgt_2_4;
		WeightsStore2[5] <= Wgt_2_5;
		WeightsStore2[6] <= Wgt_2_6;
		WeightsStore2[7] <= Wgt_2_7;
		WeightsStore2[8] <= Wgt_2_8;
		WeightsStore2[9] <= Wgt_2_9;
		WeightsStore2[10] <= Wgt_2_10;
		WeightsStore2[11] <= Wgt_2_11;
		WeightsStore2[12] <= Wgt_2_12;
		WeightsStore2[13] <= Wgt_2_13;
		WeightsStore2[14] <= Wgt_2_14;
		WeightsStore2[15] <= Wgt_2_15;
		WeightsStore2[16] <= Wgt_2_16;
		WeightsStore2[17] <= Wgt_2_17;
		WeightsStore2[18] <= Wgt_2_18;
		WeightsStore2[19] <= Wgt_2_19;
		WeightsStore2[20] <= Wgt_2_20;
		WeightsStore2[21] <= Wgt_2_21;
		WeightsStore2[22] <= Wgt_2_22;
		WeightsStore2[23] <= Wgt_2_23;
		WeightsStore2[24] <= Wgt_2_24;
		WeightsStore2[25] <= Wgt_2_25;
		WeightsStore2[26] <= Wgt_2_26;
		WeightsStore2[27] <= Wgt_2_27;
		WeightsStore2[28] <= Wgt_2_28;
		WeightsStore2[29] <= Wgt_2_29;
		WeightsStore2[30] <= Wgt_2_30;
		WeightsStore2[31] <= Wgt_2_31;
		WeightsStore2[32] <= Wgt_2_32;
		WeightsStore2[33] <= Wgt_2_33;
		WeightsStore2[34] <= Wgt_2_34;
		WeightsStore2[35] <= Wgt_2_35;
		WeightsStore2[36] <= Wgt_2_36;
		WeightsStore2[37] <= Wgt_2_37;
		WeightsStore2[38] <= Wgt_2_38;
		WeightsStore2[39] <= Wgt_2_39;
		WeightsStore2[40] <= Wgt_2_40;
		WeightsStore2[41] <= Wgt_2_41;
		WeightsStore2[42] <= Wgt_2_42;
		WeightsStore2[43] <= Wgt_2_43;
		WeightsStore2[44] <= Wgt_2_44;
		WeightsStore2[45] <= Wgt_2_45;
		WeightsStore2[46] <= Wgt_2_46;
		WeightsStore2[47] <= Wgt_2_47;
		WeightsStore2[48] <= Wgt_2_48;
		WeightsStore2[49] <= Wgt_2_49;
		WeightsStore2[50] <= Wgt_2_50;
		WeightsStore2[51] <= Wgt_2_51;
		WeightsStore2[52] <= Wgt_2_52;
		WeightsStore2[53] <= Wgt_2_53;
		WeightsStore2[54] <= Wgt_2_54;
		WeightsStore2[55] <= Wgt_2_55;
		WeightsStore2[56] <= Wgt_2_56;
		WeightsStore2[57] <= Wgt_2_57;
		WeightsStore2[58] <= Wgt_2_58;
		WeightsStore2[59] <= Wgt_2_59;
		WeightsStore2[60] <= Wgt_2_60;
		WeightsStore2[61] <= Wgt_2_61;
		WeightsStore2[62] <= Wgt_2_62;
		WeightsStore2[63] <= Wgt_2_63;
		WeightsStore2[64] <= Wgt_2_64;
		WeightsStore2[65] <= Wgt_2_65;
		WeightsStore2[66] <= Wgt_2_66;
		WeightsStore2[67] <= Wgt_2_67;
		WeightsStore2[68] <= Wgt_2_68;
		WeightsStore2[69] <= Wgt_2_69;
		WeightsStore2[70] <= Wgt_2_70;
		WeightsStore2[71] <= Wgt_2_71;
		WeightsStore2[72] <= Wgt_2_72;
		WeightsStore2[73] <= Wgt_2_73;
		WeightsStore2[74] <= Wgt_2_74;
		WeightsStore2[75] <= Wgt_2_75;
		WeightsStore2[76] <= Wgt_2_76;
		WeightsStore2[77] <= Wgt_2_77;
		WeightsStore2[78] <= Wgt_2_78;
		WeightsStore2[79] <= Wgt_2_79;
		WeightsStore2[80] <= Wgt_2_80;
		WeightsStore2[81] <= Wgt_2_81;
		WeightsStore2[82] <= Wgt_2_82;
		WeightsStore2[83] <= Wgt_2_83;
		WeightsStore2[84] <= Wgt_2_84;
		WeightsStore2[85] <= Wgt_2_85;
		WeightsStore2[86] <= Wgt_2_86;
		WeightsStore2[87] <= Wgt_2_87;
		WeightsStore2[88] <= Wgt_2_88;
		WeightsStore2[89] <= Wgt_2_89;
		WeightsStore2[90] <= Wgt_2_90;
		WeightsStore2[91] <= Wgt_2_91;
		WeightsStore2[92] <= Wgt_2_92;
		WeightsStore2[93] <= Wgt_2_93;
		WeightsStore2[94] <= Wgt_2_94;
		WeightsStore2[95] <= Wgt_2_95;
		WeightsStore2[96] <= Wgt_2_96;
		WeightsStore2[97] <= Wgt_2_97;
		WeightsStore2[98] <= Wgt_2_98;
		WeightsStore2[99] <= Wgt_2_99;
		WeightsStore2[100] <= Wgt_2_100;
		WeightsStore2[101] <= Wgt_2_101;
		WeightsStore2[102] <= Wgt_2_102;
		WeightsStore2[103] <= Wgt_2_103;
		WeightsStore2[104] <= Wgt_2_104;
		WeightsStore2[105] <= Wgt_2_105;
		WeightsStore2[106] <= Wgt_2_106;
		WeightsStore2[107] <= Wgt_2_107;
		WeightsStore2[108] <= Wgt_2_108;
		WeightsStore2[109] <= Wgt_2_109;
		WeightsStore2[110] <= Wgt_2_110;
		WeightsStore2[111] <= Wgt_2_111;
		WeightsStore2[112] <= Wgt_2_112;
		WeightsStore2[113] <= Wgt_2_113;
		WeightsStore2[114] <= Wgt_2_114;
		WeightsStore2[115] <= Wgt_2_115;
		WeightsStore2[116] <= Wgt_2_116;
		WeightsStore2[117] <= Wgt_2_117;
		WeightsStore2[118] <= Wgt_2_118;
		WeightsStore2[119] <= Wgt_2_119;
		WeightsStore2[120] <= Wgt_2_120;
		WeightsStore2[121] <= Wgt_2_121;
		WeightsStore2[122] <= Wgt_2_122;
		WeightsStore2[123] <= Wgt_2_123;
		WeightsStore2[124] <= Wgt_2_124;
		WeightsStore2[125] <= Wgt_2_125;
		WeightsStore2[126] <= Wgt_2_126;
		WeightsStore2[127] <= Wgt_2_127;
		WeightsStore2[128] <= Wgt_2_128;
		WeightsStore2[129] <= Wgt_2_129;
		WeightsStore2[130] <= Wgt_2_130;
		WeightsStore2[131] <= Wgt_2_131;
		WeightsStore2[132] <= Wgt_2_132;
		WeightsStore2[133] <= Wgt_2_133;
		WeightsStore2[134] <= Wgt_2_134;
		WeightsStore2[135] <= Wgt_2_135;
		WeightsStore2[136] <= Wgt_2_136;
		WeightsStore2[137] <= Wgt_2_137;
		WeightsStore2[138] <= Wgt_2_138;
		WeightsStore2[139] <= Wgt_2_139;
		WeightsStore2[140] <= Wgt_2_140;
		WeightsStore2[141] <= Wgt_2_141;
		WeightsStore2[142] <= Wgt_2_142;
		WeightsStore2[143] <= Wgt_2_143;
		WeightsStore2[144] <= Wgt_2_144;
		WeightsStore2[145] <= Wgt_2_145;
		WeightsStore2[146] <= Wgt_2_146;
		WeightsStore2[147] <= Wgt_2_147;
		WeightsStore2[148] <= Wgt_2_148;
		WeightsStore2[149] <= Wgt_2_149;
		WeightsStore2[150] <= Wgt_2_150;
		WeightsStore2[151] <= Wgt_2_151;
		WeightsStore2[152] <= Wgt_2_152;
		WeightsStore2[153] <= Wgt_2_153;
		WeightsStore2[154] <= Wgt_2_154;
		WeightsStore2[155] <= Wgt_2_155;
		WeightsStore2[156] <= Wgt_2_156;
		WeightsStore2[157] <= Wgt_2_157;
		WeightsStore2[158] <= Wgt_2_158;
		WeightsStore2[159] <= Wgt_2_159;
		WeightsStore2[160] <= Wgt_2_160;
		WeightsStore2[161] <= Wgt_2_161;
		WeightsStore2[162] <= Wgt_2_162;
		WeightsStore2[163] <= Wgt_2_163;
		WeightsStore2[164] <= Wgt_2_164;
		WeightsStore2[165] <= Wgt_2_165;
		WeightsStore2[166] <= Wgt_2_166;
		WeightsStore2[167] <= Wgt_2_167;
		WeightsStore2[168] <= Wgt_2_168;
		WeightsStore2[169] <= Wgt_2_169;
		WeightsStore2[170] <= Wgt_2_170;
		WeightsStore2[171] <= Wgt_2_171;
		WeightsStore2[172] <= Wgt_2_172;
		WeightsStore2[173] <= Wgt_2_173;
		WeightsStore2[174] <= Wgt_2_174;
		WeightsStore2[175] <= Wgt_2_175;
		WeightsStore2[176] <= Wgt_2_176;
		WeightsStore2[177] <= Wgt_2_177;
		WeightsStore2[178] <= Wgt_2_178;
		WeightsStore2[179] <= Wgt_2_179;
		WeightsStore2[180] <= Wgt_2_180;
		WeightsStore2[181] <= Wgt_2_181;
		WeightsStore2[182] <= Wgt_2_182;
		WeightsStore2[183] <= Wgt_2_183;
		WeightsStore2[184] <= Wgt_2_184;
		WeightsStore2[185] <= Wgt_2_185;
		WeightsStore2[186] <= Wgt_2_186;
		WeightsStore2[187] <= Wgt_2_187;
		WeightsStore2[188] <= Wgt_2_188;
		WeightsStore2[189] <= Wgt_2_189;
		WeightsStore2[190] <= Wgt_2_190;
		WeightsStore2[191] <= Wgt_2_191;
		WeightsStore2[192] <= Wgt_2_192;
		WeightsStore2[193] <= Wgt_2_193;
		WeightsStore2[194] <= Wgt_2_194;
		WeightsStore2[195] <= Wgt_2_195;
		WeightsStore2[196] <= Wgt_2_196;
		WeightsStore2[197] <= Wgt_2_197;
		WeightsStore2[198] <= Wgt_2_198;
		WeightsStore2[199] <= Wgt_2_199;
		WeightsStore2[200] <= Wgt_2_200;
		WeightsStore2[201] <= Wgt_2_201;
		WeightsStore2[202] <= Wgt_2_202;
		WeightsStore2[203] <= Wgt_2_203;
		WeightsStore2[204] <= Wgt_2_204;
		WeightsStore2[205] <= Wgt_2_205;
		WeightsStore2[206] <= Wgt_2_206;
		WeightsStore2[207] <= Wgt_2_207;
		WeightsStore2[208] <= Wgt_2_208;
		WeightsStore2[209] <= Wgt_2_209;
		WeightsStore2[210] <= Wgt_2_210;
		WeightsStore2[211] <= Wgt_2_211;
		WeightsStore2[212] <= Wgt_2_212;
		WeightsStore2[213] <= Wgt_2_213;
		WeightsStore2[214] <= Wgt_2_214;
		WeightsStore2[215] <= Wgt_2_215;
		WeightsStore2[216] <= Wgt_2_216;
		WeightsStore2[217] <= Wgt_2_217;
		WeightsStore2[218] <= Wgt_2_218;
		WeightsStore2[219] <= Wgt_2_219;
		WeightsStore2[220] <= Wgt_2_220;
		WeightsStore2[221] <= Wgt_2_221;
		WeightsStore2[222] <= Wgt_2_222;
		WeightsStore2[223] <= Wgt_2_223;
		WeightsStore2[224] <= Wgt_2_224;
		WeightsStore2[225] <= Wgt_2_225;
		WeightsStore2[226] <= Wgt_2_226;
		WeightsStore2[227] <= Wgt_2_227;
		WeightsStore2[228] <= Wgt_2_228;
		WeightsStore2[229] <= Wgt_2_229;
		WeightsStore2[230] <= Wgt_2_230;
		WeightsStore2[231] <= Wgt_2_231;
		WeightsStore2[232] <= Wgt_2_232;
		WeightsStore2[233] <= Wgt_2_233;
		WeightsStore2[234] <= Wgt_2_234;
		WeightsStore2[235] <= Wgt_2_235;
		WeightsStore2[236] <= Wgt_2_236;
		WeightsStore2[237] <= Wgt_2_237;
		WeightsStore2[238] <= Wgt_2_238;
		WeightsStore2[239] <= Wgt_2_239;
		WeightsStore2[240] <= Wgt_2_240;
		WeightsStore2[241] <= Wgt_2_241;
		WeightsStore2[242] <= Wgt_2_242;
		WeightsStore2[243] <= Wgt_2_243;
		WeightsStore2[244] <= Wgt_2_244;
		WeightsStore2[245] <= Wgt_2_245;
		WeightsStore2[246] <= Wgt_2_246;
		WeightsStore2[247] <= Wgt_2_247;
		WeightsStore2[248] <= Wgt_2_248;
		WeightsStore2[249] <= Wgt_2_249;
		WeightsStore2[250] <= Wgt_2_250;
		WeightsStore2[251] <= Wgt_2_251;
		WeightsStore2[252] <= Wgt_2_252;
		WeightsStore2[253] <= Wgt_2_253;
		WeightsStore2[254] <= Wgt_2_254;
		WeightsStore2[255] <= Wgt_2_255;
		WeightsStore2[256] <= Wgt_2_256;
		WeightsStore2[257] <= Wgt_2_257;
		WeightsStore2[258] <= Wgt_2_258;
		WeightsStore2[259] <= Wgt_2_259;
		WeightsStore2[260] <= Wgt_2_260;
		WeightsStore2[261] <= Wgt_2_261;
		WeightsStore2[262] <= Wgt_2_262;
		WeightsStore2[263] <= Wgt_2_263;
		WeightsStore2[264] <= Wgt_2_264;
		WeightsStore2[265] <= Wgt_2_265;
		WeightsStore2[266] <= Wgt_2_266;
		WeightsStore2[267] <= Wgt_2_267;
		WeightsStore2[268] <= Wgt_2_268;
		WeightsStore2[269] <= Wgt_2_269;
		WeightsStore2[270] <= Wgt_2_270;
		WeightsStore2[271] <= Wgt_2_271;
		WeightsStore2[272] <= Wgt_2_272;
		WeightsStore2[273] <= Wgt_2_273;
		WeightsStore2[274] <= Wgt_2_274;
		WeightsStore2[275] <= Wgt_2_275;
		WeightsStore2[276] <= Wgt_2_276;
		WeightsStore2[277] <= Wgt_2_277;
		WeightsStore2[278] <= Wgt_2_278;
		WeightsStore2[279] <= Wgt_2_279;
		WeightsStore2[280] <= Wgt_2_280;
		WeightsStore2[281] <= Wgt_2_281;
		WeightsStore2[282] <= Wgt_2_282;
		WeightsStore2[283] <= Wgt_2_283;
		WeightsStore2[284] <= Wgt_2_284;
		WeightsStore2[285] <= Wgt_2_285;
		WeightsStore2[286] <= Wgt_2_286;
		WeightsStore2[287] <= Wgt_2_287;
		WeightsStore2[288] <= Wgt_2_288;
		WeightsStore2[289] <= Wgt_2_289;
		WeightsStore2[290] <= Wgt_2_290;
		WeightsStore2[291] <= Wgt_2_291;
		WeightsStore2[292] <= Wgt_2_292;
		WeightsStore2[293] <= Wgt_2_293;
		WeightsStore2[294] <= Wgt_2_294;
		WeightsStore2[295] <= Wgt_2_295;
		WeightsStore2[296] <= Wgt_2_296;
		WeightsStore2[297] <= Wgt_2_297;
		WeightsStore2[298] <= Wgt_2_298;
		WeightsStore2[299] <= Wgt_2_299;
		WeightsStore2[300] <= Wgt_2_300;
		WeightsStore2[301] <= Wgt_2_301;
		WeightsStore2[302] <= Wgt_2_302;
		WeightsStore2[303] <= Wgt_2_303;
		WeightsStore2[304] <= Wgt_2_304;
		WeightsStore2[305] <= Wgt_2_305;
		WeightsStore2[306] <= Wgt_2_306;
		WeightsStore2[307] <= Wgt_2_307;
		WeightsStore2[308] <= Wgt_2_308;
		WeightsStore2[309] <= Wgt_2_309;
		WeightsStore2[310] <= Wgt_2_310;
		WeightsStore2[311] <= Wgt_2_311;
		WeightsStore2[312] <= Wgt_2_312;
		WeightsStore2[313] <= Wgt_2_313;
		WeightsStore2[314] <= Wgt_2_314;
		WeightsStore2[315] <= Wgt_2_315;
		WeightsStore2[316] <= Wgt_2_316;
		WeightsStore2[317] <= Wgt_2_317;
		WeightsStore2[318] <= Wgt_2_318;
		WeightsStore2[319] <= Wgt_2_319;
		WeightsStore2[320] <= Wgt_2_320;
		WeightsStore2[321] <= Wgt_2_321;
		WeightsStore2[322] <= Wgt_2_322;
		WeightsStore2[323] <= Wgt_2_323;
		WeightsStore2[324] <= Wgt_2_324;
		WeightsStore2[325] <= Wgt_2_325;
		WeightsStore2[326] <= Wgt_2_326;
		WeightsStore2[327] <= Wgt_2_327;
		WeightsStore2[328] <= Wgt_2_328;
		WeightsStore2[329] <= Wgt_2_329;
		WeightsStore2[330] <= Wgt_2_330;
		WeightsStore2[331] <= Wgt_2_331;
		WeightsStore2[332] <= Wgt_2_332;
		WeightsStore2[333] <= Wgt_2_333;
		WeightsStore2[334] <= Wgt_2_334;
		WeightsStore2[335] <= Wgt_2_335;
		WeightsStore2[336] <= Wgt_2_336;
		WeightsStore2[337] <= Wgt_2_337;
		WeightsStore2[338] <= Wgt_2_338;
		WeightsStore2[339] <= Wgt_2_339;
		WeightsStore2[340] <= Wgt_2_340;
		WeightsStore2[341] <= Wgt_2_341;
		WeightsStore2[342] <= Wgt_2_342;
		WeightsStore2[343] <= Wgt_2_343;
		WeightsStore2[344] <= Wgt_2_344;
		WeightsStore2[345] <= Wgt_2_345;
		WeightsStore2[346] <= Wgt_2_346;
		WeightsStore2[347] <= Wgt_2_347;
		WeightsStore2[348] <= Wgt_2_348;
		WeightsStore2[349] <= Wgt_2_349;
		WeightsStore2[350] <= Wgt_2_350;
		WeightsStore2[351] <= Wgt_2_351;
		WeightsStore2[352] <= Wgt_2_352;
		WeightsStore2[353] <= Wgt_2_353;
		WeightsStore2[354] <= Wgt_2_354;
		WeightsStore2[355] <= Wgt_2_355;
		WeightsStore2[356] <= Wgt_2_356;
		WeightsStore2[357] <= Wgt_2_357;
		WeightsStore2[358] <= Wgt_2_358;
		WeightsStore2[359] <= Wgt_2_359;
		WeightsStore2[360] <= Wgt_2_360;
		WeightsStore2[361] <= Wgt_2_361;
		WeightsStore2[362] <= Wgt_2_362;
		WeightsStore2[363] <= Wgt_2_363;
		WeightsStore2[364] <= Wgt_2_364;
		WeightsStore2[365] <= Wgt_2_365;
		WeightsStore2[366] <= Wgt_2_366;
		WeightsStore2[367] <= Wgt_2_367;
		WeightsStore2[368] <= Wgt_2_368;
		WeightsStore2[369] <= Wgt_2_369;
		WeightsStore2[370] <= Wgt_2_370;
		WeightsStore2[371] <= Wgt_2_371;
		WeightsStore2[372] <= Wgt_2_372;
		WeightsStore2[373] <= Wgt_2_373;
		WeightsStore2[374] <= Wgt_2_374;
		WeightsStore2[375] <= Wgt_2_375;
		WeightsStore2[376] <= Wgt_2_376;
		WeightsStore2[377] <= Wgt_2_377;
		WeightsStore2[378] <= Wgt_2_378;
		WeightsStore2[379] <= Wgt_2_379;
		WeightsStore2[380] <= Wgt_2_380;
		WeightsStore2[381] <= Wgt_2_381;
		WeightsStore2[382] <= Wgt_2_382;
		WeightsStore2[383] <= Wgt_2_383;
		WeightsStore2[384] <= Wgt_2_384;
		WeightsStore2[385] <= Wgt_2_385;
		WeightsStore2[386] <= Wgt_2_386;
		WeightsStore2[387] <= Wgt_2_387;
		WeightsStore2[388] <= Wgt_2_388;
		WeightsStore2[389] <= Wgt_2_389;
		WeightsStore2[390] <= Wgt_2_390;
		WeightsStore2[391] <= Wgt_2_391;
		WeightsStore2[392] <= Wgt_2_392;
		WeightsStore2[393] <= Wgt_2_393;
		WeightsStore2[394] <= Wgt_2_394;
		WeightsStore2[395] <= Wgt_2_395;
		WeightsStore2[396] <= Wgt_2_396;
		WeightsStore2[397] <= Wgt_2_397;
		WeightsStore2[398] <= Wgt_2_398;
		WeightsStore2[399] <= Wgt_2_399;
		WeightsStore2[400] <= Wgt_2_400;
		WeightsStore2[401] <= Wgt_2_401;
		WeightsStore2[402] <= Wgt_2_402;
		WeightsStore2[403] <= Wgt_2_403;
		WeightsStore2[404] <= Wgt_2_404;
		WeightsStore2[405] <= Wgt_2_405;
		WeightsStore2[406] <= Wgt_2_406;
		WeightsStore2[407] <= Wgt_2_407;
		WeightsStore2[408] <= Wgt_2_408;
		WeightsStore2[409] <= Wgt_2_409;
		WeightsStore2[410] <= Wgt_2_410;
		WeightsStore2[411] <= Wgt_2_411;
		WeightsStore2[412] <= Wgt_2_412;
		WeightsStore2[413] <= Wgt_2_413;
		WeightsStore2[414] <= Wgt_2_414;
		WeightsStore2[415] <= Wgt_2_415;
		WeightsStore2[416] <= Wgt_2_416;
		WeightsStore2[417] <= Wgt_2_417;
		WeightsStore2[418] <= Wgt_2_418;
		WeightsStore2[419] <= Wgt_2_419;
		WeightsStore2[420] <= Wgt_2_420;
		WeightsStore2[421] <= Wgt_2_421;
		WeightsStore2[422] <= Wgt_2_422;
		WeightsStore2[423] <= Wgt_2_423;
		WeightsStore2[424] <= Wgt_2_424;
		WeightsStore2[425] <= Wgt_2_425;
		WeightsStore2[426] <= Wgt_2_426;
		WeightsStore2[427] <= Wgt_2_427;
		WeightsStore2[428] <= Wgt_2_428;
		WeightsStore2[429] <= Wgt_2_429;
		WeightsStore2[430] <= Wgt_2_430;
		WeightsStore2[431] <= Wgt_2_431;
		WeightsStore2[432] <= Wgt_2_432;
		WeightsStore2[433] <= Wgt_2_433;
		WeightsStore2[434] <= Wgt_2_434;
		WeightsStore2[435] <= Wgt_2_435;
		WeightsStore2[436] <= Wgt_2_436;
		WeightsStore2[437] <= Wgt_2_437;
		WeightsStore2[438] <= Wgt_2_438;
		WeightsStore2[439] <= Wgt_2_439;
		WeightsStore2[440] <= Wgt_2_440;
		WeightsStore2[441] <= Wgt_2_441;
		WeightsStore2[442] <= Wgt_2_442;
		WeightsStore2[443] <= Wgt_2_443;
		WeightsStore2[444] <= Wgt_2_444;
		WeightsStore2[445] <= Wgt_2_445;
		WeightsStore2[446] <= Wgt_2_446;
		WeightsStore2[447] <= Wgt_2_447;
		WeightsStore2[448] <= Wgt_2_448;
		WeightsStore2[449] <= Wgt_2_449;
		WeightsStore2[450] <= Wgt_2_450;
		WeightsStore2[451] <= Wgt_2_451;
		WeightsStore2[452] <= Wgt_2_452;
		WeightsStore2[453] <= Wgt_2_453;
		WeightsStore2[454] <= Wgt_2_454;
		WeightsStore2[455] <= Wgt_2_455;
		WeightsStore2[456] <= Wgt_2_456;
		WeightsStore2[457] <= Wgt_2_457;
		WeightsStore2[458] <= Wgt_2_458;
		WeightsStore2[459] <= Wgt_2_459;
		WeightsStore2[460] <= Wgt_2_460;
		WeightsStore2[461] <= Wgt_2_461;
		WeightsStore2[462] <= Wgt_2_462;
		WeightsStore2[463] <= Wgt_2_463;
		WeightsStore2[464] <= Wgt_2_464;
		WeightsStore2[465] <= Wgt_2_465;
		WeightsStore2[466] <= Wgt_2_466;
		WeightsStore2[467] <= Wgt_2_467;
		WeightsStore2[468] <= Wgt_2_468;
		WeightsStore2[469] <= Wgt_2_469;
		WeightsStore2[470] <= Wgt_2_470;
		WeightsStore2[471] <= Wgt_2_471;
		WeightsStore2[472] <= Wgt_2_472;
		WeightsStore2[473] <= Wgt_2_473;
		WeightsStore2[474] <= Wgt_2_474;
		WeightsStore2[475] <= Wgt_2_475;
		WeightsStore2[476] <= Wgt_2_476;
		WeightsStore2[477] <= Wgt_2_477;
		WeightsStore2[478] <= Wgt_2_478;
		WeightsStore2[479] <= Wgt_2_479;
		WeightsStore2[480] <= Wgt_2_480;
		WeightsStore2[481] <= Wgt_2_481;
		WeightsStore2[482] <= Wgt_2_482;
		WeightsStore2[483] <= Wgt_2_483;
		WeightsStore2[484] <= Wgt_2_484;
		WeightsStore2[485] <= Wgt_2_485;
		WeightsStore2[486] <= Wgt_2_486;
		WeightsStore2[487] <= Wgt_2_487;
		WeightsStore2[488] <= Wgt_2_488;
		WeightsStore2[489] <= Wgt_2_489;
		WeightsStore2[490] <= Wgt_2_490;
		WeightsStore2[491] <= Wgt_2_491;
		WeightsStore2[492] <= Wgt_2_492;
		WeightsStore2[493] <= Wgt_2_493;
		WeightsStore2[494] <= Wgt_2_494;
		WeightsStore2[495] <= Wgt_2_495;
		WeightsStore2[496] <= Wgt_2_496;
		WeightsStore2[497] <= Wgt_2_497;
		WeightsStore2[498] <= Wgt_2_498;
		WeightsStore2[499] <= Wgt_2_499;
		WeightsStore2[500] <= Wgt_2_500;
		WeightsStore2[501] <= Wgt_2_501;
		WeightsStore2[502] <= Wgt_2_502;
		WeightsStore2[503] <= Wgt_2_503;
		WeightsStore2[504] <= Wgt_2_504;
		WeightsStore2[505] <= Wgt_2_505;
		WeightsStore2[506] <= Wgt_2_506;
		WeightsStore2[507] <= Wgt_2_507;
		WeightsStore2[508] <= Wgt_2_508;
		WeightsStore2[509] <= Wgt_2_509;
		WeightsStore2[510] <= Wgt_2_510;
		WeightsStore2[511] <= Wgt_2_511;
		WeightsStore2[512] <= Wgt_2_512;
		WeightsStore2[513] <= Wgt_2_513;
		WeightsStore2[514] <= Wgt_2_514;
		WeightsStore2[515] <= Wgt_2_515;
		WeightsStore2[516] <= Wgt_2_516;
		WeightsStore2[517] <= Wgt_2_517;
		WeightsStore2[518] <= Wgt_2_518;
		WeightsStore2[519] <= Wgt_2_519;
		WeightsStore2[520] <= Wgt_2_520;
		WeightsStore2[521] <= Wgt_2_521;
		WeightsStore2[522] <= Wgt_2_522;
		WeightsStore2[523] <= Wgt_2_523;
		WeightsStore2[524] <= Wgt_2_524;
		WeightsStore2[525] <= Wgt_2_525;
		WeightsStore2[526] <= Wgt_2_526;
		WeightsStore2[527] <= Wgt_2_527;
		WeightsStore2[528] <= Wgt_2_528;
		WeightsStore2[529] <= Wgt_2_529;
		WeightsStore2[530] <= Wgt_2_530;
		WeightsStore2[531] <= Wgt_2_531;
		WeightsStore2[532] <= Wgt_2_532;
		WeightsStore2[533] <= Wgt_2_533;
		WeightsStore2[534] <= Wgt_2_534;
		WeightsStore2[535] <= Wgt_2_535;
		WeightsStore2[536] <= Wgt_2_536;
		WeightsStore2[537] <= Wgt_2_537;
		WeightsStore2[538] <= Wgt_2_538;
		WeightsStore2[539] <= Wgt_2_539;
		WeightsStore2[540] <= Wgt_2_540;
		WeightsStore2[541] <= Wgt_2_541;
		WeightsStore2[542] <= Wgt_2_542;
		WeightsStore2[543] <= Wgt_2_543;
		WeightsStore2[544] <= Wgt_2_544;
		WeightsStore2[545] <= Wgt_2_545;
		WeightsStore2[546] <= Wgt_2_546;
		WeightsStore2[547] <= Wgt_2_547;
		WeightsStore2[548] <= Wgt_2_548;
		WeightsStore2[549] <= Wgt_2_549;
		WeightsStore2[550] <= Wgt_2_550;
		WeightsStore2[551] <= Wgt_2_551;
		WeightsStore2[552] <= Wgt_2_552;
		WeightsStore2[553] <= Wgt_2_553;
		WeightsStore2[554] <= Wgt_2_554;
		WeightsStore2[555] <= Wgt_2_555;
		WeightsStore2[556] <= Wgt_2_556;
		WeightsStore2[557] <= Wgt_2_557;
		WeightsStore2[558] <= Wgt_2_558;
		WeightsStore2[559] <= Wgt_2_559;
		WeightsStore2[560] <= Wgt_2_560;
		WeightsStore2[561] <= Wgt_2_561;
		WeightsStore2[562] <= Wgt_2_562;
		WeightsStore2[563] <= Wgt_2_563;
		WeightsStore2[564] <= Wgt_2_564;
		WeightsStore2[565] <= Wgt_2_565;
		WeightsStore2[566] <= Wgt_2_566;
		WeightsStore2[567] <= Wgt_2_567;
		WeightsStore2[568] <= Wgt_2_568;
		WeightsStore2[569] <= Wgt_2_569;
		WeightsStore2[570] <= Wgt_2_570;
		WeightsStore2[571] <= Wgt_2_571;
		WeightsStore2[572] <= Wgt_2_572;
		WeightsStore2[573] <= Wgt_2_573;
		WeightsStore2[574] <= Wgt_2_574;
		WeightsStore2[575] <= Wgt_2_575;
		WeightsStore2[576] <= Wgt_2_576;
		WeightsStore2[577] <= Wgt_2_577;
		WeightsStore2[578] <= Wgt_2_578;
		WeightsStore2[579] <= Wgt_2_579;
		WeightsStore2[580] <= Wgt_2_580;
		WeightsStore2[581] <= Wgt_2_581;
		WeightsStore2[582] <= Wgt_2_582;
		WeightsStore2[583] <= Wgt_2_583;
		WeightsStore2[584] <= Wgt_2_584;
		WeightsStore2[585] <= Wgt_2_585;
		WeightsStore2[586] <= Wgt_2_586;
		WeightsStore2[587] <= Wgt_2_587;
		WeightsStore2[588] <= Wgt_2_588;
		WeightsStore2[589] <= Wgt_2_589;
		WeightsStore2[590] <= Wgt_2_590;
		WeightsStore2[591] <= Wgt_2_591;
		WeightsStore2[592] <= Wgt_2_592;
		WeightsStore2[593] <= Wgt_2_593;
		WeightsStore2[594] <= Wgt_2_594;
		WeightsStore2[595] <= Wgt_2_595;
		WeightsStore2[596] <= Wgt_2_596;
		WeightsStore2[597] <= Wgt_2_597;
		WeightsStore2[598] <= Wgt_2_598;
		WeightsStore2[599] <= Wgt_2_599;
		WeightsStore2[600] <= Wgt_2_600;
		WeightsStore2[601] <= Wgt_2_601;
		WeightsStore2[602] <= Wgt_2_602;
		WeightsStore2[603] <= Wgt_2_603;
		WeightsStore2[604] <= Wgt_2_604;
		WeightsStore2[605] <= Wgt_2_605;
		WeightsStore2[606] <= Wgt_2_606;
		WeightsStore2[607] <= Wgt_2_607;
		WeightsStore2[608] <= Wgt_2_608;
		WeightsStore2[609] <= Wgt_2_609;
		WeightsStore2[610] <= Wgt_2_610;
		WeightsStore2[611] <= Wgt_2_611;
		WeightsStore2[612] <= Wgt_2_612;
		WeightsStore2[613] <= Wgt_2_613;
		WeightsStore2[614] <= Wgt_2_614;
		WeightsStore2[615] <= Wgt_2_615;
		WeightsStore2[616] <= Wgt_2_616;
		WeightsStore2[617] <= Wgt_2_617;
		WeightsStore2[618] <= Wgt_2_618;
		WeightsStore2[619] <= Wgt_2_619;
		WeightsStore2[620] <= Wgt_2_620;
		WeightsStore2[621] <= Wgt_2_621;
		WeightsStore2[622] <= Wgt_2_622;
		WeightsStore2[623] <= Wgt_2_623;
		WeightsStore2[624] <= Wgt_2_624;
		WeightsStore2[625] <= Wgt_2_625;
		WeightsStore2[626] <= Wgt_2_626;
		WeightsStore2[627] <= Wgt_2_627;
		WeightsStore2[628] <= Wgt_2_628;
		WeightsStore2[629] <= Wgt_2_629;
		WeightsStore2[630] <= Wgt_2_630;
		WeightsStore2[631] <= Wgt_2_631;
		WeightsStore2[632] <= Wgt_2_632;
		WeightsStore2[633] <= Wgt_2_633;
		WeightsStore2[634] <= Wgt_2_634;
		WeightsStore2[635] <= Wgt_2_635;
		WeightsStore2[636] <= Wgt_2_636;
		WeightsStore2[637] <= Wgt_2_637;
		WeightsStore2[638] <= Wgt_2_638;
		WeightsStore2[639] <= Wgt_2_639;
		WeightsStore2[640] <= Wgt_2_640;
		WeightsStore2[641] <= Wgt_2_641;
		WeightsStore2[642] <= Wgt_2_642;
		WeightsStore2[643] <= Wgt_2_643;
		WeightsStore2[644] <= Wgt_2_644;
		WeightsStore2[645] <= Wgt_2_645;
		WeightsStore2[646] <= Wgt_2_646;
		WeightsStore2[647] <= Wgt_2_647;
		WeightsStore2[648] <= Wgt_2_648;
		WeightsStore2[649] <= Wgt_2_649;
		WeightsStore2[650] <= Wgt_2_650;
		WeightsStore2[651] <= Wgt_2_651;
		WeightsStore2[652] <= Wgt_2_652;
		WeightsStore2[653] <= Wgt_2_653;
		WeightsStore2[654] <= Wgt_2_654;
		WeightsStore2[655] <= Wgt_2_655;
		WeightsStore2[656] <= Wgt_2_656;
		WeightsStore2[657] <= Wgt_2_657;
		WeightsStore2[658] <= Wgt_2_658;
		WeightsStore2[659] <= Wgt_2_659;
		WeightsStore2[660] <= Wgt_2_660;
		WeightsStore2[661] <= Wgt_2_661;
		WeightsStore2[662] <= Wgt_2_662;
		WeightsStore2[663] <= Wgt_2_663;
		WeightsStore2[664] <= Wgt_2_664;
		WeightsStore2[665] <= Wgt_2_665;
		WeightsStore2[666] <= Wgt_2_666;
		WeightsStore2[667] <= Wgt_2_667;
		WeightsStore2[668] <= Wgt_2_668;
		WeightsStore2[669] <= Wgt_2_669;
		WeightsStore2[670] <= Wgt_2_670;
		WeightsStore2[671] <= Wgt_2_671;
		WeightsStore2[672] <= Wgt_2_672;
		WeightsStore2[673] <= Wgt_2_673;
		WeightsStore2[674] <= Wgt_2_674;
		WeightsStore2[675] <= Wgt_2_675;
		WeightsStore2[676] <= Wgt_2_676;
		WeightsStore2[677] <= Wgt_2_677;
		WeightsStore2[678] <= Wgt_2_678;
		WeightsStore2[679] <= Wgt_2_679;
		WeightsStore2[680] <= Wgt_2_680;
		WeightsStore2[681] <= Wgt_2_681;
		WeightsStore2[682] <= Wgt_2_682;
		WeightsStore2[683] <= Wgt_2_683;
		WeightsStore2[684] <= Wgt_2_684;
		WeightsStore2[685] <= Wgt_2_685;
		WeightsStore2[686] <= Wgt_2_686;
		WeightsStore2[687] <= Wgt_2_687;
		WeightsStore2[688] <= Wgt_2_688;
		WeightsStore2[689] <= Wgt_2_689;
		WeightsStore2[690] <= Wgt_2_690;
		WeightsStore2[691] <= Wgt_2_691;
		WeightsStore2[692] <= Wgt_2_692;
		WeightsStore2[693] <= Wgt_2_693;
		WeightsStore2[694] <= Wgt_2_694;
		WeightsStore2[695] <= Wgt_2_695;
		WeightsStore2[696] <= Wgt_2_696;
		WeightsStore2[697] <= Wgt_2_697;
		WeightsStore2[698] <= Wgt_2_698;
		WeightsStore2[699] <= Wgt_2_699;
		WeightsStore2[700] <= Wgt_2_700;
		WeightsStore2[701] <= Wgt_2_701;
		WeightsStore2[702] <= Wgt_2_702;
		WeightsStore2[703] <= Wgt_2_703;
		WeightsStore2[704] <= Wgt_2_704;
		WeightsStore2[705] <= Wgt_2_705;
		WeightsStore2[706] <= Wgt_2_706;
		WeightsStore2[707] <= Wgt_2_707;
		WeightsStore2[708] <= Wgt_2_708;
		WeightsStore2[709] <= Wgt_2_709;
		WeightsStore2[710] <= Wgt_2_710;
		WeightsStore2[711] <= Wgt_2_711;
		WeightsStore2[712] <= Wgt_2_712;
		WeightsStore2[713] <= Wgt_2_713;
		WeightsStore2[714] <= Wgt_2_714;
		WeightsStore2[715] <= Wgt_2_715;
		WeightsStore2[716] <= Wgt_2_716;
		WeightsStore2[717] <= Wgt_2_717;
		WeightsStore2[718] <= Wgt_2_718;
		WeightsStore2[719] <= Wgt_2_719;
		WeightsStore2[720] <= Wgt_2_720;
		WeightsStore2[721] <= Wgt_2_721;
		WeightsStore2[722] <= Wgt_2_722;
		WeightsStore2[723] <= Wgt_2_723;
		WeightsStore2[724] <= Wgt_2_724;
		WeightsStore2[725] <= Wgt_2_725;
		WeightsStore2[726] <= Wgt_2_726;
		WeightsStore2[727] <= Wgt_2_727;
		WeightsStore2[728] <= Wgt_2_728;
		WeightsStore2[729] <= Wgt_2_729;
		WeightsStore2[730] <= Wgt_2_730;
		WeightsStore2[731] <= Wgt_2_731;
		WeightsStore2[732] <= Wgt_2_732;
		WeightsStore2[733] <= Wgt_2_733;
		WeightsStore2[734] <= Wgt_2_734;
		WeightsStore2[735] <= Wgt_2_735;
		WeightsStore2[736] <= Wgt_2_736;
		WeightsStore2[737] <= Wgt_2_737;
		WeightsStore2[738] <= Wgt_2_738;
		WeightsStore2[739] <= Wgt_2_739;
		WeightsStore2[740] <= Wgt_2_740;
		WeightsStore2[741] <= Wgt_2_741;
		WeightsStore2[742] <= Wgt_2_742;
		WeightsStore2[743] <= Wgt_2_743;
		WeightsStore2[744] <= Wgt_2_744;
		WeightsStore2[745] <= Wgt_2_745;
		WeightsStore2[746] <= Wgt_2_746;
		WeightsStore2[747] <= Wgt_2_747;
		WeightsStore2[748] <= Wgt_2_748;
		WeightsStore2[749] <= Wgt_2_749;
		WeightsStore2[750] <= Wgt_2_750;
		WeightsStore2[751] <= Wgt_2_751;
		WeightsStore2[752] <= Wgt_2_752;
		WeightsStore2[753] <= Wgt_2_753;
		WeightsStore2[754] <= Wgt_2_754;
		WeightsStore2[755] <= Wgt_2_755;
		WeightsStore2[756] <= Wgt_2_756;
		WeightsStore2[757] <= Wgt_2_757;
		WeightsStore2[758] <= Wgt_2_758;
		WeightsStore2[759] <= Wgt_2_759;
		WeightsStore2[760] <= Wgt_2_760;
		WeightsStore2[761] <= Wgt_2_761;
		WeightsStore2[762] <= Wgt_2_762;
		WeightsStore2[763] <= Wgt_2_763;
		WeightsStore2[764] <= Wgt_2_764;
		WeightsStore2[765] <= Wgt_2_765;
		WeightsStore2[766] <= Wgt_2_766;
		WeightsStore2[767] <= Wgt_2_767;
		WeightsStore2[768] <= Wgt_2_768;
		WeightsStore2[769] <= Wgt_2_769;
		WeightsStore2[770] <= Wgt_2_770;
		WeightsStore2[771] <= Wgt_2_771;
		WeightsStore2[772] <= Wgt_2_772;
		WeightsStore2[773] <= Wgt_2_773;
		WeightsStore2[774] <= Wgt_2_774;
		WeightsStore2[775] <= Wgt_2_775;
		WeightsStore2[776] <= Wgt_2_776;
		WeightsStore2[777] <= Wgt_2_777;
		WeightsStore2[778] <= Wgt_2_778;
		WeightsStore2[779] <= Wgt_2_779;
		WeightsStore2[780] <= Wgt_2_780;
		WeightsStore2[781] <= Wgt_2_781;
		WeightsStore2[782] <= Wgt_2_782;
		WeightsStore2[783] <= Wgt_2_783;
		WeightsStore2[784] <= Wgt_2_784;
		WeightsStore3[0] <= Wgt_3_0;
		WeightsStore3[1] <= Wgt_3_1;
		WeightsStore3[2] <= Wgt_3_2;
		WeightsStore3[3] <= Wgt_3_3;
		WeightsStore3[4] <= Wgt_3_4;
		WeightsStore3[5] <= Wgt_3_5;
		WeightsStore3[6] <= Wgt_3_6;
		WeightsStore3[7] <= Wgt_3_7;
		WeightsStore3[8] <= Wgt_3_8;
		WeightsStore3[9] <= Wgt_3_9;
		WeightsStore3[10] <= Wgt_3_10;
		WeightsStore3[11] <= Wgt_3_11;
		WeightsStore3[12] <= Wgt_3_12;
		WeightsStore3[13] <= Wgt_3_13;
		WeightsStore3[14] <= Wgt_3_14;
		WeightsStore3[15] <= Wgt_3_15;
		WeightsStore3[16] <= Wgt_3_16;
		WeightsStore3[17] <= Wgt_3_17;
		WeightsStore3[18] <= Wgt_3_18;
		WeightsStore3[19] <= Wgt_3_19;
		WeightsStore3[20] <= Wgt_3_20;
		WeightsStore3[21] <= Wgt_3_21;
		WeightsStore3[22] <= Wgt_3_22;
		WeightsStore3[23] <= Wgt_3_23;
		WeightsStore3[24] <= Wgt_3_24;
		WeightsStore3[25] <= Wgt_3_25;
		WeightsStore3[26] <= Wgt_3_26;
		WeightsStore3[27] <= Wgt_3_27;
		WeightsStore3[28] <= Wgt_3_28;
		WeightsStore3[29] <= Wgt_3_29;
		WeightsStore3[30] <= Wgt_3_30;
		WeightsStore3[31] <= Wgt_3_31;
		WeightsStore3[32] <= Wgt_3_32;
		WeightsStore3[33] <= Wgt_3_33;
		WeightsStore3[34] <= Wgt_3_34;
		WeightsStore3[35] <= Wgt_3_35;
		WeightsStore3[36] <= Wgt_3_36;
		WeightsStore3[37] <= Wgt_3_37;
		WeightsStore3[38] <= Wgt_3_38;
		WeightsStore3[39] <= Wgt_3_39;
		WeightsStore3[40] <= Wgt_3_40;
		WeightsStore3[41] <= Wgt_3_41;
		WeightsStore3[42] <= Wgt_3_42;
		WeightsStore3[43] <= Wgt_3_43;
		WeightsStore3[44] <= Wgt_3_44;
		WeightsStore3[45] <= Wgt_3_45;
		WeightsStore3[46] <= Wgt_3_46;
		WeightsStore3[47] <= Wgt_3_47;
		WeightsStore3[48] <= Wgt_3_48;
		WeightsStore3[49] <= Wgt_3_49;
		WeightsStore3[50] <= Wgt_3_50;
		WeightsStore3[51] <= Wgt_3_51;
		WeightsStore3[52] <= Wgt_3_52;
		WeightsStore3[53] <= Wgt_3_53;
		WeightsStore3[54] <= Wgt_3_54;
		WeightsStore3[55] <= Wgt_3_55;
		WeightsStore3[56] <= Wgt_3_56;
		WeightsStore3[57] <= Wgt_3_57;
		WeightsStore3[58] <= Wgt_3_58;
		WeightsStore3[59] <= Wgt_3_59;
		WeightsStore3[60] <= Wgt_3_60;
		WeightsStore3[61] <= Wgt_3_61;
		WeightsStore3[62] <= Wgt_3_62;
		WeightsStore3[63] <= Wgt_3_63;
		WeightsStore3[64] <= Wgt_3_64;
		WeightsStore3[65] <= Wgt_3_65;
		WeightsStore3[66] <= Wgt_3_66;
		WeightsStore3[67] <= Wgt_3_67;
		WeightsStore3[68] <= Wgt_3_68;
		WeightsStore3[69] <= Wgt_3_69;
		WeightsStore3[70] <= Wgt_3_70;
		WeightsStore3[71] <= Wgt_3_71;
		WeightsStore3[72] <= Wgt_3_72;
		WeightsStore3[73] <= Wgt_3_73;
		WeightsStore3[74] <= Wgt_3_74;
		WeightsStore3[75] <= Wgt_3_75;
		WeightsStore3[76] <= Wgt_3_76;
		WeightsStore3[77] <= Wgt_3_77;
		WeightsStore3[78] <= Wgt_3_78;
		WeightsStore3[79] <= Wgt_3_79;
		WeightsStore3[80] <= Wgt_3_80;
		WeightsStore3[81] <= Wgt_3_81;
		WeightsStore3[82] <= Wgt_3_82;
		WeightsStore3[83] <= Wgt_3_83;
		WeightsStore3[84] <= Wgt_3_84;
		WeightsStore3[85] <= Wgt_3_85;
		WeightsStore3[86] <= Wgt_3_86;
		WeightsStore3[87] <= Wgt_3_87;
		WeightsStore3[88] <= Wgt_3_88;
		WeightsStore3[89] <= Wgt_3_89;
		WeightsStore3[90] <= Wgt_3_90;
		WeightsStore3[91] <= Wgt_3_91;
		WeightsStore3[92] <= Wgt_3_92;
		WeightsStore3[93] <= Wgt_3_93;
		WeightsStore3[94] <= Wgt_3_94;
		WeightsStore3[95] <= Wgt_3_95;
		WeightsStore3[96] <= Wgt_3_96;
		WeightsStore3[97] <= Wgt_3_97;
		WeightsStore3[98] <= Wgt_3_98;
		WeightsStore3[99] <= Wgt_3_99;
		WeightsStore3[100] <= Wgt_3_100;
		WeightsStore3[101] <= Wgt_3_101;
		WeightsStore3[102] <= Wgt_3_102;
		WeightsStore3[103] <= Wgt_3_103;
		WeightsStore3[104] <= Wgt_3_104;
		WeightsStore3[105] <= Wgt_3_105;
		WeightsStore3[106] <= Wgt_3_106;
		WeightsStore3[107] <= Wgt_3_107;
		WeightsStore3[108] <= Wgt_3_108;
		WeightsStore3[109] <= Wgt_3_109;
		WeightsStore3[110] <= Wgt_3_110;
		WeightsStore3[111] <= Wgt_3_111;
		WeightsStore3[112] <= Wgt_3_112;
		WeightsStore3[113] <= Wgt_3_113;
		WeightsStore3[114] <= Wgt_3_114;
		WeightsStore3[115] <= Wgt_3_115;
		WeightsStore3[116] <= Wgt_3_116;
		WeightsStore3[117] <= Wgt_3_117;
		WeightsStore3[118] <= Wgt_3_118;
		WeightsStore3[119] <= Wgt_3_119;
		WeightsStore3[120] <= Wgt_3_120;
		WeightsStore3[121] <= Wgt_3_121;
		WeightsStore3[122] <= Wgt_3_122;
		WeightsStore3[123] <= Wgt_3_123;
		WeightsStore3[124] <= Wgt_3_124;
		WeightsStore3[125] <= Wgt_3_125;
		WeightsStore3[126] <= Wgt_3_126;
		WeightsStore3[127] <= Wgt_3_127;
		WeightsStore3[128] <= Wgt_3_128;
		WeightsStore3[129] <= Wgt_3_129;
		WeightsStore3[130] <= Wgt_3_130;
		WeightsStore3[131] <= Wgt_3_131;
		WeightsStore3[132] <= Wgt_3_132;
		WeightsStore3[133] <= Wgt_3_133;
		WeightsStore3[134] <= Wgt_3_134;
		WeightsStore3[135] <= Wgt_3_135;
		WeightsStore3[136] <= Wgt_3_136;
		WeightsStore3[137] <= Wgt_3_137;
		WeightsStore3[138] <= Wgt_3_138;
		WeightsStore3[139] <= Wgt_3_139;
		WeightsStore3[140] <= Wgt_3_140;
		WeightsStore3[141] <= Wgt_3_141;
		WeightsStore3[142] <= Wgt_3_142;
		WeightsStore3[143] <= Wgt_3_143;
		WeightsStore3[144] <= Wgt_3_144;
		WeightsStore3[145] <= Wgt_3_145;
		WeightsStore3[146] <= Wgt_3_146;
		WeightsStore3[147] <= Wgt_3_147;
		WeightsStore3[148] <= Wgt_3_148;
		WeightsStore3[149] <= Wgt_3_149;
		WeightsStore3[150] <= Wgt_3_150;
		WeightsStore3[151] <= Wgt_3_151;
		WeightsStore3[152] <= Wgt_3_152;
		WeightsStore3[153] <= Wgt_3_153;
		WeightsStore3[154] <= Wgt_3_154;
		WeightsStore3[155] <= Wgt_3_155;
		WeightsStore3[156] <= Wgt_3_156;
		WeightsStore3[157] <= Wgt_3_157;
		WeightsStore3[158] <= Wgt_3_158;
		WeightsStore3[159] <= Wgt_3_159;
		WeightsStore3[160] <= Wgt_3_160;
		WeightsStore3[161] <= Wgt_3_161;
		WeightsStore3[162] <= Wgt_3_162;
		WeightsStore3[163] <= Wgt_3_163;
		WeightsStore3[164] <= Wgt_3_164;
		WeightsStore3[165] <= Wgt_3_165;
		WeightsStore3[166] <= Wgt_3_166;
		WeightsStore3[167] <= Wgt_3_167;
		WeightsStore3[168] <= Wgt_3_168;
		WeightsStore3[169] <= Wgt_3_169;
		WeightsStore3[170] <= Wgt_3_170;
		WeightsStore3[171] <= Wgt_3_171;
		WeightsStore3[172] <= Wgt_3_172;
		WeightsStore3[173] <= Wgt_3_173;
		WeightsStore3[174] <= Wgt_3_174;
		WeightsStore3[175] <= Wgt_3_175;
		WeightsStore3[176] <= Wgt_3_176;
		WeightsStore3[177] <= Wgt_3_177;
		WeightsStore3[178] <= Wgt_3_178;
		WeightsStore3[179] <= Wgt_3_179;
		WeightsStore3[180] <= Wgt_3_180;
		WeightsStore3[181] <= Wgt_3_181;
		WeightsStore3[182] <= Wgt_3_182;
		WeightsStore3[183] <= Wgt_3_183;
		WeightsStore3[184] <= Wgt_3_184;
		WeightsStore3[185] <= Wgt_3_185;
		WeightsStore3[186] <= Wgt_3_186;
		WeightsStore3[187] <= Wgt_3_187;
		WeightsStore3[188] <= Wgt_3_188;
		WeightsStore3[189] <= Wgt_3_189;
		WeightsStore3[190] <= Wgt_3_190;
		WeightsStore3[191] <= Wgt_3_191;
		WeightsStore3[192] <= Wgt_3_192;
		WeightsStore3[193] <= Wgt_3_193;
		WeightsStore3[194] <= Wgt_3_194;
		WeightsStore3[195] <= Wgt_3_195;
		WeightsStore3[196] <= Wgt_3_196;
		WeightsStore3[197] <= Wgt_3_197;
		WeightsStore3[198] <= Wgt_3_198;
		WeightsStore3[199] <= Wgt_3_199;
		WeightsStore3[200] <= Wgt_3_200;
		WeightsStore3[201] <= Wgt_3_201;
		WeightsStore3[202] <= Wgt_3_202;
		WeightsStore3[203] <= Wgt_3_203;
		WeightsStore3[204] <= Wgt_3_204;
		WeightsStore3[205] <= Wgt_3_205;
		WeightsStore3[206] <= Wgt_3_206;
		WeightsStore3[207] <= Wgt_3_207;
		WeightsStore3[208] <= Wgt_3_208;
		WeightsStore3[209] <= Wgt_3_209;
		WeightsStore3[210] <= Wgt_3_210;
		WeightsStore3[211] <= Wgt_3_211;
		WeightsStore3[212] <= Wgt_3_212;
		WeightsStore3[213] <= Wgt_3_213;
		WeightsStore3[214] <= Wgt_3_214;
		WeightsStore3[215] <= Wgt_3_215;
		WeightsStore3[216] <= Wgt_3_216;
		WeightsStore3[217] <= Wgt_3_217;
		WeightsStore3[218] <= Wgt_3_218;
		WeightsStore3[219] <= Wgt_3_219;
		WeightsStore3[220] <= Wgt_3_220;
		WeightsStore3[221] <= Wgt_3_221;
		WeightsStore3[222] <= Wgt_3_222;
		WeightsStore3[223] <= Wgt_3_223;
		WeightsStore3[224] <= Wgt_3_224;
		WeightsStore3[225] <= Wgt_3_225;
		WeightsStore3[226] <= Wgt_3_226;
		WeightsStore3[227] <= Wgt_3_227;
		WeightsStore3[228] <= Wgt_3_228;
		WeightsStore3[229] <= Wgt_3_229;
		WeightsStore3[230] <= Wgt_3_230;
		WeightsStore3[231] <= Wgt_3_231;
		WeightsStore3[232] <= Wgt_3_232;
		WeightsStore3[233] <= Wgt_3_233;
		WeightsStore3[234] <= Wgt_3_234;
		WeightsStore3[235] <= Wgt_3_235;
		WeightsStore3[236] <= Wgt_3_236;
		WeightsStore3[237] <= Wgt_3_237;
		WeightsStore3[238] <= Wgt_3_238;
		WeightsStore3[239] <= Wgt_3_239;
		WeightsStore3[240] <= Wgt_3_240;
		WeightsStore3[241] <= Wgt_3_241;
		WeightsStore3[242] <= Wgt_3_242;
		WeightsStore3[243] <= Wgt_3_243;
		WeightsStore3[244] <= Wgt_3_244;
		WeightsStore3[245] <= Wgt_3_245;
		WeightsStore3[246] <= Wgt_3_246;
		WeightsStore3[247] <= Wgt_3_247;
		WeightsStore3[248] <= Wgt_3_248;
		WeightsStore3[249] <= Wgt_3_249;
		WeightsStore3[250] <= Wgt_3_250;
		WeightsStore3[251] <= Wgt_3_251;
		WeightsStore3[252] <= Wgt_3_252;
		WeightsStore3[253] <= Wgt_3_253;
		WeightsStore3[254] <= Wgt_3_254;
		WeightsStore3[255] <= Wgt_3_255;
		WeightsStore3[256] <= Wgt_3_256;
		WeightsStore3[257] <= Wgt_3_257;
		WeightsStore3[258] <= Wgt_3_258;
		WeightsStore3[259] <= Wgt_3_259;
		WeightsStore3[260] <= Wgt_3_260;
		WeightsStore3[261] <= Wgt_3_261;
		WeightsStore3[262] <= Wgt_3_262;
		WeightsStore3[263] <= Wgt_3_263;
		WeightsStore3[264] <= Wgt_3_264;
		WeightsStore3[265] <= Wgt_3_265;
		WeightsStore3[266] <= Wgt_3_266;
		WeightsStore3[267] <= Wgt_3_267;
		WeightsStore3[268] <= Wgt_3_268;
		WeightsStore3[269] <= Wgt_3_269;
		WeightsStore3[270] <= Wgt_3_270;
		WeightsStore3[271] <= Wgt_3_271;
		WeightsStore3[272] <= Wgt_3_272;
		WeightsStore3[273] <= Wgt_3_273;
		WeightsStore3[274] <= Wgt_3_274;
		WeightsStore3[275] <= Wgt_3_275;
		WeightsStore3[276] <= Wgt_3_276;
		WeightsStore3[277] <= Wgt_3_277;
		WeightsStore3[278] <= Wgt_3_278;
		WeightsStore3[279] <= Wgt_3_279;
		WeightsStore3[280] <= Wgt_3_280;
		WeightsStore3[281] <= Wgt_3_281;
		WeightsStore3[282] <= Wgt_3_282;
		WeightsStore3[283] <= Wgt_3_283;
		WeightsStore3[284] <= Wgt_3_284;
		WeightsStore3[285] <= Wgt_3_285;
		WeightsStore3[286] <= Wgt_3_286;
		WeightsStore3[287] <= Wgt_3_287;
		WeightsStore3[288] <= Wgt_3_288;
		WeightsStore3[289] <= Wgt_3_289;
		WeightsStore3[290] <= Wgt_3_290;
		WeightsStore3[291] <= Wgt_3_291;
		WeightsStore3[292] <= Wgt_3_292;
		WeightsStore3[293] <= Wgt_3_293;
		WeightsStore3[294] <= Wgt_3_294;
		WeightsStore3[295] <= Wgt_3_295;
		WeightsStore3[296] <= Wgt_3_296;
		WeightsStore3[297] <= Wgt_3_297;
		WeightsStore3[298] <= Wgt_3_298;
		WeightsStore3[299] <= Wgt_3_299;
		WeightsStore3[300] <= Wgt_3_300;
		WeightsStore3[301] <= Wgt_3_301;
		WeightsStore3[302] <= Wgt_3_302;
		WeightsStore3[303] <= Wgt_3_303;
		WeightsStore3[304] <= Wgt_3_304;
		WeightsStore3[305] <= Wgt_3_305;
		WeightsStore3[306] <= Wgt_3_306;
		WeightsStore3[307] <= Wgt_3_307;
		WeightsStore3[308] <= Wgt_3_308;
		WeightsStore3[309] <= Wgt_3_309;
		WeightsStore3[310] <= Wgt_3_310;
		WeightsStore3[311] <= Wgt_3_311;
		WeightsStore3[312] <= Wgt_3_312;
		WeightsStore3[313] <= Wgt_3_313;
		WeightsStore3[314] <= Wgt_3_314;
		WeightsStore3[315] <= Wgt_3_315;
		WeightsStore3[316] <= Wgt_3_316;
		WeightsStore3[317] <= Wgt_3_317;
		WeightsStore3[318] <= Wgt_3_318;
		WeightsStore3[319] <= Wgt_3_319;
		WeightsStore3[320] <= Wgt_3_320;
		WeightsStore3[321] <= Wgt_3_321;
		WeightsStore3[322] <= Wgt_3_322;
		WeightsStore3[323] <= Wgt_3_323;
		WeightsStore3[324] <= Wgt_3_324;
		WeightsStore3[325] <= Wgt_3_325;
		WeightsStore3[326] <= Wgt_3_326;
		WeightsStore3[327] <= Wgt_3_327;
		WeightsStore3[328] <= Wgt_3_328;
		WeightsStore3[329] <= Wgt_3_329;
		WeightsStore3[330] <= Wgt_3_330;
		WeightsStore3[331] <= Wgt_3_331;
		WeightsStore3[332] <= Wgt_3_332;
		WeightsStore3[333] <= Wgt_3_333;
		WeightsStore3[334] <= Wgt_3_334;
		WeightsStore3[335] <= Wgt_3_335;
		WeightsStore3[336] <= Wgt_3_336;
		WeightsStore3[337] <= Wgt_3_337;
		WeightsStore3[338] <= Wgt_3_338;
		WeightsStore3[339] <= Wgt_3_339;
		WeightsStore3[340] <= Wgt_3_340;
		WeightsStore3[341] <= Wgt_3_341;
		WeightsStore3[342] <= Wgt_3_342;
		WeightsStore3[343] <= Wgt_3_343;
		WeightsStore3[344] <= Wgt_3_344;
		WeightsStore3[345] <= Wgt_3_345;
		WeightsStore3[346] <= Wgt_3_346;
		WeightsStore3[347] <= Wgt_3_347;
		WeightsStore3[348] <= Wgt_3_348;
		WeightsStore3[349] <= Wgt_3_349;
		WeightsStore3[350] <= Wgt_3_350;
		WeightsStore3[351] <= Wgt_3_351;
		WeightsStore3[352] <= Wgt_3_352;
		WeightsStore3[353] <= Wgt_3_353;
		WeightsStore3[354] <= Wgt_3_354;
		WeightsStore3[355] <= Wgt_3_355;
		WeightsStore3[356] <= Wgt_3_356;
		WeightsStore3[357] <= Wgt_3_357;
		WeightsStore3[358] <= Wgt_3_358;
		WeightsStore3[359] <= Wgt_3_359;
		WeightsStore3[360] <= Wgt_3_360;
		WeightsStore3[361] <= Wgt_3_361;
		WeightsStore3[362] <= Wgt_3_362;
		WeightsStore3[363] <= Wgt_3_363;
		WeightsStore3[364] <= Wgt_3_364;
		WeightsStore3[365] <= Wgt_3_365;
		WeightsStore3[366] <= Wgt_3_366;
		WeightsStore3[367] <= Wgt_3_367;
		WeightsStore3[368] <= Wgt_3_368;
		WeightsStore3[369] <= Wgt_3_369;
		WeightsStore3[370] <= Wgt_3_370;
		WeightsStore3[371] <= Wgt_3_371;
		WeightsStore3[372] <= Wgt_3_372;
		WeightsStore3[373] <= Wgt_3_373;
		WeightsStore3[374] <= Wgt_3_374;
		WeightsStore3[375] <= Wgt_3_375;
		WeightsStore3[376] <= Wgt_3_376;
		WeightsStore3[377] <= Wgt_3_377;
		WeightsStore3[378] <= Wgt_3_378;
		WeightsStore3[379] <= Wgt_3_379;
		WeightsStore3[380] <= Wgt_3_380;
		WeightsStore3[381] <= Wgt_3_381;
		WeightsStore3[382] <= Wgt_3_382;
		WeightsStore3[383] <= Wgt_3_383;
		WeightsStore3[384] <= Wgt_3_384;
		WeightsStore3[385] <= Wgt_3_385;
		WeightsStore3[386] <= Wgt_3_386;
		WeightsStore3[387] <= Wgt_3_387;
		WeightsStore3[388] <= Wgt_3_388;
		WeightsStore3[389] <= Wgt_3_389;
		WeightsStore3[390] <= Wgt_3_390;
		WeightsStore3[391] <= Wgt_3_391;
		WeightsStore3[392] <= Wgt_3_392;
		WeightsStore3[393] <= Wgt_3_393;
		WeightsStore3[394] <= Wgt_3_394;
		WeightsStore3[395] <= Wgt_3_395;
		WeightsStore3[396] <= Wgt_3_396;
		WeightsStore3[397] <= Wgt_3_397;
		WeightsStore3[398] <= Wgt_3_398;
		WeightsStore3[399] <= Wgt_3_399;
		WeightsStore3[400] <= Wgt_3_400;
		WeightsStore3[401] <= Wgt_3_401;
		WeightsStore3[402] <= Wgt_3_402;
		WeightsStore3[403] <= Wgt_3_403;
		WeightsStore3[404] <= Wgt_3_404;
		WeightsStore3[405] <= Wgt_3_405;
		WeightsStore3[406] <= Wgt_3_406;
		WeightsStore3[407] <= Wgt_3_407;
		WeightsStore3[408] <= Wgt_3_408;
		WeightsStore3[409] <= Wgt_3_409;
		WeightsStore3[410] <= Wgt_3_410;
		WeightsStore3[411] <= Wgt_3_411;
		WeightsStore3[412] <= Wgt_3_412;
		WeightsStore3[413] <= Wgt_3_413;
		WeightsStore3[414] <= Wgt_3_414;
		WeightsStore3[415] <= Wgt_3_415;
		WeightsStore3[416] <= Wgt_3_416;
		WeightsStore3[417] <= Wgt_3_417;
		WeightsStore3[418] <= Wgt_3_418;
		WeightsStore3[419] <= Wgt_3_419;
		WeightsStore3[420] <= Wgt_3_420;
		WeightsStore3[421] <= Wgt_3_421;
		WeightsStore3[422] <= Wgt_3_422;
		WeightsStore3[423] <= Wgt_3_423;
		WeightsStore3[424] <= Wgt_3_424;
		WeightsStore3[425] <= Wgt_3_425;
		WeightsStore3[426] <= Wgt_3_426;
		WeightsStore3[427] <= Wgt_3_427;
		WeightsStore3[428] <= Wgt_3_428;
		WeightsStore3[429] <= Wgt_3_429;
		WeightsStore3[430] <= Wgt_3_430;
		WeightsStore3[431] <= Wgt_3_431;
		WeightsStore3[432] <= Wgt_3_432;
		WeightsStore3[433] <= Wgt_3_433;
		WeightsStore3[434] <= Wgt_3_434;
		WeightsStore3[435] <= Wgt_3_435;
		WeightsStore3[436] <= Wgt_3_436;
		WeightsStore3[437] <= Wgt_3_437;
		WeightsStore3[438] <= Wgt_3_438;
		WeightsStore3[439] <= Wgt_3_439;
		WeightsStore3[440] <= Wgt_3_440;
		WeightsStore3[441] <= Wgt_3_441;
		WeightsStore3[442] <= Wgt_3_442;
		WeightsStore3[443] <= Wgt_3_443;
		WeightsStore3[444] <= Wgt_3_444;
		WeightsStore3[445] <= Wgt_3_445;
		WeightsStore3[446] <= Wgt_3_446;
		WeightsStore3[447] <= Wgt_3_447;
		WeightsStore3[448] <= Wgt_3_448;
		WeightsStore3[449] <= Wgt_3_449;
		WeightsStore3[450] <= Wgt_3_450;
		WeightsStore3[451] <= Wgt_3_451;
		WeightsStore3[452] <= Wgt_3_452;
		WeightsStore3[453] <= Wgt_3_453;
		WeightsStore3[454] <= Wgt_3_454;
		WeightsStore3[455] <= Wgt_3_455;
		WeightsStore3[456] <= Wgt_3_456;
		WeightsStore3[457] <= Wgt_3_457;
		WeightsStore3[458] <= Wgt_3_458;
		WeightsStore3[459] <= Wgt_3_459;
		WeightsStore3[460] <= Wgt_3_460;
		WeightsStore3[461] <= Wgt_3_461;
		WeightsStore3[462] <= Wgt_3_462;
		WeightsStore3[463] <= Wgt_3_463;
		WeightsStore3[464] <= Wgt_3_464;
		WeightsStore3[465] <= Wgt_3_465;
		WeightsStore3[466] <= Wgt_3_466;
		WeightsStore3[467] <= Wgt_3_467;
		WeightsStore3[468] <= Wgt_3_468;
		WeightsStore3[469] <= Wgt_3_469;
		WeightsStore3[470] <= Wgt_3_470;
		WeightsStore3[471] <= Wgt_3_471;
		WeightsStore3[472] <= Wgt_3_472;
		WeightsStore3[473] <= Wgt_3_473;
		WeightsStore3[474] <= Wgt_3_474;
		WeightsStore3[475] <= Wgt_3_475;
		WeightsStore3[476] <= Wgt_3_476;
		WeightsStore3[477] <= Wgt_3_477;
		WeightsStore3[478] <= Wgt_3_478;
		WeightsStore3[479] <= Wgt_3_479;
		WeightsStore3[480] <= Wgt_3_480;
		WeightsStore3[481] <= Wgt_3_481;
		WeightsStore3[482] <= Wgt_3_482;
		WeightsStore3[483] <= Wgt_3_483;
		WeightsStore3[484] <= Wgt_3_484;
		WeightsStore3[485] <= Wgt_3_485;
		WeightsStore3[486] <= Wgt_3_486;
		WeightsStore3[487] <= Wgt_3_487;
		WeightsStore3[488] <= Wgt_3_488;
		WeightsStore3[489] <= Wgt_3_489;
		WeightsStore3[490] <= Wgt_3_490;
		WeightsStore3[491] <= Wgt_3_491;
		WeightsStore3[492] <= Wgt_3_492;
		WeightsStore3[493] <= Wgt_3_493;
		WeightsStore3[494] <= Wgt_3_494;
		WeightsStore3[495] <= Wgt_3_495;
		WeightsStore3[496] <= Wgt_3_496;
		WeightsStore3[497] <= Wgt_3_497;
		WeightsStore3[498] <= Wgt_3_498;
		WeightsStore3[499] <= Wgt_3_499;
		WeightsStore3[500] <= Wgt_3_500;
		WeightsStore3[501] <= Wgt_3_501;
		WeightsStore3[502] <= Wgt_3_502;
		WeightsStore3[503] <= Wgt_3_503;
		WeightsStore3[504] <= Wgt_3_504;
		WeightsStore3[505] <= Wgt_3_505;
		WeightsStore3[506] <= Wgt_3_506;
		WeightsStore3[507] <= Wgt_3_507;
		WeightsStore3[508] <= Wgt_3_508;
		WeightsStore3[509] <= Wgt_3_509;
		WeightsStore3[510] <= Wgt_3_510;
		WeightsStore3[511] <= Wgt_3_511;
		WeightsStore3[512] <= Wgt_3_512;
		WeightsStore3[513] <= Wgt_3_513;
		WeightsStore3[514] <= Wgt_3_514;
		WeightsStore3[515] <= Wgt_3_515;
		WeightsStore3[516] <= Wgt_3_516;
		WeightsStore3[517] <= Wgt_3_517;
		WeightsStore3[518] <= Wgt_3_518;
		WeightsStore3[519] <= Wgt_3_519;
		WeightsStore3[520] <= Wgt_3_520;
		WeightsStore3[521] <= Wgt_3_521;
		WeightsStore3[522] <= Wgt_3_522;
		WeightsStore3[523] <= Wgt_3_523;
		WeightsStore3[524] <= Wgt_3_524;
		WeightsStore3[525] <= Wgt_3_525;
		WeightsStore3[526] <= Wgt_3_526;
		WeightsStore3[527] <= Wgt_3_527;
		WeightsStore3[528] <= Wgt_3_528;
		WeightsStore3[529] <= Wgt_3_529;
		WeightsStore3[530] <= Wgt_3_530;
		WeightsStore3[531] <= Wgt_3_531;
		WeightsStore3[532] <= Wgt_3_532;
		WeightsStore3[533] <= Wgt_3_533;
		WeightsStore3[534] <= Wgt_3_534;
		WeightsStore3[535] <= Wgt_3_535;
		WeightsStore3[536] <= Wgt_3_536;
		WeightsStore3[537] <= Wgt_3_537;
		WeightsStore3[538] <= Wgt_3_538;
		WeightsStore3[539] <= Wgt_3_539;
		WeightsStore3[540] <= Wgt_3_540;
		WeightsStore3[541] <= Wgt_3_541;
		WeightsStore3[542] <= Wgt_3_542;
		WeightsStore3[543] <= Wgt_3_543;
		WeightsStore3[544] <= Wgt_3_544;
		WeightsStore3[545] <= Wgt_3_545;
		WeightsStore3[546] <= Wgt_3_546;
		WeightsStore3[547] <= Wgt_3_547;
		WeightsStore3[548] <= Wgt_3_548;
		WeightsStore3[549] <= Wgt_3_549;
		WeightsStore3[550] <= Wgt_3_550;
		WeightsStore3[551] <= Wgt_3_551;
		WeightsStore3[552] <= Wgt_3_552;
		WeightsStore3[553] <= Wgt_3_553;
		WeightsStore3[554] <= Wgt_3_554;
		WeightsStore3[555] <= Wgt_3_555;
		WeightsStore3[556] <= Wgt_3_556;
		WeightsStore3[557] <= Wgt_3_557;
		WeightsStore3[558] <= Wgt_3_558;
		WeightsStore3[559] <= Wgt_3_559;
		WeightsStore3[560] <= Wgt_3_560;
		WeightsStore3[561] <= Wgt_3_561;
		WeightsStore3[562] <= Wgt_3_562;
		WeightsStore3[563] <= Wgt_3_563;
		WeightsStore3[564] <= Wgt_3_564;
		WeightsStore3[565] <= Wgt_3_565;
		WeightsStore3[566] <= Wgt_3_566;
		WeightsStore3[567] <= Wgt_3_567;
		WeightsStore3[568] <= Wgt_3_568;
		WeightsStore3[569] <= Wgt_3_569;
		WeightsStore3[570] <= Wgt_3_570;
		WeightsStore3[571] <= Wgt_3_571;
		WeightsStore3[572] <= Wgt_3_572;
		WeightsStore3[573] <= Wgt_3_573;
		WeightsStore3[574] <= Wgt_3_574;
		WeightsStore3[575] <= Wgt_3_575;
		WeightsStore3[576] <= Wgt_3_576;
		WeightsStore3[577] <= Wgt_3_577;
		WeightsStore3[578] <= Wgt_3_578;
		WeightsStore3[579] <= Wgt_3_579;
		WeightsStore3[580] <= Wgt_3_580;
		WeightsStore3[581] <= Wgt_3_581;
		WeightsStore3[582] <= Wgt_3_582;
		WeightsStore3[583] <= Wgt_3_583;
		WeightsStore3[584] <= Wgt_3_584;
		WeightsStore3[585] <= Wgt_3_585;
		WeightsStore3[586] <= Wgt_3_586;
		WeightsStore3[587] <= Wgt_3_587;
		WeightsStore3[588] <= Wgt_3_588;
		WeightsStore3[589] <= Wgt_3_589;
		WeightsStore3[590] <= Wgt_3_590;
		WeightsStore3[591] <= Wgt_3_591;
		WeightsStore3[592] <= Wgt_3_592;
		WeightsStore3[593] <= Wgt_3_593;
		WeightsStore3[594] <= Wgt_3_594;
		WeightsStore3[595] <= Wgt_3_595;
		WeightsStore3[596] <= Wgt_3_596;
		WeightsStore3[597] <= Wgt_3_597;
		WeightsStore3[598] <= Wgt_3_598;
		WeightsStore3[599] <= Wgt_3_599;
		WeightsStore3[600] <= Wgt_3_600;
		WeightsStore3[601] <= Wgt_3_601;
		WeightsStore3[602] <= Wgt_3_602;
		WeightsStore3[603] <= Wgt_3_603;
		WeightsStore3[604] <= Wgt_3_604;
		WeightsStore3[605] <= Wgt_3_605;
		WeightsStore3[606] <= Wgt_3_606;
		WeightsStore3[607] <= Wgt_3_607;
		WeightsStore3[608] <= Wgt_3_608;
		WeightsStore3[609] <= Wgt_3_609;
		WeightsStore3[610] <= Wgt_3_610;
		WeightsStore3[611] <= Wgt_3_611;
		WeightsStore3[612] <= Wgt_3_612;
		WeightsStore3[613] <= Wgt_3_613;
		WeightsStore3[614] <= Wgt_3_614;
		WeightsStore3[615] <= Wgt_3_615;
		WeightsStore3[616] <= Wgt_3_616;
		WeightsStore3[617] <= Wgt_3_617;
		WeightsStore3[618] <= Wgt_3_618;
		WeightsStore3[619] <= Wgt_3_619;
		WeightsStore3[620] <= Wgt_3_620;
		WeightsStore3[621] <= Wgt_3_621;
		WeightsStore3[622] <= Wgt_3_622;
		WeightsStore3[623] <= Wgt_3_623;
		WeightsStore3[624] <= Wgt_3_624;
		WeightsStore3[625] <= Wgt_3_625;
		WeightsStore3[626] <= Wgt_3_626;
		WeightsStore3[627] <= Wgt_3_627;
		WeightsStore3[628] <= Wgt_3_628;
		WeightsStore3[629] <= Wgt_3_629;
		WeightsStore3[630] <= Wgt_3_630;
		WeightsStore3[631] <= Wgt_3_631;
		WeightsStore3[632] <= Wgt_3_632;
		WeightsStore3[633] <= Wgt_3_633;
		WeightsStore3[634] <= Wgt_3_634;
		WeightsStore3[635] <= Wgt_3_635;
		WeightsStore3[636] <= Wgt_3_636;
		WeightsStore3[637] <= Wgt_3_637;
		WeightsStore3[638] <= Wgt_3_638;
		WeightsStore3[639] <= Wgt_3_639;
		WeightsStore3[640] <= Wgt_3_640;
		WeightsStore3[641] <= Wgt_3_641;
		WeightsStore3[642] <= Wgt_3_642;
		WeightsStore3[643] <= Wgt_3_643;
		WeightsStore3[644] <= Wgt_3_644;
		WeightsStore3[645] <= Wgt_3_645;
		WeightsStore3[646] <= Wgt_3_646;
		WeightsStore3[647] <= Wgt_3_647;
		WeightsStore3[648] <= Wgt_3_648;
		WeightsStore3[649] <= Wgt_3_649;
		WeightsStore3[650] <= Wgt_3_650;
		WeightsStore3[651] <= Wgt_3_651;
		WeightsStore3[652] <= Wgt_3_652;
		WeightsStore3[653] <= Wgt_3_653;
		WeightsStore3[654] <= Wgt_3_654;
		WeightsStore3[655] <= Wgt_3_655;
		WeightsStore3[656] <= Wgt_3_656;
		WeightsStore3[657] <= Wgt_3_657;
		WeightsStore3[658] <= Wgt_3_658;
		WeightsStore3[659] <= Wgt_3_659;
		WeightsStore3[660] <= Wgt_3_660;
		WeightsStore3[661] <= Wgt_3_661;
		WeightsStore3[662] <= Wgt_3_662;
		WeightsStore3[663] <= Wgt_3_663;
		WeightsStore3[664] <= Wgt_3_664;
		WeightsStore3[665] <= Wgt_3_665;
		WeightsStore3[666] <= Wgt_3_666;
		WeightsStore3[667] <= Wgt_3_667;
		WeightsStore3[668] <= Wgt_3_668;
		WeightsStore3[669] <= Wgt_3_669;
		WeightsStore3[670] <= Wgt_3_670;
		WeightsStore3[671] <= Wgt_3_671;
		WeightsStore3[672] <= Wgt_3_672;
		WeightsStore3[673] <= Wgt_3_673;
		WeightsStore3[674] <= Wgt_3_674;
		WeightsStore3[675] <= Wgt_3_675;
		WeightsStore3[676] <= Wgt_3_676;
		WeightsStore3[677] <= Wgt_3_677;
		WeightsStore3[678] <= Wgt_3_678;
		WeightsStore3[679] <= Wgt_3_679;
		WeightsStore3[680] <= Wgt_3_680;
		WeightsStore3[681] <= Wgt_3_681;
		WeightsStore3[682] <= Wgt_3_682;
		WeightsStore3[683] <= Wgt_3_683;
		WeightsStore3[684] <= Wgt_3_684;
		WeightsStore3[685] <= Wgt_3_685;
		WeightsStore3[686] <= Wgt_3_686;
		WeightsStore3[687] <= Wgt_3_687;
		WeightsStore3[688] <= Wgt_3_688;
		WeightsStore3[689] <= Wgt_3_689;
		WeightsStore3[690] <= Wgt_3_690;
		WeightsStore3[691] <= Wgt_3_691;
		WeightsStore3[692] <= Wgt_3_692;
		WeightsStore3[693] <= Wgt_3_693;
		WeightsStore3[694] <= Wgt_3_694;
		WeightsStore3[695] <= Wgt_3_695;
		WeightsStore3[696] <= Wgt_3_696;
		WeightsStore3[697] <= Wgt_3_697;
		WeightsStore3[698] <= Wgt_3_698;
		WeightsStore3[699] <= Wgt_3_699;
		WeightsStore3[700] <= Wgt_3_700;
		WeightsStore3[701] <= Wgt_3_701;
		WeightsStore3[702] <= Wgt_3_702;
		WeightsStore3[703] <= Wgt_3_703;
		WeightsStore3[704] <= Wgt_3_704;
		WeightsStore3[705] <= Wgt_3_705;
		WeightsStore3[706] <= Wgt_3_706;
		WeightsStore3[707] <= Wgt_3_707;
		WeightsStore3[708] <= Wgt_3_708;
		WeightsStore3[709] <= Wgt_3_709;
		WeightsStore3[710] <= Wgt_3_710;
		WeightsStore3[711] <= Wgt_3_711;
		WeightsStore3[712] <= Wgt_3_712;
		WeightsStore3[713] <= Wgt_3_713;
		WeightsStore3[714] <= Wgt_3_714;
		WeightsStore3[715] <= Wgt_3_715;
		WeightsStore3[716] <= Wgt_3_716;
		WeightsStore3[717] <= Wgt_3_717;
		WeightsStore3[718] <= Wgt_3_718;
		WeightsStore3[719] <= Wgt_3_719;
		WeightsStore3[720] <= Wgt_3_720;
		WeightsStore3[721] <= Wgt_3_721;
		WeightsStore3[722] <= Wgt_3_722;
		WeightsStore3[723] <= Wgt_3_723;
		WeightsStore3[724] <= Wgt_3_724;
		WeightsStore3[725] <= Wgt_3_725;
		WeightsStore3[726] <= Wgt_3_726;
		WeightsStore3[727] <= Wgt_3_727;
		WeightsStore3[728] <= Wgt_3_728;
		WeightsStore3[729] <= Wgt_3_729;
		WeightsStore3[730] <= Wgt_3_730;
		WeightsStore3[731] <= Wgt_3_731;
		WeightsStore3[732] <= Wgt_3_732;
		WeightsStore3[733] <= Wgt_3_733;
		WeightsStore3[734] <= Wgt_3_734;
		WeightsStore3[735] <= Wgt_3_735;
		WeightsStore3[736] <= Wgt_3_736;
		WeightsStore3[737] <= Wgt_3_737;
		WeightsStore3[738] <= Wgt_3_738;
		WeightsStore3[739] <= Wgt_3_739;
		WeightsStore3[740] <= Wgt_3_740;
		WeightsStore3[741] <= Wgt_3_741;
		WeightsStore3[742] <= Wgt_3_742;
		WeightsStore3[743] <= Wgt_3_743;
		WeightsStore3[744] <= Wgt_3_744;
		WeightsStore3[745] <= Wgt_3_745;
		WeightsStore3[746] <= Wgt_3_746;
		WeightsStore3[747] <= Wgt_3_747;
		WeightsStore3[748] <= Wgt_3_748;
		WeightsStore3[749] <= Wgt_3_749;
		WeightsStore3[750] <= Wgt_3_750;
		WeightsStore3[751] <= Wgt_3_751;
		WeightsStore3[752] <= Wgt_3_752;
		WeightsStore3[753] <= Wgt_3_753;
		WeightsStore3[754] <= Wgt_3_754;
		WeightsStore3[755] <= Wgt_3_755;
		WeightsStore3[756] <= Wgt_3_756;
		WeightsStore3[757] <= Wgt_3_757;
		WeightsStore3[758] <= Wgt_3_758;
		WeightsStore3[759] <= Wgt_3_759;
		WeightsStore3[760] <= Wgt_3_760;
		WeightsStore3[761] <= Wgt_3_761;
		WeightsStore3[762] <= Wgt_3_762;
		WeightsStore3[763] <= Wgt_3_763;
		WeightsStore3[764] <= Wgt_3_764;
		WeightsStore3[765] <= Wgt_3_765;
		WeightsStore3[766] <= Wgt_3_766;
		WeightsStore3[767] <= Wgt_3_767;
		WeightsStore3[768] <= Wgt_3_768;
		WeightsStore3[769] <= Wgt_3_769;
		WeightsStore3[770] <= Wgt_3_770;
		WeightsStore3[771] <= Wgt_3_771;
		WeightsStore3[772] <= Wgt_3_772;
		WeightsStore3[773] <= Wgt_3_773;
		WeightsStore3[774] <= Wgt_3_774;
		WeightsStore3[775] <= Wgt_3_775;
		WeightsStore3[776] <= Wgt_3_776;
		WeightsStore3[777] <= Wgt_3_777;
		WeightsStore3[778] <= Wgt_3_778;
		WeightsStore3[779] <= Wgt_3_779;
		WeightsStore3[780] <= Wgt_3_780;
		WeightsStore3[781] <= Wgt_3_781;
		WeightsStore3[782] <= Wgt_3_782;
		WeightsStore3[783] <= Wgt_3_783;
		WeightsStore3[784] <= Wgt_3_784;
		WeightsStore4[0] <= Wgt_4_0;
		WeightsStore4[1] <= Wgt_4_1;
		WeightsStore4[2] <= Wgt_4_2;
		WeightsStore4[3] <= Wgt_4_3;
		WeightsStore4[4] <= Wgt_4_4;
		WeightsStore4[5] <= Wgt_4_5;
		WeightsStore4[6] <= Wgt_4_6;
		WeightsStore4[7] <= Wgt_4_7;
		WeightsStore4[8] <= Wgt_4_8;
		WeightsStore4[9] <= Wgt_4_9;
		WeightsStore4[10] <= Wgt_4_10;
		WeightsStore4[11] <= Wgt_4_11;
		WeightsStore4[12] <= Wgt_4_12;
		WeightsStore4[13] <= Wgt_4_13;
		WeightsStore4[14] <= Wgt_4_14;
		WeightsStore4[15] <= Wgt_4_15;
		WeightsStore4[16] <= Wgt_4_16;
		WeightsStore4[17] <= Wgt_4_17;
		WeightsStore4[18] <= Wgt_4_18;
		WeightsStore4[19] <= Wgt_4_19;
		WeightsStore4[20] <= Wgt_4_20;
		WeightsStore4[21] <= Wgt_4_21;
		WeightsStore4[22] <= Wgt_4_22;
		WeightsStore4[23] <= Wgt_4_23;
		WeightsStore4[24] <= Wgt_4_24;
		WeightsStore4[25] <= Wgt_4_25;
		WeightsStore4[26] <= Wgt_4_26;
		WeightsStore4[27] <= Wgt_4_27;
		WeightsStore4[28] <= Wgt_4_28;
		WeightsStore4[29] <= Wgt_4_29;
		WeightsStore4[30] <= Wgt_4_30;
		WeightsStore4[31] <= Wgt_4_31;
		WeightsStore4[32] <= Wgt_4_32;
		WeightsStore4[33] <= Wgt_4_33;
		WeightsStore4[34] <= Wgt_4_34;
		WeightsStore4[35] <= Wgt_4_35;
		WeightsStore4[36] <= Wgt_4_36;
		WeightsStore4[37] <= Wgt_4_37;
		WeightsStore4[38] <= Wgt_4_38;
		WeightsStore4[39] <= Wgt_4_39;
		WeightsStore4[40] <= Wgt_4_40;
		WeightsStore4[41] <= Wgt_4_41;
		WeightsStore4[42] <= Wgt_4_42;
		WeightsStore4[43] <= Wgt_4_43;
		WeightsStore4[44] <= Wgt_4_44;
		WeightsStore4[45] <= Wgt_4_45;
		WeightsStore4[46] <= Wgt_4_46;
		WeightsStore4[47] <= Wgt_4_47;
		WeightsStore4[48] <= Wgt_4_48;
		WeightsStore4[49] <= Wgt_4_49;
		WeightsStore4[50] <= Wgt_4_50;
		WeightsStore4[51] <= Wgt_4_51;
		WeightsStore4[52] <= Wgt_4_52;
		WeightsStore4[53] <= Wgt_4_53;
		WeightsStore4[54] <= Wgt_4_54;
		WeightsStore4[55] <= Wgt_4_55;
		WeightsStore4[56] <= Wgt_4_56;
		WeightsStore4[57] <= Wgt_4_57;
		WeightsStore4[58] <= Wgt_4_58;
		WeightsStore4[59] <= Wgt_4_59;
		WeightsStore4[60] <= Wgt_4_60;
		WeightsStore4[61] <= Wgt_4_61;
		WeightsStore4[62] <= Wgt_4_62;
		WeightsStore4[63] <= Wgt_4_63;
		WeightsStore4[64] <= Wgt_4_64;
		WeightsStore4[65] <= Wgt_4_65;
		WeightsStore4[66] <= Wgt_4_66;
		WeightsStore4[67] <= Wgt_4_67;
		WeightsStore4[68] <= Wgt_4_68;
		WeightsStore4[69] <= Wgt_4_69;
		WeightsStore4[70] <= Wgt_4_70;
		WeightsStore4[71] <= Wgt_4_71;
		WeightsStore4[72] <= Wgt_4_72;
		WeightsStore4[73] <= Wgt_4_73;
		WeightsStore4[74] <= Wgt_4_74;
		WeightsStore4[75] <= Wgt_4_75;
		WeightsStore4[76] <= Wgt_4_76;
		WeightsStore4[77] <= Wgt_4_77;
		WeightsStore4[78] <= Wgt_4_78;
		WeightsStore4[79] <= Wgt_4_79;
		WeightsStore4[80] <= Wgt_4_80;
		WeightsStore4[81] <= Wgt_4_81;
		WeightsStore4[82] <= Wgt_4_82;
		WeightsStore4[83] <= Wgt_4_83;
		WeightsStore4[84] <= Wgt_4_84;
		WeightsStore4[85] <= Wgt_4_85;
		WeightsStore4[86] <= Wgt_4_86;
		WeightsStore4[87] <= Wgt_4_87;
		WeightsStore4[88] <= Wgt_4_88;
		WeightsStore4[89] <= Wgt_4_89;
		WeightsStore4[90] <= Wgt_4_90;
		WeightsStore4[91] <= Wgt_4_91;
		WeightsStore4[92] <= Wgt_4_92;
		WeightsStore4[93] <= Wgt_4_93;
		WeightsStore4[94] <= Wgt_4_94;
		WeightsStore4[95] <= Wgt_4_95;
		WeightsStore4[96] <= Wgt_4_96;
		WeightsStore4[97] <= Wgt_4_97;
		WeightsStore4[98] <= Wgt_4_98;
		WeightsStore4[99] <= Wgt_4_99;
		WeightsStore4[100] <= Wgt_4_100;
		WeightsStore4[101] <= Wgt_4_101;
		WeightsStore4[102] <= Wgt_4_102;
		WeightsStore4[103] <= Wgt_4_103;
		WeightsStore4[104] <= Wgt_4_104;
		WeightsStore4[105] <= Wgt_4_105;
		WeightsStore4[106] <= Wgt_4_106;
		WeightsStore4[107] <= Wgt_4_107;
		WeightsStore4[108] <= Wgt_4_108;
		WeightsStore4[109] <= Wgt_4_109;
		WeightsStore4[110] <= Wgt_4_110;
		WeightsStore4[111] <= Wgt_4_111;
		WeightsStore4[112] <= Wgt_4_112;
		WeightsStore4[113] <= Wgt_4_113;
		WeightsStore4[114] <= Wgt_4_114;
		WeightsStore4[115] <= Wgt_4_115;
		WeightsStore4[116] <= Wgt_4_116;
		WeightsStore4[117] <= Wgt_4_117;
		WeightsStore4[118] <= Wgt_4_118;
		WeightsStore4[119] <= Wgt_4_119;
		WeightsStore4[120] <= Wgt_4_120;
		WeightsStore4[121] <= Wgt_4_121;
		WeightsStore4[122] <= Wgt_4_122;
		WeightsStore4[123] <= Wgt_4_123;
		WeightsStore4[124] <= Wgt_4_124;
		WeightsStore4[125] <= Wgt_4_125;
		WeightsStore4[126] <= Wgt_4_126;
		WeightsStore4[127] <= Wgt_4_127;
		WeightsStore4[128] <= Wgt_4_128;
		WeightsStore4[129] <= Wgt_4_129;
		WeightsStore4[130] <= Wgt_4_130;
		WeightsStore4[131] <= Wgt_4_131;
		WeightsStore4[132] <= Wgt_4_132;
		WeightsStore4[133] <= Wgt_4_133;
		WeightsStore4[134] <= Wgt_4_134;
		WeightsStore4[135] <= Wgt_4_135;
		WeightsStore4[136] <= Wgt_4_136;
		WeightsStore4[137] <= Wgt_4_137;
		WeightsStore4[138] <= Wgt_4_138;
		WeightsStore4[139] <= Wgt_4_139;
		WeightsStore4[140] <= Wgt_4_140;
		WeightsStore4[141] <= Wgt_4_141;
		WeightsStore4[142] <= Wgt_4_142;
		WeightsStore4[143] <= Wgt_4_143;
		WeightsStore4[144] <= Wgt_4_144;
		WeightsStore4[145] <= Wgt_4_145;
		WeightsStore4[146] <= Wgt_4_146;
		WeightsStore4[147] <= Wgt_4_147;
		WeightsStore4[148] <= Wgt_4_148;
		WeightsStore4[149] <= Wgt_4_149;
		WeightsStore4[150] <= Wgt_4_150;
		WeightsStore4[151] <= Wgt_4_151;
		WeightsStore4[152] <= Wgt_4_152;
		WeightsStore4[153] <= Wgt_4_153;
		WeightsStore4[154] <= Wgt_4_154;
		WeightsStore4[155] <= Wgt_4_155;
		WeightsStore4[156] <= Wgt_4_156;
		WeightsStore4[157] <= Wgt_4_157;
		WeightsStore4[158] <= Wgt_4_158;
		WeightsStore4[159] <= Wgt_4_159;
		WeightsStore4[160] <= Wgt_4_160;
		WeightsStore4[161] <= Wgt_4_161;
		WeightsStore4[162] <= Wgt_4_162;
		WeightsStore4[163] <= Wgt_4_163;
		WeightsStore4[164] <= Wgt_4_164;
		WeightsStore4[165] <= Wgt_4_165;
		WeightsStore4[166] <= Wgt_4_166;
		WeightsStore4[167] <= Wgt_4_167;
		WeightsStore4[168] <= Wgt_4_168;
		WeightsStore4[169] <= Wgt_4_169;
		WeightsStore4[170] <= Wgt_4_170;
		WeightsStore4[171] <= Wgt_4_171;
		WeightsStore4[172] <= Wgt_4_172;
		WeightsStore4[173] <= Wgt_4_173;
		WeightsStore4[174] <= Wgt_4_174;
		WeightsStore4[175] <= Wgt_4_175;
		WeightsStore4[176] <= Wgt_4_176;
		WeightsStore4[177] <= Wgt_4_177;
		WeightsStore4[178] <= Wgt_4_178;
		WeightsStore4[179] <= Wgt_4_179;
		WeightsStore4[180] <= Wgt_4_180;
		WeightsStore4[181] <= Wgt_4_181;
		WeightsStore4[182] <= Wgt_4_182;
		WeightsStore4[183] <= Wgt_4_183;
		WeightsStore4[184] <= Wgt_4_184;
		WeightsStore4[185] <= Wgt_4_185;
		WeightsStore4[186] <= Wgt_4_186;
		WeightsStore4[187] <= Wgt_4_187;
		WeightsStore4[188] <= Wgt_4_188;
		WeightsStore4[189] <= Wgt_4_189;
		WeightsStore4[190] <= Wgt_4_190;
		WeightsStore4[191] <= Wgt_4_191;
		WeightsStore4[192] <= Wgt_4_192;
		WeightsStore4[193] <= Wgt_4_193;
		WeightsStore4[194] <= Wgt_4_194;
		WeightsStore4[195] <= Wgt_4_195;
		WeightsStore4[196] <= Wgt_4_196;
		WeightsStore4[197] <= Wgt_4_197;
		WeightsStore4[198] <= Wgt_4_198;
		WeightsStore4[199] <= Wgt_4_199;
		WeightsStore4[200] <= Wgt_4_200;
		WeightsStore4[201] <= Wgt_4_201;
		WeightsStore4[202] <= Wgt_4_202;
		WeightsStore4[203] <= Wgt_4_203;
		WeightsStore4[204] <= Wgt_4_204;
		WeightsStore4[205] <= Wgt_4_205;
		WeightsStore4[206] <= Wgt_4_206;
		WeightsStore4[207] <= Wgt_4_207;
		WeightsStore4[208] <= Wgt_4_208;
		WeightsStore4[209] <= Wgt_4_209;
		WeightsStore4[210] <= Wgt_4_210;
		WeightsStore4[211] <= Wgt_4_211;
		WeightsStore4[212] <= Wgt_4_212;
		WeightsStore4[213] <= Wgt_4_213;
		WeightsStore4[214] <= Wgt_4_214;
		WeightsStore4[215] <= Wgt_4_215;
		WeightsStore4[216] <= Wgt_4_216;
		WeightsStore4[217] <= Wgt_4_217;
		WeightsStore4[218] <= Wgt_4_218;
		WeightsStore4[219] <= Wgt_4_219;
		WeightsStore4[220] <= Wgt_4_220;
		WeightsStore4[221] <= Wgt_4_221;
		WeightsStore4[222] <= Wgt_4_222;
		WeightsStore4[223] <= Wgt_4_223;
		WeightsStore4[224] <= Wgt_4_224;
		WeightsStore4[225] <= Wgt_4_225;
		WeightsStore4[226] <= Wgt_4_226;
		WeightsStore4[227] <= Wgt_4_227;
		WeightsStore4[228] <= Wgt_4_228;
		WeightsStore4[229] <= Wgt_4_229;
		WeightsStore4[230] <= Wgt_4_230;
		WeightsStore4[231] <= Wgt_4_231;
		WeightsStore4[232] <= Wgt_4_232;
		WeightsStore4[233] <= Wgt_4_233;
		WeightsStore4[234] <= Wgt_4_234;
		WeightsStore4[235] <= Wgt_4_235;
		WeightsStore4[236] <= Wgt_4_236;
		WeightsStore4[237] <= Wgt_4_237;
		WeightsStore4[238] <= Wgt_4_238;
		WeightsStore4[239] <= Wgt_4_239;
		WeightsStore4[240] <= Wgt_4_240;
		WeightsStore4[241] <= Wgt_4_241;
		WeightsStore4[242] <= Wgt_4_242;
		WeightsStore4[243] <= Wgt_4_243;
		WeightsStore4[244] <= Wgt_4_244;
		WeightsStore4[245] <= Wgt_4_245;
		WeightsStore4[246] <= Wgt_4_246;
		WeightsStore4[247] <= Wgt_4_247;
		WeightsStore4[248] <= Wgt_4_248;
		WeightsStore4[249] <= Wgt_4_249;
		WeightsStore4[250] <= Wgt_4_250;
		WeightsStore4[251] <= Wgt_4_251;
		WeightsStore4[252] <= Wgt_4_252;
		WeightsStore4[253] <= Wgt_4_253;
		WeightsStore4[254] <= Wgt_4_254;
		WeightsStore4[255] <= Wgt_4_255;
		WeightsStore4[256] <= Wgt_4_256;
		WeightsStore4[257] <= Wgt_4_257;
		WeightsStore4[258] <= Wgt_4_258;
		WeightsStore4[259] <= Wgt_4_259;
		WeightsStore4[260] <= Wgt_4_260;
		WeightsStore4[261] <= Wgt_4_261;
		WeightsStore4[262] <= Wgt_4_262;
		WeightsStore4[263] <= Wgt_4_263;
		WeightsStore4[264] <= Wgt_4_264;
		WeightsStore4[265] <= Wgt_4_265;
		WeightsStore4[266] <= Wgt_4_266;
		WeightsStore4[267] <= Wgt_4_267;
		WeightsStore4[268] <= Wgt_4_268;
		WeightsStore4[269] <= Wgt_4_269;
		WeightsStore4[270] <= Wgt_4_270;
		WeightsStore4[271] <= Wgt_4_271;
		WeightsStore4[272] <= Wgt_4_272;
		WeightsStore4[273] <= Wgt_4_273;
		WeightsStore4[274] <= Wgt_4_274;
		WeightsStore4[275] <= Wgt_4_275;
		WeightsStore4[276] <= Wgt_4_276;
		WeightsStore4[277] <= Wgt_4_277;
		WeightsStore4[278] <= Wgt_4_278;
		WeightsStore4[279] <= Wgt_4_279;
		WeightsStore4[280] <= Wgt_4_280;
		WeightsStore4[281] <= Wgt_4_281;
		WeightsStore4[282] <= Wgt_4_282;
		WeightsStore4[283] <= Wgt_4_283;
		WeightsStore4[284] <= Wgt_4_284;
		WeightsStore4[285] <= Wgt_4_285;
		WeightsStore4[286] <= Wgt_4_286;
		WeightsStore4[287] <= Wgt_4_287;
		WeightsStore4[288] <= Wgt_4_288;
		WeightsStore4[289] <= Wgt_4_289;
		WeightsStore4[290] <= Wgt_4_290;
		WeightsStore4[291] <= Wgt_4_291;
		WeightsStore4[292] <= Wgt_4_292;
		WeightsStore4[293] <= Wgt_4_293;
		WeightsStore4[294] <= Wgt_4_294;
		WeightsStore4[295] <= Wgt_4_295;
		WeightsStore4[296] <= Wgt_4_296;
		WeightsStore4[297] <= Wgt_4_297;
		WeightsStore4[298] <= Wgt_4_298;
		WeightsStore4[299] <= Wgt_4_299;
		WeightsStore4[300] <= Wgt_4_300;
		WeightsStore4[301] <= Wgt_4_301;
		WeightsStore4[302] <= Wgt_4_302;
		WeightsStore4[303] <= Wgt_4_303;
		WeightsStore4[304] <= Wgt_4_304;
		WeightsStore4[305] <= Wgt_4_305;
		WeightsStore4[306] <= Wgt_4_306;
		WeightsStore4[307] <= Wgt_4_307;
		WeightsStore4[308] <= Wgt_4_308;
		WeightsStore4[309] <= Wgt_4_309;
		WeightsStore4[310] <= Wgt_4_310;
		WeightsStore4[311] <= Wgt_4_311;
		WeightsStore4[312] <= Wgt_4_312;
		WeightsStore4[313] <= Wgt_4_313;
		WeightsStore4[314] <= Wgt_4_314;
		WeightsStore4[315] <= Wgt_4_315;
		WeightsStore4[316] <= Wgt_4_316;
		WeightsStore4[317] <= Wgt_4_317;
		WeightsStore4[318] <= Wgt_4_318;
		WeightsStore4[319] <= Wgt_4_319;
		WeightsStore4[320] <= Wgt_4_320;
		WeightsStore4[321] <= Wgt_4_321;
		WeightsStore4[322] <= Wgt_4_322;
		WeightsStore4[323] <= Wgt_4_323;
		WeightsStore4[324] <= Wgt_4_324;
		WeightsStore4[325] <= Wgt_4_325;
		WeightsStore4[326] <= Wgt_4_326;
		WeightsStore4[327] <= Wgt_4_327;
		WeightsStore4[328] <= Wgt_4_328;
		WeightsStore4[329] <= Wgt_4_329;
		WeightsStore4[330] <= Wgt_4_330;
		WeightsStore4[331] <= Wgt_4_331;
		WeightsStore4[332] <= Wgt_4_332;
		WeightsStore4[333] <= Wgt_4_333;
		WeightsStore4[334] <= Wgt_4_334;
		WeightsStore4[335] <= Wgt_4_335;
		WeightsStore4[336] <= Wgt_4_336;
		WeightsStore4[337] <= Wgt_4_337;
		WeightsStore4[338] <= Wgt_4_338;
		WeightsStore4[339] <= Wgt_4_339;
		WeightsStore4[340] <= Wgt_4_340;
		WeightsStore4[341] <= Wgt_4_341;
		WeightsStore4[342] <= Wgt_4_342;
		WeightsStore4[343] <= Wgt_4_343;
		WeightsStore4[344] <= Wgt_4_344;
		WeightsStore4[345] <= Wgt_4_345;
		WeightsStore4[346] <= Wgt_4_346;
		WeightsStore4[347] <= Wgt_4_347;
		WeightsStore4[348] <= Wgt_4_348;
		WeightsStore4[349] <= Wgt_4_349;
		WeightsStore4[350] <= Wgt_4_350;
		WeightsStore4[351] <= Wgt_4_351;
		WeightsStore4[352] <= Wgt_4_352;
		WeightsStore4[353] <= Wgt_4_353;
		WeightsStore4[354] <= Wgt_4_354;
		WeightsStore4[355] <= Wgt_4_355;
		WeightsStore4[356] <= Wgt_4_356;
		WeightsStore4[357] <= Wgt_4_357;
		WeightsStore4[358] <= Wgt_4_358;
		WeightsStore4[359] <= Wgt_4_359;
		WeightsStore4[360] <= Wgt_4_360;
		WeightsStore4[361] <= Wgt_4_361;
		WeightsStore4[362] <= Wgt_4_362;
		WeightsStore4[363] <= Wgt_4_363;
		WeightsStore4[364] <= Wgt_4_364;
		WeightsStore4[365] <= Wgt_4_365;
		WeightsStore4[366] <= Wgt_4_366;
		WeightsStore4[367] <= Wgt_4_367;
		WeightsStore4[368] <= Wgt_4_368;
		WeightsStore4[369] <= Wgt_4_369;
		WeightsStore4[370] <= Wgt_4_370;
		WeightsStore4[371] <= Wgt_4_371;
		WeightsStore4[372] <= Wgt_4_372;
		WeightsStore4[373] <= Wgt_4_373;
		WeightsStore4[374] <= Wgt_4_374;
		WeightsStore4[375] <= Wgt_4_375;
		WeightsStore4[376] <= Wgt_4_376;
		WeightsStore4[377] <= Wgt_4_377;
		WeightsStore4[378] <= Wgt_4_378;
		WeightsStore4[379] <= Wgt_4_379;
		WeightsStore4[380] <= Wgt_4_380;
		WeightsStore4[381] <= Wgt_4_381;
		WeightsStore4[382] <= Wgt_4_382;
		WeightsStore4[383] <= Wgt_4_383;
		WeightsStore4[384] <= Wgt_4_384;
		WeightsStore4[385] <= Wgt_4_385;
		WeightsStore4[386] <= Wgt_4_386;
		WeightsStore4[387] <= Wgt_4_387;
		WeightsStore4[388] <= Wgt_4_388;
		WeightsStore4[389] <= Wgt_4_389;
		WeightsStore4[390] <= Wgt_4_390;
		WeightsStore4[391] <= Wgt_4_391;
		WeightsStore4[392] <= Wgt_4_392;
		WeightsStore4[393] <= Wgt_4_393;
		WeightsStore4[394] <= Wgt_4_394;
		WeightsStore4[395] <= Wgt_4_395;
		WeightsStore4[396] <= Wgt_4_396;
		WeightsStore4[397] <= Wgt_4_397;
		WeightsStore4[398] <= Wgt_4_398;
		WeightsStore4[399] <= Wgt_4_399;
		WeightsStore4[400] <= Wgt_4_400;
		WeightsStore4[401] <= Wgt_4_401;
		WeightsStore4[402] <= Wgt_4_402;
		WeightsStore4[403] <= Wgt_4_403;
		WeightsStore4[404] <= Wgt_4_404;
		WeightsStore4[405] <= Wgt_4_405;
		WeightsStore4[406] <= Wgt_4_406;
		WeightsStore4[407] <= Wgt_4_407;
		WeightsStore4[408] <= Wgt_4_408;
		WeightsStore4[409] <= Wgt_4_409;
		WeightsStore4[410] <= Wgt_4_410;
		WeightsStore4[411] <= Wgt_4_411;
		WeightsStore4[412] <= Wgt_4_412;
		WeightsStore4[413] <= Wgt_4_413;
		WeightsStore4[414] <= Wgt_4_414;
		WeightsStore4[415] <= Wgt_4_415;
		WeightsStore4[416] <= Wgt_4_416;
		WeightsStore4[417] <= Wgt_4_417;
		WeightsStore4[418] <= Wgt_4_418;
		WeightsStore4[419] <= Wgt_4_419;
		WeightsStore4[420] <= Wgt_4_420;
		WeightsStore4[421] <= Wgt_4_421;
		WeightsStore4[422] <= Wgt_4_422;
		WeightsStore4[423] <= Wgt_4_423;
		WeightsStore4[424] <= Wgt_4_424;
		WeightsStore4[425] <= Wgt_4_425;
		WeightsStore4[426] <= Wgt_4_426;
		WeightsStore4[427] <= Wgt_4_427;
		WeightsStore4[428] <= Wgt_4_428;
		WeightsStore4[429] <= Wgt_4_429;
		WeightsStore4[430] <= Wgt_4_430;
		WeightsStore4[431] <= Wgt_4_431;
		WeightsStore4[432] <= Wgt_4_432;
		WeightsStore4[433] <= Wgt_4_433;
		WeightsStore4[434] <= Wgt_4_434;
		WeightsStore4[435] <= Wgt_4_435;
		WeightsStore4[436] <= Wgt_4_436;
		WeightsStore4[437] <= Wgt_4_437;
		WeightsStore4[438] <= Wgt_4_438;
		WeightsStore4[439] <= Wgt_4_439;
		WeightsStore4[440] <= Wgt_4_440;
		WeightsStore4[441] <= Wgt_4_441;
		WeightsStore4[442] <= Wgt_4_442;
		WeightsStore4[443] <= Wgt_4_443;
		WeightsStore4[444] <= Wgt_4_444;
		WeightsStore4[445] <= Wgt_4_445;
		WeightsStore4[446] <= Wgt_4_446;
		WeightsStore4[447] <= Wgt_4_447;
		WeightsStore4[448] <= Wgt_4_448;
		WeightsStore4[449] <= Wgt_4_449;
		WeightsStore4[450] <= Wgt_4_450;
		WeightsStore4[451] <= Wgt_4_451;
		WeightsStore4[452] <= Wgt_4_452;
		WeightsStore4[453] <= Wgt_4_453;
		WeightsStore4[454] <= Wgt_4_454;
		WeightsStore4[455] <= Wgt_4_455;
		WeightsStore4[456] <= Wgt_4_456;
		WeightsStore4[457] <= Wgt_4_457;
		WeightsStore4[458] <= Wgt_4_458;
		WeightsStore4[459] <= Wgt_4_459;
		WeightsStore4[460] <= Wgt_4_460;
		WeightsStore4[461] <= Wgt_4_461;
		WeightsStore4[462] <= Wgt_4_462;
		WeightsStore4[463] <= Wgt_4_463;
		WeightsStore4[464] <= Wgt_4_464;
		WeightsStore4[465] <= Wgt_4_465;
		WeightsStore4[466] <= Wgt_4_466;
		WeightsStore4[467] <= Wgt_4_467;
		WeightsStore4[468] <= Wgt_4_468;
		WeightsStore4[469] <= Wgt_4_469;
		WeightsStore4[470] <= Wgt_4_470;
		WeightsStore4[471] <= Wgt_4_471;
		WeightsStore4[472] <= Wgt_4_472;
		WeightsStore4[473] <= Wgt_4_473;
		WeightsStore4[474] <= Wgt_4_474;
		WeightsStore4[475] <= Wgt_4_475;
		WeightsStore4[476] <= Wgt_4_476;
		WeightsStore4[477] <= Wgt_4_477;
		WeightsStore4[478] <= Wgt_4_478;
		WeightsStore4[479] <= Wgt_4_479;
		WeightsStore4[480] <= Wgt_4_480;
		WeightsStore4[481] <= Wgt_4_481;
		WeightsStore4[482] <= Wgt_4_482;
		WeightsStore4[483] <= Wgt_4_483;
		WeightsStore4[484] <= Wgt_4_484;
		WeightsStore4[485] <= Wgt_4_485;
		WeightsStore4[486] <= Wgt_4_486;
		WeightsStore4[487] <= Wgt_4_487;
		WeightsStore4[488] <= Wgt_4_488;
		WeightsStore4[489] <= Wgt_4_489;
		WeightsStore4[490] <= Wgt_4_490;
		WeightsStore4[491] <= Wgt_4_491;
		WeightsStore4[492] <= Wgt_4_492;
		WeightsStore4[493] <= Wgt_4_493;
		WeightsStore4[494] <= Wgt_4_494;
		WeightsStore4[495] <= Wgt_4_495;
		WeightsStore4[496] <= Wgt_4_496;
		WeightsStore4[497] <= Wgt_4_497;
		WeightsStore4[498] <= Wgt_4_498;
		WeightsStore4[499] <= Wgt_4_499;
		WeightsStore4[500] <= Wgt_4_500;
		WeightsStore4[501] <= Wgt_4_501;
		WeightsStore4[502] <= Wgt_4_502;
		WeightsStore4[503] <= Wgt_4_503;
		WeightsStore4[504] <= Wgt_4_504;
		WeightsStore4[505] <= Wgt_4_505;
		WeightsStore4[506] <= Wgt_4_506;
		WeightsStore4[507] <= Wgt_4_507;
		WeightsStore4[508] <= Wgt_4_508;
		WeightsStore4[509] <= Wgt_4_509;
		WeightsStore4[510] <= Wgt_4_510;
		WeightsStore4[511] <= Wgt_4_511;
		WeightsStore4[512] <= Wgt_4_512;
		WeightsStore4[513] <= Wgt_4_513;
		WeightsStore4[514] <= Wgt_4_514;
		WeightsStore4[515] <= Wgt_4_515;
		WeightsStore4[516] <= Wgt_4_516;
		WeightsStore4[517] <= Wgt_4_517;
		WeightsStore4[518] <= Wgt_4_518;
		WeightsStore4[519] <= Wgt_4_519;
		WeightsStore4[520] <= Wgt_4_520;
		WeightsStore4[521] <= Wgt_4_521;
		WeightsStore4[522] <= Wgt_4_522;
		WeightsStore4[523] <= Wgt_4_523;
		WeightsStore4[524] <= Wgt_4_524;
		WeightsStore4[525] <= Wgt_4_525;
		WeightsStore4[526] <= Wgt_4_526;
		WeightsStore4[527] <= Wgt_4_527;
		WeightsStore4[528] <= Wgt_4_528;
		WeightsStore4[529] <= Wgt_4_529;
		WeightsStore4[530] <= Wgt_4_530;
		WeightsStore4[531] <= Wgt_4_531;
		WeightsStore4[532] <= Wgt_4_532;
		WeightsStore4[533] <= Wgt_4_533;
		WeightsStore4[534] <= Wgt_4_534;
		WeightsStore4[535] <= Wgt_4_535;
		WeightsStore4[536] <= Wgt_4_536;
		WeightsStore4[537] <= Wgt_4_537;
		WeightsStore4[538] <= Wgt_4_538;
		WeightsStore4[539] <= Wgt_4_539;
		WeightsStore4[540] <= Wgt_4_540;
		WeightsStore4[541] <= Wgt_4_541;
		WeightsStore4[542] <= Wgt_4_542;
		WeightsStore4[543] <= Wgt_4_543;
		WeightsStore4[544] <= Wgt_4_544;
		WeightsStore4[545] <= Wgt_4_545;
		WeightsStore4[546] <= Wgt_4_546;
		WeightsStore4[547] <= Wgt_4_547;
		WeightsStore4[548] <= Wgt_4_548;
		WeightsStore4[549] <= Wgt_4_549;
		WeightsStore4[550] <= Wgt_4_550;
		WeightsStore4[551] <= Wgt_4_551;
		WeightsStore4[552] <= Wgt_4_552;
		WeightsStore4[553] <= Wgt_4_553;
		WeightsStore4[554] <= Wgt_4_554;
		WeightsStore4[555] <= Wgt_4_555;
		WeightsStore4[556] <= Wgt_4_556;
		WeightsStore4[557] <= Wgt_4_557;
		WeightsStore4[558] <= Wgt_4_558;
		WeightsStore4[559] <= Wgt_4_559;
		WeightsStore4[560] <= Wgt_4_560;
		WeightsStore4[561] <= Wgt_4_561;
		WeightsStore4[562] <= Wgt_4_562;
		WeightsStore4[563] <= Wgt_4_563;
		WeightsStore4[564] <= Wgt_4_564;
		WeightsStore4[565] <= Wgt_4_565;
		WeightsStore4[566] <= Wgt_4_566;
		WeightsStore4[567] <= Wgt_4_567;
		WeightsStore4[568] <= Wgt_4_568;
		WeightsStore4[569] <= Wgt_4_569;
		WeightsStore4[570] <= Wgt_4_570;
		WeightsStore4[571] <= Wgt_4_571;
		WeightsStore4[572] <= Wgt_4_572;
		WeightsStore4[573] <= Wgt_4_573;
		WeightsStore4[574] <= Wgt_4_574;
		WeightsStore4[575] <= Wgt_4_575;
		WeightsStore4[576] <= Wgt_4_576;
		WeightsStore4[577] <= Wgt_4_577;
		WeightsStore4[578] <= Wgt_4_578;
		WeightsStore4[579] <= Wgt_4_579;
		WeightsStore4[580] <= Wgt_4_580;
		WeightsStore4[581] <= Wgt_4_581;
		WeightsStore4[582] <= Wgt_4_582;
		WeightsStore4[583] <= Wgt_4_583;
		WeightsStore4[584] <= Wgt_4_584;
		WeightsStore4[585] <= Wgt_4_585;
		WeightsStore4[586] <= Wgt_4_586;
		WeightsStore4[587] <= Wgt_4_587;
		WeightsStore4[588] <= Wgt_4_588;
		WeightsStore4[589] <= Wgt_4_589;
		WeightsStore4[590] <= Wgt_4_590;
		WeightsStore4[591] <= Wgt_4_591;
		WeightsStore4[592] <= Wgt_4_592;
		WeightsStore4[593] <= Wgt_4_593;
		WeightsStore4[594] <= Wgt_4_594;
		WeightsStore4[595] <= Wgt_4_595;
		WeightsStore4[596] <= Wgt_4_596;
		WeightsStore4[597] <= Wgt_4_597;
		WeightsStore4[598] <= Wgt_4_598;
		WeightsStore4[599] <= Wgt_4_599;
		WeightsStore4[600] <= Wgt_4_600;
		WeightsStore4[601] <= Wgt_4_601;
		WeightsStore4[602] <= Wgt_4_602;
		WeightsStore4[603] <= Wgt_4_603;
		WeightsStore4[604] <= Wgt_4_604;
		WeightsStore4[605] <= Wgt_4_605;
		WeightsStore4[606] <= Wgt_4_606;
		WeightsStore4[607] <= Wgt_4_607;
		WeightsStore4[608] <= Wgt_4_608;
		WeightsStore4[609] <= Wgt_4_609;
		WeightsStore4[610] <= Wgt_4_610;
		WeightsStore4[611] <= Wgt_4_611;
		WeightsStore4[612] <= Wgt_4_612;
		WeightsStore4[613] <= Wgt_4_613;
		WeightsStore4[614] <= Wgt_4_614;
		WeightsStore4[615] <= Wgt_4_615;
		WeightsStore4[616] <= Wgt_4_616;
		WeightsStore4[617] <= Wgt_4_617;
		WeightsStore4[618] <= Wgt_4_618;
		WeightsStore4[619] <= Wgt_4_619;
		WeightsStore4[620] <= Wgt_4_620;
		WeightsStore4[621] <= Wgt_4_621;
		WeightsStore4[622] <= Wgt_4_622;
		WeightsStore4[623] <= Wgt_4_623;
		WeightsStore4[624] <= Wgt_4_624;
		WeightsStore4[625] <= Wgt_4_625;
		WeightsStore4[626] <= Wgt_4_626;
		WeightsStore4[627] <= Wgt_4_627;
		WeightsStore4[628] <= Wgt_4_628;
		WeightsStore4[629] <= Wgt_4_629;
		WeightsStore4[630] <= Wgt_4_630;
		WeightsStore4[631] <= Wgt_4_631;
		WeightsStore4[632] <= Wgt_4_632;
		WeightsStore4[633] <= Wgt_4_633;
		WeightsStore4[634] <= Wgt_4_634;
		WeightsStore4[635] <= Wgt_4_635;
		WeightsStore4[636] <= Wgt_4_636;
		WeightsStore4[637] <= Wgt_4_637;
		WeightsStore4[638] <= Wgt_4_638;
		WeightsStore4[639] <= Wgt_4_639;
		WeightsStore4[640] <= Wgt_4_640;
		WeightsStore4[641] <= Wgt_4_641;
		WeightsStore4[642] <= Wgt_4_642;
		WeightsStore4[643] <= Wgt_4_643;
		WeightsStore4[644] <= Wgt_4_644;
		WeightsStore4[645] <= Wgt_4_645;
		WeightsStore4[646] <= Wgt_4_646;
		WeightsStore4[647] <= Wgt_4_647;
		WeightsStore4[648] <= Wgt_4_648;
		WeightsStore4[649] <= Wgt_4_649;
		WeightsStore4[650] <= Wgt_4_650;
		WeightsStore4[651] <= Wgt_4_651;
		WeightsStore4[652] <= Wgt_4_652;
		WeightsStore4[653] <= Wgt_4_653;
		WeightsStore4[654] <= Wgt_4_654;
		WeightsStore4[655] <= Wgt_4_655;
		WeightsStore4[656] <= Wgt_4_656;
		WeightsStore4[657] <= Wgt_4_657;
		WeightsStore4[658] <= Wgt_4_658;
		WeightsStore4[659] <= Wgt_4_659;
		WeightsStore4[660] <= Wgt_4_660;
		WeightsStore4[661] <= Wgt_4_661;
		WeightsStore4[662] <= Wgt_4_662;
		WeightsStore4[663] <= Wgt_4_663;
		WeightsStore4[664] <= Wgt_4_664;
		WeightsStore4[665] <= Wgt_4_665;
		WeightsStore4[666] <= Wgt_4_666;
		WeightsStore4[667] <= Wgt_4_667;
		WeightsStore4[668] <= Wgt_4_668;
		WeightsStore4[669] <= Wgt_4_669;
		WeightsStore4[670] <= Wgt_4_670;
		WeightsStore4[671] <= Wgt_4_671;
		WeightsStore4[672] <= Wgt_4_672;
		WeightsStore4[673] <= Wgt_4_673;
		WeightsStore4[674] <= Wgt_4_674;
		WeightsStore4[675] <= Wgt_4_675;
		WeightsStore4[676] <= Wgt_4_676;
		WeightsStore4[677] <= Wgt_4_677;
		WeightsStore4[678] <= Wgt_4_678;
		WeightsStore4[679] <= Wgt_4_679;
		WeightsStore4[680] <= Wgt_4_680;
		WeightsStore4[681] <= Wgt_4_681;
		WeightsStore4[682] <= Wgt_4_682;
		WeightsStore4[683] <= Wgt_4_683;
		WeightsStore4[684] <= Wgt_4_684;
		WeightsStore4[685] <= Wgt_4_685;
		WeightsStore4[686] <= Wgt_4_686;
		WeightsStore4[687] <= Wgt_4_687;
		WeightsStore4[688] <= Wgt_4_688;
		WeightsStore4[689] <= Wgt_4_689;
		WeightsStore4[690] <= Wgt_4_690;
		WeightsStore4[691] <= Wgt_4_691;
		WeightsStore4[692] <= Wgt_4_692;
		WeightsStore4[693] <= Wgt_4_693;
		WeightsStore4[694] <= Wgt_4_694;
		WeightsStore4[695] <= Wgt_4_695;
		WeightsStore4[696] <= Wgt_4_696;
		WeightsStore4[697] <= Wgt_4_697;
		WeightsStore4[698] <= Wgt_4_698;
		WeightsStore4[699] <= Wgt_4_699;
		WeightsStore4[700] <= Wgt_4_700;
		WeightsStore4[701] <= Wgt_4_701;
		WeightsStore4[702] <= Wgt_4_702;
		WeightsStore4[703] <= Wgt_4_703;
		WeightsStore4[704] <= Wgt_4_704;
		WeightsStore4[705] <= Wgt_4_705;
		WeightsStore4[706] <= Wgt_4_706;
		WeightsStore4[707] <= Wgt_4_707;
		WeightsStore4[708] <= Wgt_4_708;
		WeightsStore4[709] <= Wgt_4_709;
		WeightsStore4[710] <= Wgt_4_710;
		WeightsStore4[711] <= Wgt_4_711;
		WeightsStore4[712] <= Wgt_4_712;
		WeightsStore4[713] <= Wgt_4_713;
		WeightsStore4[714] <= Wgt_4_714;
		WeightsStore4[715] <= Wgt_4_715;
		WeightsStore4[716] <= Wgt_4_716;
		WeightsStore4[717] <= Wgt_4_717;
		WeightsStore4[718] <= Wgt_4_718;
		WeightsStore4[719] <= Wgt_4_719;
		WeightsStore4[720] <= Wgt_4_720;
		WeightsStore4[721] <= Wgt_4_721;
		WeightsStore4[722] <= Wgt_4_722;
		WeightsStore4[723] <= Wgt_4_723;
		WeightsStore4[724] <= Wgt_4_724;
		WeightsStore4[725] <= Wgt_4_725;
		WeightsStore4[726] <= Wgt_4_726;
		WeightsStore4[727] <= Wgt_4_727;
		WeightsStore4[728] <= Wgt_4_728;
		WeightsStore4[729] <= Wgt_4_729;
		WeightsStore4[730] <= Wgt_4_730;
		WeightsStore4[731] <= Wgt_4_731;
		WeightsStore4[732] <= Wgt_4_732;
		WeightsStore4[733] <= Wgt_4_733;
		WeightsStore4[734] <= Wgt_4_734;
		WeightsStore4[735] <= Wgt_4_735;
		WeightsStore4[736] <= Wgt_4_736;
		WeightsStore4[737] <= Wgt_4_737;
		WeightsStore4[738] <= Wgt_4_738;
		WeightsStore4[739] <= Wgt_4_739;
		WeightsStore4[740] <= Wgt_4_740;
		WeightsStore4[741] <= Wgt_4_741;
		WeightsStore4[742] <= Wgt_4_742;
		WeightsStore4[743] <= Wgt_4_743;
		WeightsStore4[744] <= Wgt_4_744;
		WeightsStore4[745] <= Wgt_4_745;
		WeightsStore4[746] <= Wgt_4_746;
		WeightsStore4[747] <= Wgt_4_747;
		WeightsStore4[748] <= Wgt_4_748;
		WeightsStore4[749] <= Wgt_4_749;
		WeightsStore4[750] <= Wgt_4_750;
		WeightsStore4[751] <= Wgt_4_751;
		WeightsStore4[752] <= Wgt_4_752;
		WeightsStore4[753] <= Wgt_4_753;
		WeightsStore4[754] <= Wgt_4_754;
		WeightsStore4[755] <= Wgt_4_755;
		WeightsStore4[756] <= Wgt_4_756;
		WeightsStore4[757] <= Wgt_4_757;
		WeightsStore4[758] <= Wgt_4_758;
		WeightsStore4[759] <= Wgt_4_759;
		WeightsStore4[760] <= Wgt_4_760;
		WeightsStore4[761] <= Wgt_4_761;
		WeightsStore4[762] <= Wgt_4_762;
		WeightsStore4[763] <= Wgt_4_763;
		WeightsStore4[764] <= Wgt_4_764;
		WeightsStore4[765] <= Wgt_4_765;
		WeightsStore4[766] <= Wgt_4_766;
		WeightsStore4[767] <= Wgt_4_767;
		WeightsStore4[768] <= Wgt_4_768;
		WeightsStore4[769] <= Wgt_4_769;
		WeightsStore4[770] <= Wgt_4_770;
		WeightsStore4[771] <= Wgt_4_771;
		WeightsStore4[772] <= Wgt_4_772;
		WeightsStore4[773] <= Wgt_4_773;
		WeightsStore4[774] <= Wgt_4_774;
		WeightsStore4[775] <= Wgt_4_775;
		WeightsStore4[776] <= Wgt_4_776;
		WeightsStore4[777] <= Wgt_4_777;
		WeightsStore4[778] <= Wgt_4_778;
		WeightsStore4[779] <= Wgt_4_779;
		WeightsStore4[780] <= Wgt_4_780;
		WeightsStore4[781] <= Wgt_4_781;
		WeightsStore4[782] <= Wgt_4_782;
		WeightsStore4[783] <= Wgt_4_783;
		WeightsStore4[784] <= Wgt_4_784;
		WeightsStore5[0] <= Wgt_5_0;
		WeightsStore5[1] <= Wgt_5_1;
		WeightsStore5[2] <= Wgt_5_2;
		WeightsStore5[3] <= Wgt_5_3;
		WeightsStore5[4] <= Wgt_5_4;
		WeightsStore5[5] <= Wgt_5_5;
		WeightsStore5[6] <= Wgt_5_6;
		WeightsStore5[7] <= Wgt_5_7;
		WeightsStore5[8] <= Wgt_5_8;
		WeightsStore5[9] <= Wgt_5_9;
		WeightsStore5[10] <= Wgt_5_10;
		WeightsStore5[11] <= Wgt_5_11;
		WeightsStore5[12] <= Wgt_5_12;
		WeightsStore5[13] <= Wgt_5_13;
		WeightsStore5[14] <= Wgt_5_14;
		WeightsStore5[15] <= Wgt_5_15;
		WeightsStore5[16] <= Wgt_5_16;
		WeightsStore5[17] <= Wgt_5_17;
		WeightsStore5[18] <= Wgt_5_18;
		WeightsStore5[19] <= Wgt_5_19;
		WeightsStore5[20] <= Wgt_5_20;
		WeightsStore5[21] <= Wgt_5_21;
		WeightsStore5[22] <= Wgt_5_22;
		WeightsStore5[23] <= Wgt_5_23;
		WeightsStore5[24] <= Wgt_5_24;
		WeightsStore5[25] <= Wgt_5_25;
		WeightsStore5[26] <= Wgt_5_26;
		WeightsStore5[27] <= Wgt_5_27;
		WeightsStore5[28] <= Wgt_5_28;
		WeightsStore5[29] <= Wgt_5_29;
		WeightsStore5[30] <= Wgt_5_30;
		WeightsStore5[31] <= Wgt_5_31;
		WeightsStore5[32] <= Wgt_5_32;
		WeightsStore5[33] <= Wgt_5_33;
		WeightsStore5[34] <= Wgt_5_34;
		WeightsStore5[35] <= Wgt_5_35;
		WeightsStore5[36] <= Wgt_5_36;
		WeightsStore5[37] <= Wgt_5_37;
		WeightsStore5[38] <= Wgt_5_38;
		WeightsStore5[39] <= Wgt_5_39;
		WeightsStore5[40] <= Wgt_5_40;
		WeightsStore5[41] <= Wgt_5_41;
		WeightsStore5[42] <= Wgt_5_42;
		WeightsStore5[43] <= Wgt_5_43;
		WeightsStore5[44] <= Wgt_5_44;
		WeightsStore5[45] <= Wgt_5_45;
		WeightsStore5[46] <= Wgt_5_46;
		WeightsStore5[47] <= Wgt_5_47;
		WeightsStore5[48] <= Wgt_5_48;
		WeightsStore5[49] <= Wgt_5_49;
		WeightsStore5[50] <= Wgt_5_50;
		WeightsStore5[51] <= Wgt_5_51;
		WeightsStore5[52] <= Wgt_5_52;
		WeightsStore5[53] <= Wgt_5_53;
		WeightsStore5[54] <= Wgt_5_54;
		WeightsStore5[55] <= Wgt_5_55;
		WeightsStore5[56] <= Wgt_5_56;
		WeightsStore5[57] <= Wgt_5_57;
		WeightsStore5[58] <= Wgt_5_58;
		WeightsStore5[59] <= Wgt_5_59;
		WeightsStore5[60] <= Wgt_5_60;
		WeightsStore5[61] <= Wgt_5_61;
		WeightsStore5[62] <= Wgt_5_62;
		WeightsStore5[63] <= Wgt_5_63;
		WeightsStore5[64] <= Wgt_5_64;
		WeightsStore5[65] <= Wgt_5_65;
		WeightsStore5[66] <= Wgt_5_66;
		WeightsStore5[67] <= Wgt_5_67;
		WeightsStore5[68] <= Wgt_5_68;
		WeightsStore5[69] <= Wgt_5_69;
		WeightsStore5[70] <= Wgt_5_70;
		WeightsStore5[71] <= Wgt_5_71;
		WeightsStore5[72] <= Wgt_5_72;
		WeightsStore5[73] <= Wgt_5_73;
		WeightsStore5[74] <= Wgt_5_74;
		WeightsStore5[75] <= Wgt_5_75;
		WeightsStore5[76] <= Wgt_5_76;
		WeightsStore5[77] <= Wgt_5_77;
		WeightsStore5[78] <= Wgt_5_78;
		WeightsStore5[79] <= Wgt_5_79;
		WeightsStore5[80] <= Wgt_5_80;
		WeightsStore5[81] <= Wgt_5_81;
		WeightsStore5[82] <= Wgt_5_82;
		WeightsStore5[83] <= Wgt_5_83;
		WeightsStore5[84] <= Wgt_5_84;
		WeightsStore5[85] <= Wgt_5_85;
		WeightsStore5[86] <= Wgt_5_86;
		WeightsStore5[87] <= Wgt_5_87;
		WeightsStore5[88] <= Wgt_5_88;
		WeightsStore5[89] <= Wgt_5_89;
		WeightsStore5[90] <= Wgt_5_90;
		WeightsStore5[91] <= Wgt_5_91;
		WeightsStore5[92] <= Wgt_5_92;
		WeightsStore5[93] <= Wgt_5_93;
		WeightsStore5[94] <= Wgt_5_94;
		WeightsStore5[95] <= Wgt_5_95;
		WeightsStore5[96] <= Wgt_5_96;
		WeightsStore5[97] <= Wgt_5_97;
		WeightsStore5[98] <= Wgt_5_98;
		WeightsStore5[99] <= Wgt_5_99;
		WeightsStore5[100] <= Wgt_5_100;
		WeightsStore5[101] <= Wgt_5_101;
		WeightsStore5[102] <= Wgt_5_102;
		WeightsStore5[103] <= Wgt_5_103;
		WeightsStore5[104] <= Wgt_5_104;
		WeightsStore5[105] <= Wgt_5_105;
		WeightsStore5[106] <= Wgt_5_106;
		WeightsStore5[107] <= Wgt_5_107;
		WeightsStore5[108] <= Wgt_5_108;
		WeightsStore5[109] <= Wgt_5_109;
		WeightsStore5[110] <= Wgt_5_110;
		WeightsStore5[111] <= Wgt_5_111;
		WeightsStore5[112] <= Wgt_5_112;
		WeightsStore5[113] <= Wgt_5_113;
		WeightsStore5[114] <= Wgt_5_114;
		WeightsStore5[115] <= Wgt_5_115;
		WeightsStore5[116] <= Wgt_5_116;
		WeightsStore5[117] <= Wgt_5_117;
		WeightsStore5[118] <= Wgt_5_118;
		WeightsStore5[119] <= Wgt_5_119;
		WeightsStore5[120] <= Wgt_5_120;
		WeightsStore5[121] <= Wgt_5_121;
		WeightsStore5[122] <= Wgt_5_122;
		WeightsStore5[123] <= Wgt_5_123;
		WeightsStore5[124] <= Wgt_5_124;
		WeightsStore5[125] <= Wgt_5_125;
		WeightsStore5[126] <= Wgt_5_126;
		WeightsStore5[127] <= Wgt_5_127;
		WeightsStore5[128] <= Wgt_5_128;
		WeightsStore5[129] <= Wgt_5_129;
		WeightsStore5[130] <= Wgt_5_130;
		WeightsStore5[131] <= Wgt_5_131;
		WeightsStore5[132] <= Wgt_5_132;
		WeightsStore5[133] <= Wgt_5_133;
		WeightsStore5[134] <= Wgt_5_134;
		WeightsStore5[135] <= Wgt_5_135;
		WeightsStore5[136] <= Wgt_5_136;
		WeightsStore5[137] <= Wgt_5_137;
		WeightsStore5[138] <= Wgt_5_138;
		WeightsStore5[139] <= Wgt_5_139;
		WeightsStore5[140] <= Wgt_5_140;
		WeightsStore5[141] <= Wgt_5_141;
		WeightsStore5[142] <= Wgt_5_142;
		WeightsStore5[143] <= Wgt_5_143;
		WeightsStore5[144] <= Wgt_5_144;
		WeightsStore5[145] <= Wgt_5_145;
		WeightsStore5[146] <= Wgt_5_146;
		WeightsStore5[147] <= Wgt_5_147;
		WeightsStore5[148] <= Wgt_5_148;
		WeightsStore5[149] <= Wgt_5_149;
		WeightsStore5[150] <= Wgt_5_150;
		WeightsStore5[151] <= Wgt_5_151;
		WeightsStore5[152] <= Wgt_5_152;
		WeightsStore5[153] <= Wgt_5_153;
		WeightsStore5[154] <= Wgt_5_154;
		WeightsStore5[155] <= Wgt_5_155;
		WeightsStore5[156] <= Wgt_5_156;
		WeightsStore5[157] <= Wgt_5_157;
		WeightsStore5[158] <= Wgt_5_158;
		WeightsStore5[159] <= Wgt_5_159;
		WeightsStore5[160] <= Wgt_5_160;
		WeightsStore5[161] <= Wgt_5_161;
		WeightsStore5[162] <= Wgt_5_162;
		WeightsStore5[163] <= Wgt_5_163;
		WeightsStore5[164] <= Wgt_5_164;
		WeightsStore5[165] <= Wgt_5_165;
		WeightsStore5[166] <= Wgt_5_166;
		WeightsStore5[167] <= Wgt_5_167;
		WeightsStore5[168] <= Wgt_5_168;
		WeightsStore5[169] <= Wgt_5_169;
		WeightsStore5[170] <= Wgt_5_170;
		WeightsStore5[171] <= Wgt_5_171;
		WeightsStore5[172] <= Wgt_5_172;
		WeightsStore5[173] <= Wgt_5_173;
		WeightsStore5[174] <= Wgt_5_174;
		WeightsStore5[175] <= Wgt_5_175;
		WeightsStore5[176] <= Wgt_5_176;
		WeightsStore5[177] <= Wgt_5_177;
		WeightsStore5[178] <= Wgt_5_178;
		WeightsStore5[179] <= Wgt_5_179;
		WeightsStore5[180] <= Wgt_5_180;
		WeightsStore5[181] <= Wgt_5_181;
		WeightsStore5[182] <= Wgt_5_182;
		WeightsStore5[183] <= Wgt_5_183;
		WeightsStore5[184] <= Wgt_5_184;
		WeightsStore5[185] <= Wgt_5_185;
		WeightsStore5[186] <= Wgt_5_186;
		WeightsStore5[187] <= Wgt_5_187;
		WeightsStore5[188] <= Wgt_5_188;
		WeightsStore5[189] <= Wgt_5_189;
		WeightsStore5[190] <= Wgt_5_190;
		WeightsStore5[191] <= Wgt_5_191;
		WeightsStore5[192] <= Wgt_5_192;
		WeightsStore5[193] <= Wgt_5_193;
		WeightsStore5[194] <= Wgt_5_194;
		WeightsStore5[195] <= Wgt_5_195;
		WeightsStore5[196] <= Wgt_5_196;
		WeightsStore5[197] <= Wgt_5_197;
		WeightsStore5[198] <= Wgt_5_198;
		WeightsStore5[199] <= Wgt_5_199;
		WeightsStore5[200] <= Wgt_5_200;
		WeightsStore5[201] <= Wgt_5_201;
		WeightsStore5[202] <= Wgt_5_202;
		WeightsStore5[203] <= Wgt_5_203;
		WeightsStore5[204] <= Wgt_5_204;
		WeightsStore5[205] <= Wgt_5_205;
		WeightsStore5[206] <= Wgt_5_206;
		WeightsStore5[207] <= Wgt_5_207;
		WeightsStore5[208] <= Wgt_5_208;
		WeightsStore5[209] <= Wgt_5_209;
		WeightsStore5[210] <= Wgt_5_210;
		WeightsStore5[211] <= Wgt_5_211;
		WeightsStore5[212] <= Wgt_5_212;
		WeightsStore5[213] <= Wgt_5_213;
		WeightsStore5[214] <= Wgt_5_214;
		WeightsStore5[215] <= Wgt_5_215;
		WeightsStore5[216] <= Wgt_5_216;
		WeightsStore5[217] <= Wgt_5_217;
		WeightsStore5[218] <= Wgt_5_218;
		WeightsStore5[219] <= Wgt_5_219;
		WeightsStore5[220] <= Wgt_5_220;
		WeightsStore5[221] <= Wgt_5_221;
		WeightsStore5[222] <= Wgt_5_222;
		WeightsStore5[223] <= Wgt_5_223;
		WeightsStore5[224] <= Wgt_5_224;
		WeightsStore5[225] <= Wgt_5_225;
		WeightsStore5[226] <= Wgt_5_226;
		WeightsStore5[227] <= Wgt_5_227;
		WeightsStore5[228] <= Wgt_5_228;
		WeightsStore5[229] <= Wgt_5_229;
		WeightsStore5[230] <= Wgt_5_230;
		WeightsStore5[231] <= Wgt_5_231;
		WeightsStore5[232] <= Wgt_5_232;
		WeightsStore5[233] <= Wgt_5_233;
		WeightsStore5[234] <= Wgt_5_234;
		WeightsStore5[235] <= Wgt_5_235;
		WeightsStore5[236] <= Wgt_5_236;
		WeightsStore5[237] <= Wgt_5_237;
		WeightsStore5[238] <= Wgt_5_238;
		WeightsStore5[239] <= Wgt_5_239;
		WeightsStore5[240] <= Wgt_5_240;
		WeightsStore5[241] <= Wgt_5_241;
		WeightsStore5[242] <= Wgt_5_242;
		WeightsStore5[243] <= Wgt_5_243;
		WeightsStore5[244] <= Wgt_5_244;
		WeightsStore5[245] <= Wgt_5_245;
		WeightsStore5[246] <= Wgt_5_246;
		WeightsStore5[247] <= Wgt_5_247;
		WeightsStore5[248] <= Wgt_5_248;
		WeightsStore5[249] <= Wgt_5_249;
		WeightsStore5[250] <= Wgt_5_250;
		WeightsStore5[251] <= Wgt_5_251;
		WeightsStore5[252] <= Wgt_5_252;
		WeightsStore5[253] <= Wgt_5_253;
		WeightsStore5[254] <= Wgt_5_254;
		WeightsStore5[255] <= Wgt_5_255;
		WeightsStore5[256] <= Wgt_5_256;
		WeightsStore5[257] <= Wgt_5_257;
		WeightsStore5[258] <= Wgt_5_258;
		WeightsStore5[259] <= Wgt_5_259;
		WeightsStore5[260] <= Wgt_5_260;
		WeightsStore5[261] <= Wgt_5_261;
		WeightsStore5[262] <= Wgt_5_262;
		WeightsStore5[263] <= Wgt_5_263;
		WeightsStore5[264] <= Wgt_5_264;
		WeightsStore5[265] <= Wgt_5_265;
		WeightsStore5[266] <= Wgt_5_266;
		WeightsStore5[267] <= Wgt_5_267;
		WeightsStore5[268] <= Wgt_5_268;
		WeightsStore5[269] <= Wgt_5_269;
		WeightsStore5[270] <= Wgt_5_270;
		WeightsStore5[271] <= Wgt_5_271;
		WeightsStore5[272] <= Wgt_5_272;
		WeightsStore5[273] <= Wgt_5_273;
		WeightsStore5[274] <= Wgt_5_274;
		WeightsStore5[275] <= Wgt_5_275;
		WeightsStore5[276] <= Wgt_5_276;
		WeightsStore5[277] <= Wgt_5_277;
		WeightsStore5[278] <= Wgt_5_278;
		WeightsStore5[279] <= Wgt_5_279;
		WeightsStore5[280] <= Wgt_5_280;
		WeightsStore5[281] <= Wgt_5_281;
		WeightsStore5[282] <= Wgt_5_282;
		WeightsStore5[283] <= Wgt_5_283;
		WeightsStore5[284] <= Wgt_5_284;
		WeightsStore5[285] <= Wgt_5_285;
		WeightsStore5[286] <= Wgt_5_286;
		WeightsStore5[287] <= Wgt_5_287;
		WeightsStore5[288] <= Wgt_5_288;
		WeightsStore5[289] <= Wgt_5_289;
		WeightsStore5[290] <= Wgt_5_290;
		WeightsStore5[291] <= Wgt_5_291;
		WeightsStore5[292] <= Wgt_5_292;
		WeightsStore5[293] <= Wgt_5_293;
		WeightsStore5[294] <= Wgt_5_294;
		WeightsStore5[295] <= Wgt_5_295;
		WeightsStore5[296] <= Wgt_5_296;
		WeightsStore5[297] <= Wgt_5_297;
		WeightsStore5[298] <= Wgt_5_298;
		WeightsStore5[299] <= Wgt_5_299;
		WeightsStore5[300] <= Wgt_5_300;
		WeightsStore5[301] <= Wgt_5_301;
		WeightsStore5[302] <= Wgt_5_302;
		WeightsStore5[303] <= Wgt_5_303;
		WeightsStore5[304] <= Wgt_5_304;
		WeightsStore5[305] <= Wgt_5_305;
		WeightsStore5[306] <= Wgt_5_306;
		WeightsStore5[307] <= Wgt_5_307;
		WeightsStore5[308] <= Wgt_5_308;
		WeightsStore5[309] <= Wgt_5_309;
		WeightsStore5[310] <= Wgt_5_310;
		WeightsStore5[311] <= Wgt_5_311;
		WeightsStore5[312] <= Wgt_5_312;
		WeightsStore5[313] <= Wgt_5_313;
		WeightsStore5[314] <= Wgt_5_314;
		WeightsStore5[315] <= Wgt_5_315;
		WeightsStore5[316] <= Wgt_5_316;
		WeightsStore5[317] <= Wgt_5_317;
		WeightsStore5[318] <= Wgt_5_318;
		WeightsStore5[319] <= Wgt_5_319;
		WeightsStore5[320] <= Wgt_5_320;
		WeightsStore5[321] <= Wgt_5_321;
		WeightsStore5[322] <= Wgt_5_322;
		WeightsStore5[323] <= Wgt_5_323;
		WeightsStore5[324] <= Wgt_5_324;
		WeightsStore5[325] <= Wgt_5_325;
		WeightsStore5[326] <= Wgt_5_326;
		WeightsStore5[327] <= Wgt_5_327;
		WeightsStore5[328] <= Wgt_5_328;
		WeightsStore5[329] <= Wgt_5_329;
		WeightsStore5[330] <= Wgt_5_330;
		WeightsStore5[331] <= Wgt_5_331;
		WeightsStore5[332] <= Wgt_5_332;
		WeightsStore5[333] <= Wgt_5_333;
		WeightsStore5[334] <= Wgt_5_334;
		WeightsStore5[335] <= Wgt_5_335;
		WeightsStore5[336] <= Wgt_5_336;
		WeightsStore5[337] <= Wgt_5_337;
		WeightsStore5[338] <= Wgt_5_338;
		WeightsStore5[339] <= Wgt_5_339;
		WeightsStore5[340] <= Wgt_5_340;
		WeightsStore5[341] <= Wgt_5_341;
		WeightsStore5[342] <= Wgt_5_342;
		WeightsStore5[343] <= Wgt_5_343;
		WeightsStore5[344] <= Wgt_5_344;
		WeightsStore5[345] <= Wgt_5_345;
		WeightsStore5[346] <= Wgt_5_346;
		WeightsStore5[347] <= Wgt_5_347;
		WeightsStore5[348] <= Wgt_5_348;
		WeightsStore5[349] <= Wgt_5_349;
		WeightsStore5[350] <= Wgt_5_350;
		WeightsStore5[351] <= Wgt_5_351;
		WeightsStore5[352] <= Wgt_5_352;
		WeightsStore5[353] <= Wgt_5_353;
		WeightsStore5[354] <= Wgt_5_354;
		WeightsStore5[355] <= Wgt_5_355;
		WeightsStore5[356] <= Wgt_5_356;
		WeightsStore5[357] <= Wgt_5_357;
		WeightsStore5[358] <= Wgt_5_358;
		WeightsStore5[359] <= Wgt_5_359;
		WeightsStore5[360] <= Wgt_5_360;
		WeightsStore5[361] <= Wgt_5_361;
		WeightsStore5[362] <= Wgt_5_362;
		WeightsStore5[363] <= Wgt_5_363;
		WeightsStore5[364] <= Wgt_5_364;
		WeightsStore5[365] <= Wgt_5_365;
		WeightsStore5[366] <= Wgt_5_366;
		WeightsStore5[367] <= Wgt_5_367;
		WeightsStore5[368] <= Wgt_5_368;
		WeightsStore5[369] <= Wgt_5_369;
		WeightsStore5[370] <= Wgt_5_370;
		WeightsStore5[371] <= Wgt_5_371;
		WeightsStore5[372] <= Wgt_5_372;
		WeightsStore5[373] <= Wgt_5_373;
		WeightsStore5[374] <= Wgt_5_374;
		WeightsStore5[375] <= Wgt_5_375;
		WeightsStore5[376] <= Wgt_5_376;
		WeightsStore5[377] <= Wgt_5_377;
		WeightsStore5[378] <= Wgt_5_378;
		WeightsStore5[379] <= Wgt_5_379;
		WeightsStore5[380] <= Wgt_5_380;
		WeightsStore5[381] <= Wgt_5_381;
		WeightsStore5[382] <= Wgt_5_382;
		WeightsStore5[383] <= Wgt_5_383;
		WeightsStore5[384] <= Wgt_5_384;
		WeightsStore5[385] <= Wgt_5_385;
		WeightsStore5[386] <= Wgt_5_386;
		WeightsStore5[387] <= Wgt_5_387;
		WeightsStore5[388] <= Wgt_5_388;
		WeightsStore5[389] <= Wgt_5_389;
		WeightsStore5[390] <= Wgt_5_390;
		WeightsStore5[391] <= Wgt_5_391;
		WeightsStore5[392] <= Wgt_5_392;
		WeightsStore5[393] <= Wgt_5_393;
		WeightsStore5[394] <= Wgt_5_394;
		WeightsStore5[395] <= Wgt_5_395;
		WeightsStore5[396] <= Wgt_5_396;
		WeightsStore5[397] <= Wgt_5_397;
		WeightsStore5[398] <= Wgt_5_398;
		WeightsStore5[399] <= Wgt_5_399;
		WeightsStore5[400] <= Wgt_5_400;
		WeightsStore5[401] <= Wgt_5_401;
		WeightsStore5[402] <= Wgt_5_402;
		WeightsStore5[403] <= Wgt_5_403;
		WeightsStore5[404] <= Wgt_5_404;
		WeightsStore5[405] <= Wgt_5_405;
		WeightsStore5[406] <= Wgt_5_406;
		WeightsStore5[407] <= Wgt_5_407;
		WeightsStore5[408] <= Wgt_5_408;
		WeightsStore5[409] <= Wgt_5_409;
		WeightsStore5[410] <= Wgt_5_410;
		WeightsStore5[411] <= Wgt_5_411;
		WeightsStore5[412] <= Wgt_5_412;
		WeightsStore5[413] <= Wgt_5_413;
		WeightsStore5[414] <= Wgt_5_414;
		WeightsStore5[415] <= Wgt_5_415;
		WeightsStore5[416] <= Wgt_5_416;
		WeightsStore5[417] <= Wgt_5_417;
		WeightsStore5[418] <= Wgt_5_418;
		WeightsStore5[419] <= Wgt_5_419;
		WeightsStore5[420] <= Wgt_5_420;
		WeightsStore5[421] <= Wgt_5_421;
		WeightsStore5[422] <= Wgt_5_422;
		WeightsStore5[423] <= Wgt_5_423;
		WeightsStore5[424] <= Wgt_5_424;
		WeightsStore5[425] <= Wgt_5_425;
		WeightsStore5[426] <= Wgt_5_426;
		WeightsStore5[427] <= Wgt_5_427;
		WeightsStore5[428] <= Wgt_5_428;
		WeightsStore5[429] <= Wgt_5_429;
		WeightsStore5[430] <= Wgt_5_430;
		WeightsStore5[431] <= Wgt_5_431;
		WeightsStore5[432] <= Wgt_5_432;
		WeightsStore5[433] <= Wgt_5_433;
		WeightsStore5[434] <= Wgt_5_434;
		WeightsStore5[435] <= Wgt_5_435;
		WeightsStore5[436] <= Wgt_5_436;
		WeightsStore5[437] <= Wgt_5_437;
		WeightsStore5[438] <= Wgt_5_438;
		WeightsStore5[439] <= Wgt_5_439;
		WeightsStore5[440] <= Wgt_5_440;
		WeightsStore5[441] <= Wgt_5_441;
		WeightsStore5[442] <= Wgt_5_442;
		WeightsStore5[443] <= Wgt_5_443;
		WeightsStore5[444] <= Wgt_5_444;
		WeightsStore5[445] <= Wgt_5_445;
		WeightsStore5[446] <= Wgt_5_446;
		WeightsStore5[447] <= Wgt_5_447;
		WeightsStore5[448] <= Wgt_5_448;
		WeightsStore5[449] <= Wgt_5_449;
		WeightsStore5[450] <= Wgt_5_450;
		WeightsStore5[451] <= Wgt_5_451;
		WeightsStore5[452] <= Wgt_5_452;
		WeightsStore5[453] <= Wgt_5_453;
		WeightsStore5[454] <= Wgt_5_454;
		WeightsStore5[455] <= Wgt_5_455;
		WeightsStore5[456] <= Wgt_5_456;
		WeightsStore5[457] <= Wgt_5_457;
		WeightsStore5[458] <= Wgt_5_458;
		WeightsStore5[459] <= Wgt_5_459;
		WeightsStore5[460] <= Wgt_5_460;
		WeightsStore5[461] <= Wgt_5_461;
		WeightsStore5[462] <= Wgt_5_462;
		WeightsStore5[463] <= Wgt_5_463;
		WeightsStore5[464] <= Wgt_5_464;
		WeightsStore5[465] <= Wgt_5_465;
		WeightsStore5[466] <= Wgt_5_466;
		WeightsStore5[467] <= Wgt_5_467;
		WeightsStore5[468] <= Wgt_5_468;
		WeightsStore5[469] <= Wgt_5_469;
		WeightsStore5[470] <= Wgt_5_470;
		WeightsStore5[471] <= Wgt_5_471;
		WeightsStore5[472] <= Wgt_5_472;
		WeightsStore5[473] <= Wgt_5_473;
		WeightsStore5[474] <= Wgt_5_474;
		WeightsStore5[475] <= Wgt_5_475;
		WeightsStore5[476] <= Wgt_5_476;
		WeightsStore5[477] <= Wgt_5_477;
		WeightsStore5[478] <= Wgt_5_478;
		WeightsStore5[479] <= Wgt_5_479;
		WeightsStore5[480] <= Wgt_5_480;
		WeightsStore5[481] <= Wgt_5_481;
		WeightsStore5[482] <= Wgt_5_482;
		WeightsStore5[483] <= Wgt_5_483;
		WeightsStore5[484] <= Wgt_5_484;
		WeightsStore5[485] <= Wgt_5_485;
		WeightsStore5[486] <= Wgt_5_486;
		WeightsStore5[487] <= Wgt_5_487;
		WeightsStore5[488] <= Wgt_5_488;
		WeightsStore5[489] <= Wgt_5_489;
		WeightsStore5[490] <= Wgt_5_490;
		WeightsStore5[491] <= Wgt_5_491;
		WeightsStore5[492] <= Wgt_5_492;
		WeightsStore5[493] <= Wgt_5_493;
		WeightsStore5[494] <= Wgt_5_494;
		WeightsStore5[495] <= Wgt_5_495;
		WeightsStore5[496] <= Wgt_5_496;
		WeightsStore5[497] <= Wgt_5_497;
		WeightsStore5[498] <= Wgt_5_498;
		WeightsStore5[499] <= Wgt_5_499;
		WeightsStore5[500] <= Wgt_5_500;
		WeightsStore5[501] <= Wgt_5_501;
		WeightsStore5[502] <= Wgt_5_502;
		WeightsStore5[503] <= Wgt_5_503;
		WeightsStore5[504] <= Wgt_5_504;
		WeightsStore5[505] <= Wgt_5_505;
		WeightsStore5[506] <= Wgt_5_506;
		WeightsStore5[507] <= Wgt_5_507;
		WeightsStore5[508] <= Wgt_5_508;
		WeightsStore5[509] <= Wgt_5_509;
		WeightsStore5[510] <= Wgt_5_510;
		WeightsStore5[511] <= Wgt_5_511;
		WeightsStore5[512] <= Wgt_5_512;
		WeightsStore5[513] <= Wgt_5_513;
		WeightsStore5[514] <= Wgt_5_514;
		WeightsStore5[515] <= Wgt_5_515;
		WeightsStore5[516] <= Wgt_5_516;
		WeightsStore5[517] <= Wgt_5_517;
		WeightsStore5[518] <= Wgt_5_518;
		WeightsStore5[519] <= Wgt_5_519;
		WeightsStore5[520] <= Wgt_5_520;
		WeightsStore5[521] <= Wgt_5_521;
		WeightsStore5[522] <= Wgt_5_522;
		WeightsStore5[523] <= Wgt_5_523;
		WeightsStore5[524] <= Wgt_5_524;
		WeightsStore5[525] <= Wgt_5_525;
		WeightsStore5[526] <= Wgt_5_526;
		WeightsStore5[527] <= Wgt_5_527;
		WeightsStore5[528] <= Wgt_5_528;
		WeightsStore5[529] <= Wgt_5_529;
		WeightsStore5[530] <= Wgt_5_530;
		WeightsStore5[531] <= Wgt_5_531;
		WeightsStore5[532] <= Wgt_5_532;
		WeightsStore5[533] <= Wgt_5_533;
		WeightsStore5[534] <= Wgt_5_534;
		WeightsStore5[535] <= Wgt_5_535;
		WeightsStore5[536] <= Wgt_5_536;
		WeightsStore5[537] <= Wgt_5_537;
		WeightsStore5[538] <= Wgt_5_538;
		WeightsStore5[539] <= Wgt_5_539;
		WeightsStore5[540] <= Wgt_5_540;
		WeightsStore5[541] <= Wgt_5_541;
		WeightsStore5[542] <= Wgt_5_542;
		WeightsStore5[543] <= Wgt_5_543;
		WeightsStore5[544] <= Wgt_5_544;
		WeightsStore5[545] <= Wgt_5_545;
		WeightsStore5[546] <= Wgt_5_546;
		WeightsStore5[547] <= Wgt_5_547;
		WeightsStore5[548] <= Wgt_5_548;
		WeightsStore5[549] <= Wgt_5_549;
		WeightsStore5[550] <= Wgt_5_550;
		WeightsStore5[551] <= Wgt_5_551;
		WeightsStore5[552] <= Wgt_5_552;
		WeightsStore5[553] <= Wgt_5_553;
		WeightsStore5[554] <= Wgt_5_554;
		WeightsStore5[555] <= Wgt_5_555;
		WeightsStore5[556] <= Wgt_5_556;
		WeightsStore5[557] <= Wgt_5_557;
		WeightsStore5[558] <= Wgt_5_558;
		WeightsStore5[559] <= Wgt_5_559;
		WeightsStore5[560] <= Wgt_5_560;
		WeightsStore5[561] <= Wgt_5_561;
		WeightsStore5[562] <= Wgt_5_562;
		WeightsStore5[563] <= Wgt_5_563;
		WeightsStore5[564] <= Wgt_5_564;
		WeightsStore5[565] <= Wgt_5_565;
		WeightsStore5[566] <= Wgt_5_566;
		WeightsStore5[567] <= Wgt_5_567;
		WeightsStore5[568] <= Wgt_5_568;
		WeightsStore5[569] <= Wgt_5_569;
		WeightsStore5[570] <= Wgt_5_570;
		WeightsStore5[571] <= Wgt_5_571;
		WeightsStore5[572] <= Wgt_5_572;
		WeightsStore5[573] <= Wgt_5_573;
		WeightsStore5[574] <= Wgt_5_574;
		WeightsStore5[575] <= Wgt_5_575;
		WeightsStore5[576] <= Wgt_5_576;
		WeightsStore5[577] <= Wgt_5_577;
		WeightsStore5[578] <= Wgt_5_578;
		WeightsStore5[579] <= Wgt_5_579;
		WeightsStore5[580] <= Wgt_5_580;
		WeightsStore5[581] <= Wgt_5_581;
		WeightsStore5[582] <= Wgt_5_582;
		WeightsStore5[583] <= Wgt_5_583;
		WeightsStore5[584] <= Wgt_5_584;
		WeightsStore5[585] <= Wgt_5_585;
		WeightsStore5[586] <= Wgt_5_586;
		WeightsStore5[587] <= Wgt_5_587;
		WeightsStore5[588] <= Wgt_5_588;
		WeightsStore5[589] <= Wgt_5_589;
		WeightsStore5[590] <= Wgt_5_590;
		WeightsStore5[591] <= Wgt_5_591;
		WeightsStore5[592] <= Wgt_5_592;
		WeightsStore5[593] <= Wgt_5_593;
		WeightsStore5[594] <= Wgt_5_594;
		WeightsStore5[595] <= Wgt_5_595;
		WeightsStore5[596] <= Wgt_5_596;
		WeightsStore5[597] <= Wgt_5_597;
		WeightsStore5[598] <= Wgt_5_598;
		WeightsStore5[599] <= Wgt_5_599;
		WeightsStore5[600] <= Wgt_5_600;
		WeightsStore5[601] <= Wgt_5_601;
		WeightsStore5[602] <= Wgt_5_602;
		WeightsStore5[603] <= Wgt_5_603;
		WeightsStore5[604] <= Wgt_5_604;
		WeightsStore5[605] <= Wgt_5_605;
		WeightsStore5[606] <= Wgt_5_606;
		WeightsStore5[607] <= Wgt_5_607;
		WeightsStore5[608] <= Wgt_5_608;
		WeightsStore5[609] <= Wgt_5_609;
		WeightsStore5[610] <= Wgt_5_610;
		WeightsStore5[611] <= Wgt_5_611;
		WeightsStore5[612] <= Wgt_5_612;
		WeightsStore5[613] <= Wgt_5_613;
		WeightsStore5[614] <= Wgt_5_614;
		WeightsStore5[615] <= Wgt_5_615;
		WeightsStore5[616] <= Wgt_5_616;
		WeightsStore5[617] <= Wgt_5_617;
		WeightsStore5[618] <= Wgt_5_618;
		WeightsStore5[619] <= Wgt_5_619;
		WeightsStore5[620] <= Wgt_5_620;
		WeightsStore5[621] <= Wgt_5_621;
		WeightsStore5[622] <= Wgt_5_622;
		WeightsStore5[623] <= Wgt_5_623;
		WeightsStore5[624] <= Wgt_5_624;
		WeightsStore5[625] <= Wgt_5_625;
		WeightsStore5[626] <= Wgt_5_626;
		WeightsStore5[627] <= Wgt_5_627;
		WeightsStore5[628] <= Wgt_5_628;
		WeightsStore5[629] <= Wgt_5_629;
		WeightsStore5[630] <= Wgt_5_630;
		WeightsStore5[631] <= Wgt_5_631;
		WeightsStore5[632] <= Wgt_5_632;
		WeightsStore5[633] <= Wgt_5_633;
		WeightsStore5[634] <= Wgt_5_634;
		WeightsStore5[635] <= Wgt_5_635;
		WeightsStore5[636] <= Wgt_5_636;
		WeightsStore5[637] <= Wgt_5_637;
		WeightsStore5[638] <= Wgt_5_638;
		WeightsStore5[639] <= Wgt_5_639;
		WeightsStore5[640] <= Wgt_5_640;
		WeightsStore5[641] <= Wgt_5_641;
		WeightsStore5[642] <= Wgt_5_642;
		WeightsStore5[643] <= Wgt_5_643;
		WeightsStore5[644] <= Wgt_5_644;
		WeightsStore5[645] <= Wgt_5_645;
		WeightsStore5[646] <= Wgt_5_646;
		WeightsStore5[647] <= Wgt_5_647;
		WeightsStore5[648] <= Wgt_5_648;
		WeightsStore5[649] <= Wgt_5_649;
		WeightsStore5[650] <= Wgt_5_650;
		WeightsStore5[651] <= Wgt_5_651;
		WeightsStore5[652] <= Wgt_5_652;
		WeightsStore5[653] <= Wgt_5_653;
		WeightsStore5[654] <= Wgt_5_654;
		WeightsStore5[655] <= Wgt_5_655;
		WeightsStore5[656] <= Wgt_5_656;
		WeightsStore5[657] <= Wgt_5_657;
		WeightsStore5[658] <= Wgt_5_658;
		WeightsStore5[659] <= Wgt_5_659;
		WeightsStore5[660] <= Wgt_5_660;
		WeightsStore5[661] <= Wgt_5_661;
		WeightsStore5[662] <= Wgt_5_662;
		WeightsStore5[663] <= Wgt_5_663;
		WeightsStore5[664] <= Wgt_5_664;
		WeightsStore5[665] <= Wgt_5_665;
		WeightsStore5[666] <= Wgt_5_666;
		WeightsStore5[667] <= Wgt_5_667;
		WeightsStore5[668] <= Wgt_5_668;
		WeightsStore5[669] <= Wgt_5_669;
		WeightsStore5[670] <= Wgt_5_670;
		WeightsStore5[671] <= Wgt_5_671;
		WeightsStore5[672] <= Wgt_5_672;
		WeightsStore5[673] <= Wgt_5_673;
		WeightsStore5[674] <= Wgt_5_674;
		WeightsStore5[675] <= Wgt_5_675;
		WeightsStore5[676] <= Wgt_5_676;
		WeightsStore5[677] <= Wgt_5_677;
		WeightsStore5[678] <= Wgt_5_678;
		WeightsStore5[679] <= Wgt_5_679;
		WeightsStore5[680] <= Wgt_5_680;
		WeightsStore5[681] <= Wgt_5_681;
		WeightsStore5[682] <= Wgt_5_682;
		WeightsStore5[683] <= Wgt_5_683;
		WeightsStore5[684] <= Wgt_5_684;
		WeightsStore5[685] <= Wgt_5_685;
		WeightsStore5[686] <= Wgt_5_686;
		WeightsStore5[687] <= Wgt_5_687;
		WeightsStore5[688] <= Wgt_5_688;
		WeightsStore5[689] <= Wgt_5_689;
		WeightsStore5[690] <= Wgt_5_690;
		WeightsStore5[691] <= Wgt_5_691;
		WeightsStore5[692] <= Wgt_5_692;
		WeightsStore5[693] <= Wgt_5_693;
		WeightsStore5[694] <= Wgt_5_694;
		WeightsStore5[695] <= Wgt_5_695;
		WeightsStore5[696] <= Wgt_5_696;
		WeightsStore5[697] <= Wgt_5_697;
		WeightsStore5[698] <= Wgt_5_698;
		WeightsStore5[699] <= Wgt_5_699;
		WeightsStore5[700] <= Wgt_5_700;
		WeightsStore5[701] <= Wgt_5_701;
		WeightsStore5[702] <= Wgt_5_702;
		WeightsStore5[703] <= Wgt_5_703;
		WeightsStore5[704] <= Wgt_5_704;
		WeightsStore5[705] <= Wgt_5_705;
		WeightsStore5[706] <= Wgt_5_706;
		WeightsStore5[707] <= Wgt_5_707;
		WeightsStore5[708] <= Wgt_5_708;
		WeightsStore5[709] <= Wgt_5_709;
		WeightsStore5[710] <= Wgt_5_710;
		WeightsStore5[711] <= Wgt_5_711;
		WeightsStore5[712] <= Wgt_5_712;
		WeightsStore5[713] <= Wgt_5_713;
		WeightsStore5[714] <= Wgt_5_714;
		WeightsStore5[715] <= Wgt_5_715;
		WeightsStore5[716] <= Wgt_5_716;
		WeightsStore5[717] <= Wgt_5_717;
		WeightsStore5[718] <= Wgt_5_718;
		WeightsStore5[719] <= Wgt_5_719;
		WeightsStore5[720] <= Wgt_5_720;
		WeightsStore5[721] <= Wgt_5_721;
		WeightsStore5[722] <= Wgt_5_722;
		WeightsStore5[723] <= Wgt_5_723;
		WeightsStore5[724] <= Wgt_5_724;
		WeightsStore5[725] <= Wgt_5_725;
		WeightsStore5[726] <= Wgt_5_726;
		WeightsStore5[727] <= Wgt_5_727;
		WeightsStore5[728] <= Wgt_5_728;
		WeightsStore5[729] <= Wgt_5_729;
		WeightsStore5[730] <= Wgt_5_730;
		WeightsStore5[731] <= Wgt_5_731;
		WeightsStore5[732] <= Wgt_5_732;
		WeightsStore5[733] <= Wgt_5_733;
		WeightsStore5[734] <= Wgt_5_734;
		WeightsStore5[735] <= Wgt_5_735;
		WeightsStore5[736] <= Wgt_5_736;
		WeightsStore5[737] <= Wgt_5_737;
		WeightsStore5[738] <= Wgt_5_738;
		WeightsStore5[739] <= Wgt_5_739;
		WeightsStore5[740] <= Wgt_5_740;
		WeightsStore5[741] <= Wgt_5_741;
		WeightsStore5[742] <= Wgt_5_742;
		WeightsStore5[743] <= Wgt_5_743;
		WeightsStore5[744] <= Wgt_5_744;
		WeightsStore5[745] <= Wgt_5_745;
		WeightsStore5[746] <= Wgt_5_746;
		WeightsStore5[747] <= Wgt_5_747;
		WeightsStore5[748] <= Wgt_5_748;
		WeightsStore5[749] <= Wgt_5_749;
		WeightsStore5[750] <= Wgt_5_750;
		WeightsStore5[751] <= Wgt_5_751;
		WeightsStore5[752] <= Wgt_5_752;
		WeightsStore5[753] <= Wgt_5_753;
		WeightsStore5[754] <= Wgt_5_754;
		WeightsStore5[755] <= Wgt_5_755;
		WeightsStore5[756] <= Wgt_5_756;
		WeightsStore5[757] <= Wgt_5_757;
		WeightsStore5[758] <= Wgt_5_758;
		WeightsStore5[759] <= Wgt_5_759;
		WeightsStore5[760] <= Wgt_5_760;
		WeightsStore5[761] <= Wgt_5_761;
		WeightsStore5[762] <= Wgt_5_762;
		WeightsStore5[763] <= Wgt_5_763;
		WeightsStore5[764] <= Wgt_5_764;
		WeightsStore5[765] <= Wgt_5_765;
		WeightsStore5[766] <= Wgt_5_766;
		WeightsStore5[767] <= Wgt_5_767;
		WeightsStore5[768] <= Wgt_5_768;
		WeightsStore5[769] <= Wgt_5_769;
		WeightsStore5[770] <= Wgt_5_770;
		WeightsStore5[771] <= Wgt_5_771;
		WeightsStore5[772] <= Wgt_5_772;
		WeightsStore5[773] <= Wgt_5_773;
		WeightsStore5[774] <= Wgt_5_774;
		WeightsStore5[775] <= Wgt_5_775;
		WeightsStore5[776] <= Wgt_5_776;
		WeightsStore5[777] <= Wgt_5_777;
		WeightsStore5[778] <= Wgt_5_778;
		WeightsStore5[779] <= Wgt_5_779;
		WeightsStore5[780] <= Wgt_5_780;
		WeightsStore5[781] <= Wgt_5_781;
		WeightsStore5[782] <= Wgt_5_782;
		WeightsStore5[783] <= Wgt_5_783;
		WeightsStore5[784] <= Wgt_5_784;
		WeightsStore6[0] <= Wgt_6_0;
		WeightsStore6[1] <= Wgt_6_1;
		WeightsStore6[2] <= Wgt_6_2;
		WeightsStore6[3] <= Wgt_6_3;
		WeightsStore6[4] <= Wgt_6_4;
		WeightsStore6[5] <= Wgt_6_5;
		WeightsStore6[6] <= Wgt_6_6;
		WeightsStore6[7] <= Wgt_6_7;
		WeightsStore6[8] <= Wgt_6_8;
		WeightsStore6[9] <= Wgt_6_9;
		WeightsStore6[10] <= Wgt_6_10;
		WeightsStore6[11] <= Wgt_6_11;
		WeightsStore6[12] <= Wgt_6_12;
		WeightsStore6[13] <= Wgt_6_13;
		WeightsStore6[14] <= Wgt_6_14;
		WeightsStore6[15] <= Wgt_6_15;
		WeightsStore6[16] <= Wgt_6_16;
		WeightsStore6[17] <= Wgt_6_17;
		WeightsStore6[18] <= Wgt_6_18;
		WeightsStore6[19] <= Wgt_6_19;
		WeightsStore6[20] <= Wgt_6_20;
		WeightsStore6[21] <= Wgt_6_21;
		WeightsStore6[22] <= Wgt_6_22;
		WeightsStore6[23] <= Wgt_6_23;
		WeightsStore6[24] <= Wgt_6_24;
		WeightsStore6[25] <= Wgt_6_25;
		WeightsStore6[26] <= Wgt_6_26;
		WeightsStore6[27] <= Wgt_6_27;
		WeightsStore6[28] <= Wgt_6_28;
		WeightsStore6[29] <= Wgt_6_29;
		WeightsStore6[30] <= Wgt_6_30;
		WeightsStore6[31] <= Wgt_6_31;
		WeightsStore6[32] <= Wgt_6_32;
		WeightsStore6[33] <= Wgt_6_33;
		WeightsStore6[34] <= Wgt_6_34;
		WeightsStore6[35] <= Wgt_6_35;
		WeightsStore6[36] <= Wgt_6_36;
		WeightsStore6[37] <= Wgt_6_37;
		WeightsStore6[38] <= Wgt_6_38;
		WeightsStore6[39] <= Wgt_6_39;
		WeightsStore6[40] <= Wgt_6_40;
		WeightsStore6[41] <= Wgt_6_41;
		WeightsStore6[42] <= Wgt_6_42;
		WeightsStore6[43] <= Wgt_6_43;
		WeightsStore6[44] <= Wgt_6_44;
		WeightsStore6[45] <= Wgt_6_45;
		WeightsStore6[46] <= Wgt_6_46;
		WeightsStore6[47] <= Wgt_6_47;
		WeightsStore6[48] <= Wgt_6_48;
		WeightsStore6[49] <= Wgt_6_49;
		WeightsStore6[50] <= Wgt_6_50;
		WeightsStore6[51] <= Wgt_6_51;
		WeightsStore6[52] <= Wgt_6_52;
		WeightsStore6[53] <= Wgt_6_53;
		WeightsStore6[54] <= Wgt_6_54;
		WeightsStore6[55] <= Wgt_6_55;
		WeightsStore6[56] <= Wgt_6_56;
		WeightsStore6[57] <= Wgt_6_57;
		WeightsStore6[58] <= Wgt_6_58;
		WeightsStore6[59] <= Wgt_6_59;
		WeightsStore6[60] <= Wgt_6_60;
		WeightsStore6[61] <= Wgt_6_61;
		WeightsStore6[62] <= Wgt_6_62;
		WeightsStore6[63] <= Wgt_6_63;
		WeightsStore6[64] <= Wgt_6_64;
		WeightsStore6[65] <= Wgt_6_65;
		WeightsStore6[66] <= Wgt_6_66;
		WeightsStore6[67] <= Wgt_6_67;
		WeightsStore6[68] <= Wgt_6_68;
		WeightsStore6[69] <= Wgt_6_69;
		WeightsStore6[70] <= Wgt_6_70;
		WeightsStore6[71] <= Wgt_6_71;
		WeightsStore6[72] <= Wgt_6_72;
		WeightsStore6[73] <= Wgt_6_73;
		WeightsStore6[74] <= Wgt_6_74;
		WeightsStore6[75] <= Wgt_6_75;
		WeightsStore6[76] <= Wgt_6_76;
		WeightsStore6[77] <= Wgt_6_77;
		WeightsStore6[78] <= Wgt_6_78;
		WeightsStore6[79] <= Wgt_6_79;
		WeightsStore6[80] <= Wgt_6_80;
		WeightsStore6[81] <= Wgt_6_81;
		WeightsStore6[82] <= Wgt_6_82;
		WeightsStore6[83] <= Wgt_6_83;
		WeightsStore6[84] <= Wgt_6_84;
		WeightsStore6[85] <= Wgt_6_85;
		WeightsStore6[86] <= Wgt_6_86;
		WeightsStore6[87] <= Wgt_6_87;
		WeightsStore6[88] <= Wgt_6_88;
		WeightsStore6[89] <= Wgt_6_89;
		WeightsStore6[90] <= Wgt_6_90;
		WeightsStore6[91] <= Wgt_6_91;
		WeightsStore6[92] <= Wgt_6_92;
		WeightsStore6[93] <= Wgt_6_93;
		WeightsStore6[94] <= Wgt_6_94;
		WeightsStore6[95] <= Wgt_6_95;
		WeightsStore6[96] <= Wgt_6_96;
		WeightsStore6[97] <= Wgt_6_97;
		WeightsStore6[98] <= Wgt_6_98;
		WeightsStore6[99] <= Wgt_6_99;
		WeightsStore6[100] <= Wgt_6_100;
		WeightsStore6[101] <= Wgt_6_101;
		WeightsStore6[102] <= Wgt_6_102;
		WeightsStore6[103] <= Wgt_6_103;
		WeightsStore6[104] <= Wgt_6_104;
		WeightsStore6[105] <= Wgt_6_105;
		WeightsStore6[106] <= Wgt_6_106;
		WeightsStore6[107] <= Wgt_6_107;
		WeightsStore6[108] <= Wgt_6_108;
		WeightsStore6[109] <= Wgt_6_109;
		WeightsStore6[110] <= Wgt_6_110;
		WeightsStore6[111] <= Wgt_6_111;
		WeightsStore6[112] <= Wgt_6_112;
		WeightsStore6[113] <= Wgt_6_113;
		WeightsStore6[114] <= Wgt_6_114;
		WeightsStore6[115] <= Wgt_6_115;
		WeightsStore6[116] <= Wgt_6_116;
		WeightsStore6[117] <= Wgt_6_117;
		WeightsStore6[118] <= Wgt_6_118;
		WeightsStore6[119] <= Wgt_6_119;
		WeightsStore6[120] <= Wgt_6_120;
		WeightsStore6[121] <= Wgt_6_121;
		WeightsStore6[122] <= Wgt_6_122;
		WeightsStore6[123] <= Wgt_6_123;
		WeightsStore6[124] <= Wgt_6_124;
		WeightsStore6[125] <= Wgt_6_125;
		WeightsStore6[126] <= Wgt_6_126;
		WeightsStore6[127] <= Wgt_6_127;
		WeightsStore6[128] <= Wgt_6_128;
		WeightsStore6[129] <= Wgt_6_129;
		WeightsStore6[130] <= Wgt_6_130;
		WeightsStore6[131] <= Wgt_6_131;
		WeightsStore6[132] <= Wgt_6_132;
		WeightsStore6[133] <= Wgt_6_133;
		WeightsStore6[134] <= Wgt_6_134;
		WeightsStore6[135] <= Wgt_6_135;
		WeightsStore6[136] <= Wgt_6_136;
		WeightsStore6[137] <= Wgt_6_137;
		WeightsStore6[138] <= Wgt_6_138;
		WeightsStore6[139] <= Wgt_6_139;
		WeightsStore6[140] <= Wgt_6_140;
		WeightsStore6[141] <= Wgt_6_141;
		WeightsStore6[142] <= Wgt_6_142;
		WeightsStore6[143] <= Wgt_6_143;
		WeightsStore6[144] <= Wgt_6_144;
		WeightsStore6[145] <= Wgt_6_145;
		WeightsStore6[146] <= Wgt_6_146;
		WeightsStore6[147] <= Wgt_6_147;
		WeightsStore6[148] <= Wgt_6_148;
		WeightsStore6[149] <= Wgt_6_149;
		WeightsStore6[150] <= Wgt_6_150;
		WeightsStore6[151] <= Wgt_6_151;
		WeightsStore6[152] <= Wgt_6_152;
		WeightsStore6[153] <= Wgt_6_153;
		WeightsStore6[154] <= Wgt_6_154;
		WeightsStore6[155] <= Wgt_6_155;
		WeightsStore6[156] <= Wgt_6_156;
		WeightsStore6[157] <= Wgt_6_157;
		WeightsStore6[158] <= Wgt_6_158;
		WeightsStore6[159] <= Wgt_6_159;
		WeightsStore6[160] <= Wgt_6_160;
		WeightsStore6[161] <= Wgt_6_161;
		WeightsStore6[162] <= Wgt_6_162;
		WeightsStore6[163] <= Wgt_6_163;
		WeightsStore6[164] <= Wgt_6_164;
		WeightsStore6[165] <= Wgt_6_165;
		WeightsStore6[166] <= Wgt_6_166;
		WeightsStore6[167] <= Wgt_6_167;
		WeightsStore6[168] <= Wgt_6_168;
		WeightsStore6[169] <= Wgt_6_169;
		WeightsStore6[170] <= Wgt_6_170;
		WeightsStore6[171] <= Wgt_6_171;
		WeightsStore6[172] <= Wgt_6_172;
		WeightsStore6[173] <= Wgt_6_173;
		WeightsStore6[174] <= Wgt_6_174;
		WeightsStore6[175] <= Wgt_6_175;
		WeightsStore6[176] <= Wgt_6_176;
		WeightsStore6[177] <= Wgt_6_177;
		WeightsStore6[178] <= Wgt_6_178;
		WeightsStore6[179] <= Wgt_6_179;
		WeightsStore6[180] <= Wgt_6_180;
		WeightsStore6[181] <= Wgt_6_181;
		WeightsStore6[182] <= Wgt_6_182;
		WeightsStore6[183] <= Wgt_6_183;
		WeightsStore6[184] <= Wgt_6_184;
		WeightsStore6[185] <= Wgt_6_185;
		WeightsStore6[186] <= Wgt_6_186;
		WeightsStore6[187] <= Wgt_6_187;
		WeightsStore6[188] <= Wgt_6_188;
		WeightsStore6[189] <= Wgt_6_189;
		WeightsStore6[190] <= Wgt_6_190;
		WeightsStore6[191] <= Wgt_6_191;
		WeightsStore6[192] <= Wgt_6_192;
		WeightsStore6[193] <= Wgt_6_193;
		WeightsStore6[194] <= Wgt_6_194;
		WeightsStore6[195] <= Wgt_6_195;
		WeightsStore6[196] <= Wgt_6_196;
		WeightsStore6[197] <= Wgt_6_197;
		WeightsStore6[198] <= Wgt_6_198;
		WeightsStore6[199] <= Wgt_6_199;
		WeightsStore6[200] <= Wgt_6_200;
		WeightsStore6[201] <= Wgt_6_201;
		WeightsStore6[202] <= Wgt_6_202;
		WeightsStore6[203] <= Wgt_6_203;
		WeightsStore6[204] <= Wgt_6_204;
		WeightsStore6[205] <= Wgt_6_205;
		WeightsStore6[206] <= Wgt_6_206;
		WeightsStore6[207] <= Wgt_6_207;
		WeightsStore6[208] <= Wgt_6_208;
		WeightsStore6[209] <= Wgt_6_209;
		WeightsStore6[210] <= Wgt_6_210;
		WeightsStore6[211] <= Wgt_6_211;
		WeightsStore6[212] <= Wgt_6_212;
		WeightsStore6[213] <= Wgt_6_213;
		WeightsStore6[214] <= Wgt_6_214;
		WeightsStore6[215] <= Wgt_6_215;
		WeightsStore6[216] <= Wgt_6_216;
		WeightsStore6[217] <= Wgt_6_217;
		WeightsStore6[218] <= Wgt_6_218;
		WeightsStore6[219] <= Wgt_6_219;
		WeightsStore6[220] <= Wgt_6_220;
		WeightsStore6[221] <= Wgt_6_221;
		WeightsStore6[222] <= Wgt_6_222;
		WeightsStore6[223] <= Wgt_6_223;
		WeightsStore6[224] <= Wgt_6_224;
		WeightsStore6[225] <= Wgt_6_225;
		WeightsStore6[226] <= Wgt_6_226;
		WeightsStore6[227] <= Wgt_6_227;
		WeightsStore6[228] <= Wgt_6_228;
		WeightsStore6[229] <= Wgt_6_229;
		WeightsStore6[230] <= Wgt_6_230;
		WeightsStore6[231] <= Wgt_6_231;
		WeightsStore6[232] <= Wgt_6_232;
		WeightsStore6[233] <= Wgt_6_233;
		WeightsStore6[234] <= Wgt_6_234;
		WeightsStore6[235] <= Wgt_6_235;
		WeightsStore6[236] <= Wgt_6_236;
		WeightsStore6[237] <= Wgt_6_237;
		WeightsStore6[238] <= Wgt_6_238;
		WeightsStore6[239] <= Wgt_6_239;
		WeightsStore6[240] <= Wgt_6_240;
		WeightsStore6[241] <= Wgt_6_241;
		WeightsStore6[242] <= Wgt_6_242;
		WeightsStore6[243] <= Wgt_6_243;
		WeightsStore6[244] <= Wgt_6_244;
		WeightsStore6[245] <= Wgt_6_245;
		WeightsStore6[246] <= Wgt_6_246;
		WeightsStore6[247] <= Wgt_6_247;
		WeightsStore6[248] <= Wgt_6_248;
		WeightsStore6[249] <= Wgt_6_249;
		WeightsStore6[250] <= Wgt_6_250;
		WeightsStore6[251] <= Wgt_6_251;
		WeightsStore6[252] <= Wgt_6_252;
		WeightsStore6[253] <= Wgt_6_253;
		WeightsStore6[254] <= Wgt_6_254;
		WeightsStore6[255] <= Wgt_6_255;
		WeightsStore6[256] <= Wgt_6_256;
		WeightsStore6[257] <= Wgt_6_257;
		WeightsStore6[258] <= Wgt_6_258;
		WeightsStore6[259] <= Wgt_6_259;
		WeightsStore6[260] <= Wgt_6_260;
		WeightsStore6[261] <= Wgt_6_261;
		WeightsStore6[262] <= Wgt_6_262;
		WeightsStore6[263] <= Wgt_6_263;
		WeightsStore6[264] <= Wgt_6_264;
		WeightsStore6[265] <= Wgt_6_265;
		WeightsStore6[266] <= Wgt_6_266;
		WeightsStore6[267] <= Wgt_6_267;
		WeightsStore6[268] <= Wgt_6_268;
		WeightsStore6[269] <= Wgt_6_269;
		WeightsStore6[270] <= Wgt_6_270;
		WeightsStore6[271] <= Wgt_6_271;
		WeightsStore6[272] <= Wgt_6_272;
		WeightsStore6[273] <= Wgt_6_273;
		WeightsStore6[274] <= Wgt_6_274;
		WeightsStore6[275] <= Wgt_6_275;
		WeightsStore6[276] <= Wgt_6_276;
		WeightsStore6[277] <= Wgt_6_277;
		WeightsStore6[278] <= Wgt_6_278;
		WeightsStore6[279] <= Wgt_6_279;
		WeightsStore6[280] <= Wgt_6_280;
		WeightsStore6[281] <= Wgt_6_281;
		WeightsStore6[282] <= Wgt_6_282;
		WeightsStore6[283] <= Wgt_6_283;
		WeightsStore6[284] <= Wgt_6_284;
		WeightsStore6[285] <= Wgt_6_285;
		WeightsStore6[286] <= Wgt_6_286;
		WeightsStore6[287] <= Wgt_6_287;
		WeightsStore6[288] <= Wgt_6_288;
		WeightsStore6[289] <= Wgt_6_289;
		WeightsStore6[290] <= Wgt_6_290;
		WeightsStore6[291] <= Wgt_6_291;
		WeightsStore6[292] <= Wgt_6_292;
		WeightsStore6[293] <= Wgt_6_293;
		WeightsStore6[294] <= Wgt_6_294;
		WeightsStore6[295] <= Wgt_6_295;
		WeightsStore6[296] <= Wgt_6_296;
		WeightsStore6[297] <= Wgt_6_297;
		WeightsStore6[298] <= Wgt_6_298;
		WeightsStore6[299] <= Wgt_6_299;
		WeightsStore6[300] <= Wgt_6_300;
		WeightsStore6[301] <= Wgt_6_301;
		WeightsStore6[302] <= Wgt_6_302;
		WeightsStore6[303] <= Wgt_6_303;
		WeightsStore6[304] <= Wgt_6_304;
		WeightsStore6[305] <= Wgt_6_305;
		WeightsStore6[306] <= Wgt_6_306;
		WeightsStore6[307] <= Wgt_6_307;
		WeightsStore6[308] <= Wgt_6_308;
		WeightsStore6[309] <= Wgt_6_309;
		WeightsStore6[310] <= Wgt_6_310;
		WeightsStore6[311] <= Wgt_6_311;
		WeightsStore6[312] <= Wgt_6_312;
		WeightsStore6[313] <= Wgt_6_313;
		WeightsStore6[314] <= Wgt_6_314;
		WeightsStore6[315] <= Wgt_6_315;
		WeightsStore6[316] <= Wgt_6_316;
		WeightsStore6[317] <= Wgt_6_317;
		WeightsStore6[318] <= Wgt_6_318;
		WeightsStore6[319] <= Wgt_6_319;
		WeightsStore6[320] <= Wgt_6_320;
		WeightsStore6[321] <= Wgt_6_321;
		WeightsStore6[322] <= Wgt_6_322;
		WeightsStore6[323] <= Wgt_6_323;
		WeightsStore6[324] <= Wgt_6_324;
		WeightsStore6[325] <= Wgt_6_325;
		WeightsStore6[326] <= Wgt_6_326;
		WeightsStore6[327] <= Wgt_6_327;
		WeightsStore6[328] <= Wgt_6_328;
		WeightsStore6[329] <= Wgt_6_329;
		WeightsStore6[330] <= Wgt_6_330;
		WeightsStore6[331] <= Wgt_6_331;
		WeightsStore6[332] <= Wgt_6_332;
		WeightsStore6[333] <= Wgt_6_333;
		WeightsStore6[334] <= Wgt_6_334;
		WeightsStore6[335] <= Wgt_6_335;
		WeightsStore6[336] <= Wgt_6_336;
		WeightsStore6[337] <= Wgt_6_337;
		WeightsStore6[338] <= Wgt_6_338;
		WeightsStore6[339] <= Wgt_6_339;
		WeightsStore6[340] <= Wgt_6_340;
		WeightsStore6[341] <= Wgt_6_341;
		WeightsStore6[342] <= Wgt_6_342;
		WeightsStore6[343] <= Wgt_6_343;
		WeightsStore6[344] <= Wgt_6_344;
		WeightsStore6[345] <= Wgt_6_345;
		WeightsStore6[346] <= Wgt_6_346;
		WeightsStore6[347] <= Wgt_6_347;
		WeightsStore6[348] <= Wgt_6_348;
		WeightsStore6[349] <= Wgt_6_349;
		WeightsStore6[350] <= Wgt_6_350;
		WeightsStore6[351] <= Wgt_6_351;
		WeightsStore6[352] <= Wgt_6_352;
		WeightsStore6[353] <= Wgt_6_353;
		WeightsStore6[354] <= Wgt_6_354;
		WeightsStore6[355] <= Wgt_6_355;
		WeightsStore6[356] <= Wgt_6_356;
		WeightsStore6[357] <= Wgt_6_357;
		WeightsStore6[358] <= Wgt_6_358;
		WeightsStore6[359] <= Wgt_6_359;
		WeightsStore6[360] <= Wgt_6_360;
		WeightsStore6[361] <= Wgt_6_361;
		WeightsStore6[362] <= Wgt_6_362;
		WeightsStore6[363] <= Wgt_6_363;
		WeightsStore6[364] <= Wgt_6_364;
		WeightsStore6[365] <= Wgt_6_365;
		WeightsStore6[366] <= Wgt_6_366;
		WeightsStore6[367] <= Wgt_6_367;
		WeightsStore6[368] <= Wgt_6_368;
		WeightsStore6[369] <= Wgt_6_369;
		WeightsStore6[370] <= Wgt_6_370;
		WeightsStore6[371] <= Wgt_6_371;
		WeightsStore6[372] <= Wgt_6_372;
		WeightsStore6[373] <= Wgt_6_373;
		WeightsStore6[374] <= Wgt_6_374;
		WeightsStore6[375] <= Wgt_6_375;
		WeightsStore6[376] <= Wgt_6_376;
		WeightsStore6[377] <= Wgt_6_377;
		WeightsStore6[378] <= Wgt_6_378;
		WeightsStore6[379] <= Wgt_6_379;
		WeightsStore6[380] <= Wgt_6_380;
		WeightsStore6[381] <= Wgt_6_381;
		WeightsStore6[382] <= Wgt_6_382;
		WeightsStore6[383] <= Wgt_6_383;
		WeightsStore6[384] <= Wgt_6_384;
		WeightsStore6[385] <= Wgt_6_385;
		WeightsStore6[386] <= Wgt_6_386;
		WeightsStore6[387] <= Wgt_6_387;
		WeightsStore6[388] <= Wgt_6_388;
		WeightsStore6[389] <= Wgt_6_389;
		WeightsStore6[390] <= Wgt_6_390;
		WeightsStore6[391] <= Wgt_6_391;
		WeightsStore6[392] <= Wgt_6_392;
		WeightsStore6[393] <= Wgt_6_393;
		WeightsStore6[394] <= Wgt_6_394;
		WeightsStore6[395] <= Wgt_6_395;
		WeightsStore6[396] <= Wgt_6_396;
		WeightsStore6[397] <= Wgt_6_397;
		WeightsStore6[398] <= Wgt_6_398;
		WeightsStore6[399] <= Wgt_6_399;
		WeightsStore6[400] <= Wgt_6_400;
		WeightsStore6[401] <= Wgt_6_401;
		WeightsStore6[402] <= Wgt_6_402;
		WeightsStore6[403] <= Wgt_6_403;
		WeightsStore6[404] <= Wgt_6_404;
		WeightsStore6[405] <= Wgt_6_405;
		WeightsStore6[406] <= Wgt_6_406;
		WeightsStore6[407] <= Wgt_6_407;
		WeightsStore6[408] <= Wgt_6_408;
		WeightsStore6[409] <= Wgt_6_409;
		WeightsStore6[410] <= Wgt_6_410;
		WeightsStore6[411] <= Wgt_6_411;
		WeightsStore6[412] <= Wgt_6_412;
		WeightsStore6[413] <= Wgt_6_413;
		WeightsStore6[414] <= Wgt_6_414;
		WeightsStore6[415] <= Wgt_6_415;
		WeightsStore6[416] <= Wgt_6_416;
		WeightsStore6[417] <= Wgt_6_417;
		WeightsStore6[418] <= Wgt_6_418;
		WeightsStore6[419] <= Wgt_6_419;
		WeightsStore6[420] <= Wgt_6_420;
		WeightsStore6[421] <= Wgt_6_421;
		WeightsStore6[422] <= Wgt_6_422;
		WeightsStore6[423] <= Wgt_6_423;
		WeightsStore6[424] <= Wgt_6_424;
		WeightsStore6[425] <= Wgt_6_425;
		WeightsStore6[426] <= Wgt_6_426;
		WeightsStore6[427] <= Wgt_6_427;
		WeightsStore6[428] <= Wgt_6_428;
		WeightsStore6[429] <= Wgt_6_429;
		WeightsStore6[430] <= Wgt_6_430;
		WeightsStore6[431] <= Wgt_6_431;
		WeightsStore6[432] <= Wgt_6_432;
		WeightsStore6[433] <= Wgt_6_433;
		WeightsStore6[434] <= Wgt_6_434;
		WeightsStore6[435] <= Wgt_6_435;
		WeightsStore6[436] <= Wgt_6_436;
		WeightsStore6[437] <= Wgt_6_437;
		WeightsStore6[438] <= Wgt_6_438;
		WeightsStore6[439] <= Wgt_6_439;
		WeightsStore6[440] <= Wgt_6_440;
		WeightsStore6[441] <= Wgt_6_441;
		WeightsStore6[442] <= Wgt_6_442;
		WeightsStore6[443] <= Wgt_6_443;
		WeightsStore6[444] <= Wgt_6_444;
		WeightsStore6[445] <= Wgt_6_445;
		WeightsStore6[446] <= Wgt_6_446;
		WeightsStore6[447] <= Wgt_6_447;
		WeightsStore6[448] <= Wgt_6_448;
		WeightsStore6[449] <= Wgt_6_449;
		WeightsStore6[450] <= Wgt_6_450;
		WeightsStore6[451] <= Wgt_6_451;
		WeightsStore6[452] <= Wgt_6_452;
		WeightsStore6[453] <= Wgt_6_453;
		WeightsStore6[454] <= Wgt_6_454;
		WeightsStore6[455] <= Wgt_6_455;
		WeightsStore6[456] <= Wgt_6_456;
		WeightsStore6[457] <= Wgt_6_457;
		WeightsStore6[458] <= Wgt_6_458;
		WeightsStore6[459] <= Wgt_6_459;
		WeightsStore6[460] <= Wgt_6_460;
		WeightsStore6[461] <= Wgt_6_461;
		WeightsStore6[462] <= Wgt_6_462;
		WeightsStore6[463] <= Wgt_6_463;
		WeightsStore6[464] <= Wgt_6_464;
		WeightsStore6[465] <= Wgt_6_465;
		WeightsStore6[466] <= Wgt_6_466;
		WeightsStore6[467] <= Wgt_6_467;
		WeightsStore6[468] <= Wgt_6_468;
		WeightsStore6[469] <= Wgt_6_469;
		WeightsStore6[470] <= Wgt_6_470;
		WeightsStore6[471] <= Wgt_6_471;
		WeightsStore6[472] <= Wgt_6_472;
		WeightsStore6[473] <= Wgt_6_473;
		WeightsStore6[474] <= Wgt_6_474;
		WeightsStore6[475] <= Wgt_6_475;
		WeightsStore6[476] <= Wgt_6_476;
		WeightsStore6[477] <= Wgt_6_477;
		WeightsStore6[478] <= Wgt_6_478;
		WeightsStore6[479] <= Wgt_6_479;
		WeightsStore6[480] <= Wgt_6_480;
		WeightsStore6[481] <= Wgt_6_481;
		WeightsStore6[482] <= Wgt_6_482;
		WeightsStore6[483] <= Wgt_6_483;
		WeightsStore6[484] <= Wgt_6_484;
		WeightsStore6[485] <= Wgt_6_485;
		WeightsStore6[486] <= Wgt_6_486;
		WeightsStore6[487] <= Wgt_6_487;
		WeightsStore6[488] <= Wgt_6_488;
		WeightsStore6[489] <= Wgt_6_489;
		WeightsStore6[490] <= Wgt_6_490;
		WeightsStore6[491] <= Wgt_6_491;
		WeightsStore6[492] <= Wgt_6_492;
		WeightsStore6[493] <= Wgt_6_493;
		WeightsStore6[494] <= Wgt_6_494;
		WeightsStore6[495] <= Wgt_6_495;
		WeightsStore6[496] <= Wgt_6_496;
		WeightsStore6[497] <= Wgt_6_497;
		WeightsStore6[498] <= Wgt_6_498;
		WeightsStore6[499] <= Wgt_6_499;
		WeightsStore6[500] <= Wgt_6_500;
		WeightsStore6[501] <= Wgt_6_501;
		WeightsStore6[502] <= Wgt_6_502;
		WeightsStore6[503] <= Wgt_6_503;
		WeightsStore6[504] <= Wgt_6_504;
		WeightsStore6[505] <= Wgt_6_505;
		WeightsStore6[506] <= Wgt_6_506;
		WeightsStore6[507] <= Wgt_6_507;
		WeightsStore6[508] <= Wgt_6_508;
		WeightsStore6[509] <= Wgt_6_509;
		WeightsStore6[510] <= Wgt_6_510;
		WeightsStore6[511] <= Wgt_6_511;
		WeightsStore6[512] <= Wgt_6_512;
		WeightsStore6[513] <= Wgt_6_513;
		WeightsStore6[514] <= Wgt_6_514;
		WeightsStore6[515] <= Wgt_6_515;
		WeightsStore6[516] <= Wgt_6_516;
		WeightsStore6[517] <= Wgt_6_517;
		WeightsStore6[518] <= Wgt_6_518;
		WeightsStore6[519] <= Wgt_6_519;
		WeightsStore6[520] <= Wgt_6_520;
		WeightsStore6[521] <= Wgt_6_521;
		WeightsStore6[522] <= Wgt_6_522;
		WeightsStore6[523] <= Wgt_6_523;
		WeightsStore6[524] <= Wgt_6_524;
		WeightsStore6[525] <= Wgt_6_525;
		WeightsStore6[526] <= Wgt_6_526;
		WeightsStore6[527] <= Wgt_6_527;
		WeightsStore6[528] <= Wgt_6_528;
		WeightsStore6[529] <= Wgt_6_529;
		WeightsStore6[530] <= Wgt_6_530;
		WeightsStore6[531] <= Wgt_6_531;
		WeightsStore6[532] <= Wgt_6_532;
		WeightsStore6[533] <= Wgt_6_533;
		WeightsStore6[534] <= Wgt_6_534;
		WeightsStore6[535] <= Wgt_6_535;
		WeightsStore6[536] <= Wgt_6_536;
		WeightsStore6[537] <= Wgt_6_537;
		WeightsStore6[538] <= Wgt_6_538;
		WeightsStore6[539] <= Wgt_6_539;
		WeightsStore6[540] <= Wgt_6_540;
		WeightsStore6[541] <= Wgt_6_541;
		WeightsStore6[542] <= Wgt_6_542;
		WeightsStore6[543] <= Wgt_6_543;
		WeightsStore6[544] <= Wgt_6_544;
		WeightsStore6[545] <= Wgt_6_545;
		WeightsStore6[546] <= Wgt_6_546;
		WeightsStore6[547] <= Wgt_6_547;
		WeightsStore6[548] <= Wgt_6_548;
		WeightsStore6[549] <= Wgt_6_549;
		WeightsStore6[550] <= Wgt_6_550;
		WeightsStore6[551] <= Wgt_6_551;
		WeightsStore6[552] <= Wgt_6_552;
		WeightsStore6[553] <= Wgt_6_553;
		WeightsStore6[554] <= Wgt_6_554;
		WeightsStore6[555] <= Wgt_6_555;
		WeightsStore6[556] <= Wgt_6_556;
		WeightsStore6[557] <= Wgt_6_557;
		WeightsStore6[558] <= Wgt_6_558;
		WeightsStore6[559] <= Wgt_6_559;
		WeightsStore6[560] <= Wgt_6_560;
		WeightsStore6[561] <= Wgt_6_561;
		WeightsStore6[562] <= Wgt_6_562;
		WeightsStore6[563] <= Wgt_6_563;
		WeightsStore6[564] <= Wgt_6_564;
		WeightsStore6[565] <= Wgt_6_565;
		WeightsStore6[566] <= Wgt_6_566;
		WeightsStore6[567] <= Wgt_6_567;
		WeightsStore6[568] <= Wgt_6_568;
		WeightsStore6[569] <= Wgt_6_569;
		WeightsStore6[570] <= Wgt_6_570;
		WeightsStore6[571] <= Wgt_6_571;
		WeightsStore6[572] <= Wgt_6_572;
		WeightsStore6[573] <= Wgt_6_573;
		WeightsStore6[574] <= Wgt_6_574;
		WeightsStore6[575] <= Wgt_6_575;
		WeightsStore6[576] <= Wgt_6_576;
		WeightsStore6[577] <= Wgt_6_577;
		WeightsStore6[578] <= Wgt_6_578;
		WeightsStore6[579] <= Wgt_6_579;
		WeightsStore6[580] <= Wgt_6_580;
		WeightsStore6[581] <= Wgt_6_581;
		WeightsStore6[582] <= Wgt_6_582;
		WeightsStore6[583] <= Wgt_6_583;
		WeightsStore6[584] <= Wgt_6_584;
		WeightsStore6[585] <= Wgt_6_585;
		WeightsStore6[586] <= Wgt_6_586;
		WeightsStore6[587] <= Wgt_6_587;
		WeightsStore6[588] <= Wgt_6_588;
		WeightsStore6[589] <= Wgt_6_589;
		WeightsStore6[590] <= Wgt_6_590;
		WeightsStore6[591] <= Wgt_6_591;
		WeightsStore6[592] <= Wgt_6_592;
		WeightsStore6[593] <= Wgt_6_593;
		WeightsStore6[594] <= Wgt_6_594;
		WeightsStore6[595] <= Wgt_6_595;
		WeightsStore6[596] <= Wgt_6_596;
		WeightsStore6[597] <= Wgt_6_597;
		WeightsStore6[598] <= Wgt_6_598;
		WeightsStore6[599] <= Wgt_6_599;
		WeightsStore6[600] <= Wgt_6_600;
		WeightsStore6[601] <= Wgt_6_601;
		WeightsStore6[602] <= Wgt_6_602;
		WeightsStore6[603] <= Wgt_6_603;
		WeightsStore6[604] <= Wgt_6_604;
		WeightsStore6[605] <= Wgt_6_605;
		WeightsStore6[606] <= Wgt_6_606;
		WeightsStore6[607] <= Wgt_6_607;
		WeightsStore6[608] <= Wgt_6_608;
		WeightsStore6[609] <= Wgt_6_609;
		WeightsStore6[610] <= Wgt_6_610;
		WeightsStore6[611] <= Wgt_6_611;
		WeightsStore6[612] <= Wgt_6_612;
		WeightsStore6[613] <= Wgt_6_613;
		WeightsStore6[614] <= Wgt_6_614;
		WeightsStore6[615] <= Wgt_6_615;
		WeightsStore6[616] <= Wgt_6_616;
		WeightsStore6[617] <= Wgt_6_617;
		WeightsStore6[618] <= Wgt_6_618;
		WeightsStore6[619] <= Wgt_6_619;
		WeightsStore6[620] <= Wgt_6_620;
		WeightsStore6[621] <= Wgt_6_621;
		WeightsStore6[622] <= Wgt_6_622;
		WeightsStore6[623] <= Wgt_6_623;
		WeightsStore6[624] <= Wgt_6_624;
		WeightsStore6[625] <= Wgt_6_625;
		WeightsStore6[626] <= Wgt_6_626;
		WeightsStore6[627] <= Wgt_6_627;
		WeightsStore6[628] <= Wgt_6_628;
		WeightsStore6[629] <= Wgt_6_629;
		WeightsStore6[630] <= Wgt_6_630;
		WeightsStore6[631] <= Wgt_6_631;
		WeightsStore6[632] <= Wgt_6_632;
		WeightsStore6[633] <= Wgt_6_633;
		WeightsStore6[634] <= Wgt_6_634;
		WeightsStore6[635] <= Wgt_6_635;
		WeightsStore6[636] <= Wgt_6_636;
		WeightsStore6[637] <= Wgt_6_637;
		WeightsStore6[638] <= Wgt_6_638;
		WeightsStore6[639] <= Wgt_6_639;
		WeightsStore6[640] <= Wgt_6_640;
		WeightsStore6[641] <= Wgt_6_641;
		WeightsStore6[642] <= Wgt_6_642;
		WeightsStore6[643] <= Wgt_6_643;
		WeightsStore6[644] <= Wgt_6_644;
		WeightsStore6[645] <= Wgt_6_645;
		WeightsStore6[646] <= Wgt_6_646;
		WeightsStore6[647] <= Wgt_6_647;
		WeightsStore6[648] <= Wgt_6_648;
		WeightsStore6[649] <= Wgt_6_649;
		WeightsStore6[650] <= Wgt_6_650;
		WeightsStore6[651] <= Wgt_6_651;
		WeightsStore6[652] <= Wgt_6_652;
		WeightsStore6[653] <= Wgt_6_653;
		WeightsStore6[654] <= Wgt_6_654;
		WeightsStore6[655] <= Wgt_6_655;
		WeightsStore6[656] <= Wgt_6_656;
		WeightsStore6[657] <= Wgt_6_657;
		WeightsStore6[658] <= Wgt_6_658;
		WeightsStore6[659] <= Wgt_6_659;
		WeightsStore6[660] <= Wgt_6_660;
		WeightsStore6[661] <= Wgt_6_661;
		WeightsStore6[662] <= Wgt_6_662;
		WeightsStore6[663] <= Wgt_6_663;
		WeightsStore6[664] <= Wgt_6_664;
		WeightsStore6[665] <= Wgt_6_665;
		WeightsStore6[666] <= Wgt_6_666;
		WeightsStore6[667] <= Wgt_6_667;
		WeightsStore6[668] <= Wgt_6_668;
		WeightsStore6[669] <= Wgt_6_669;
		WeightsStore6[670] <= Wgt_6_670;
		WeightsStore6[671] <= Wgt_6_671;
		WeightsStore6[672] <= Wgt_6_672;
		WeightsStore6[673] <= Wgt_6_673;
		WeightsStore6[674] <= Wgt_6_674;
		WeightsStore6[675] <= Wgt_6_675;
		WeightsStore6[676] <= Wgt_6_676;
		WeightsStore6[677] <= Wgt_6_677;
		WeightsStore6[678] <= Wgt_6_678;
		WeightsStore6[679] <= Wgt_6_679;
		WeightsStore6[680] <= Wgt_6_680;
		WeightsStore6[681] <= Wgt_6_681;
		WeightsStore6[682] <= Wgt_6_682;
		WeightsStore6[683] <= Wgt_6_683;
		WeightsStore6[684] <= Wgt_6_684;
		WeightsStore6[685] <= Wgt_6_685;
		WeightsStore6[686] <= Wgt_6_686;
		WeightsStore6[687] <= Wgt_6_687;
		WeightsStore6[688] <= Wgt_6_688;
		WeightsStore6[689] <= Wgt_6_689;
		WeightsStore6[690] <= Wgt_6_690;
		WeightsStore6[691] <= Wgt_6_691;
		WeightsStore6[692] <= Wgt_6_692;
		WeightsStore6[693] <= Wgt_6_693;
		WeightsStore6[694] <= Wgt_6_694;
		WeightsStore6[695] <= Wgt_6_695;
		WeightsStore6[696] <= Wgt_6_696;
		WeightsStore6[697] <= Wgt_6_697;
		WeightsStore6[698] <= Wgt_6_698;
		WeightsStore6[699] <= Wgt_6_699;
		WeightsStore6[700] <= Wgt_6_700;
		WeightsStore6[701] <= Wgt_6_701;
		WeightsStore6[702] <= Wgt_6_702;
		WeightsStore6[703] <= Wgt_6_703;
		WeightsStore6[704] <= Wgt_6_704;
		WeightsStore6[705] <= Wgt_6_705;
		WeightsStore6[706] <= Wgt_6_706;
		WeightsStore6[707] <= Wgt_6_707;
		WeightsStore6[708] <= Wgt_6_708;
		WeightsStore6[709] <= Wgt_6_709;
		WeightsStore6[710] <= Wgt_6_710;
		WeightsStore6[711] <= Wgt_6_711;
		WeightsStore6[712] <= Wgt_6_712;
		WeightsStore6[713] <= Wgt_6_713;
		WeightsStore6[714] <= Wgt_6_714;
		WeightsStore6[715] <= Wgt_6_715;
		WeightsStore6[716] <= Wgt_6_716;
		WeightsStore6[717] <= Wgt_6_717;
		WeightsStore6[718] <= Wgt_6_718;
		WeightsStore6[719] <= Wgt_6_719;
		WeightsStore6[720] <= Wgt_6_720;
		WeightsStore6[721] <= Wgt_6_721;
		WeightsStore6[722] <= Wgt_6_722;
		WeightsStore6[723] <= Wgt_6_723;
		WeightsStore6[724] <= Wgt_6_724;
		WeightsStore6[725] <= Wgt_6_725;
		WeightsStore6[726] <= Wgt_6_726;
		WeightsStore6[727] <= Wgt_6_727;
		WeightsStore6[728] <= Wgt_6_728;
		WeightsStore6[729] <= Wgt_6_729;
		WeightsStore6[730] <= Wgt_6_730;
		WeightsStore6[731] <= Wgt_6_731;
		WeightsStore6[732] <= Wgt_6_732;
		WeightsStore6[733] <= Wgt_6_733;
		WeightsStore6[734] <= Wgt_6_734;
		WeightsStore6[735] <= Wgt_6_735;
		WeightsStore6[736] <= Wgt_6_736;
		WeightsStore6[737] <= Wgt_6_737;
		WeightsStore6[738] <= Wgt_6_738;
		WeightsStore6[739] <= Wgt_6_739;
		WeightsStore6[740] <= Wgt_6_740;
		WeightsStore6[741] <= Wgt_6_741;
		WeightsStore6[742] <= Wgt_6_742;
		WeightsStore6[743] <= Wgt_6_743;
		WeightsStore6[744] <= Wgt_6_744;
		WeightsStore6[745] <= Wgt_6_745;
		WeightsStore6[746] <= Wgt_6_746;
		WeightsStore6[747] <= Wgt_6_747;
		WeightsStore6[748] <= Wgt_6_748;
		WeightsStore6[749] <= Wgt_6_749;
		WeightsStore6[750] <= Wgt_6_750;
		WeightsStore6[751] <= Wgt_6_751;
		WeightsStore6[752] <= Wgt_6_752;
		WeightsStore6[753] <= Wgt_6_753;
		WeightsStore6[754] <= Wgt_6_754;
		WeightsStore6[755] <= Wgt_6_755;
		WeightsStore6[756] <= Wgt_6_756;
		WeightsStore6[757] <= Wgt_6_757;
		WeightsStore6[758] <= Wgt_6_758;
		WeightsStore6[759] <= Wgt_6_759;
		WeightsStore6[760] <= Wgt_6_760;
		WeightsStore6[761] <= Wgt_6_761;
		WeightsStore6[762] <= Wgt_6_762;
		WeightsStore6[763] <= Wgt_6_763;
		WeightsStore6[764] <= Wgt_6_764;
		WeightsStore6[765] <= Wgt_6_765;
		WeightsStore6[766] <= Wgt_6_766;
		WeightsStore6[767] <= Wgt_6_767;
		WeightsStore6[768] <= Wgt_6_768;
		WeightsStore6[769] <= Wgt_6_769;
		WeightsStore6[770] <= Wgt_6_770;
		WeightsStore6[771] <= Wgt_6_771;
		WeightsStore6[772] <= Wgt_6_772;
		WeightsStore6[773] <= Wgt_6_773;
		WeightsStore6[774] <= Wgt_6_774;
		WeightsStore6[775] <= Wgt_6_775;
		WeightsStore6[776] <= Wgt_6_776;
		WeightsStore6[777] <= Wgt_6_777;
		WeightsStore6[778] <= Wgt_6_778;
		WeightsStore6[779] <= Wgt_6_779;
		WeightsStore6[780] <= Wgt_6_780;
		WeightsStore6[781] <= Wgt_6_781;
		WeightsStore6[782] <= Wgt_6_782;
		WeightsStore6[783] <= Wgt_6_783;
		WeightsStore6[784] <= Wgt_6_784;
		WeightsStore7[0] <= Wgt_7_0;
		WeightsStore7[1] <= Wgt_7_1;
		WeightsStore7[2] <= Wgt_7_2;
		WeightsStore7[3] <= Wgt_7_3;
		WeightsStore7[4] <= Wgt_7_4;
		WeightsStore7[5] <= Wgt_7_5;
		WeightsStore7[6] <= Wgt_7_6;
		WeightsStore7[7] <= Wgt_7_7;
		WeightsStore7[8] <= Wgt_7_8;
		WeightsStore7[9] <= Wgt_7_9;
		WeightsStore7[10] <= Wgt_7_10;
		WeightsStore7[11] <= Wgt_7_11;
		WeightsStore7[12] <= Wgt_7_12;
		WeightsStore7[13] <= Wgt_7_13;
		WeightsStore7[14] <= Wgt_7_14;
		WeightsStore7[15] <= Wgt_7_15;
		WeightsStore7[16] <= Wgt_7_16;
		WeightsStore7[17] <= Wgt_7_17;
		WeightsStore7[18] <= Wgt_7_18;
		WeightsStore7[19] <= Wgt_7_19;
		WeightsStore7[20] <= Wgt_7_20;
		WeightsStore7[21] <= Wgt_7_21;
		WeightsStore7[22] <= Wgt_7_22;
		WeightsStore7[23] <= Wgt_7_23;
		WeightsStore7[24] <= Wgt_7_24;
		WeightsStore7[25] <= Wgt_7_25;
		WeightsStore7[26] <= Wgt_7_26;
		WeightsStore7[27] <= Wgt_7_27;
		WeightsStore7[28] <= Wgt_7_28;
		WeightsStore7[29] <= Wgt_7_29;
		WeightsStore7[30] <= Wgt_7_30;
		WeightsStore7[31] <= Wgt_7_31;
		WeightsStore7[32] <= Wgt_7_32;
		WeightsStore7[33] <= Wgt_7_33;
		WeightsStore7[34] <= Wgt_7_34;
		WeightsStore7[35] <= Wgt_7_35;
		WeightsStore7[36] <= Wgt_7_36;
		WeightsStore7[37] <= Wgt_7_37;
		WeightsStore7[38] <= Wgt_7_38;
		WeightsStore7[39] <= Wgt_7_39;
		WeightsStore7[40] <= Wgt_7_40;
		WeightsStore7[41] <= Wgt_7_41;
		WeightsStore7[42] <= Wgt_7_42;
		WeightsStore7[43] <= Wgt_7_43;
		WeightsStore7[44] <= Wgt_7_44;
		WeightsStore7[45] <= Wgt_7_45;
		WeightsStore7[46] <= Wgt_7_46;
		WeightsStore7[47] <= Wgt_7_47;
		WeightsStore7[48] <= Wgt_7_48;
		WeightsStore7[49] <= Wgt_7_49;
		WeightsStore7[50] <= Wgt_7_50;
		WeightsStore7[51] <= Wgt_7_51;
		WeightsStore7[52] <= Wgt_7_52;
		WeightsStore7[53] <= Wgt_7_53;
		WeightsStore7[54] <= Wgt_7_54;
		WeightsStore7[55] <= Wgt_7_55;
		WeightsStore7[56] <= Wgt_7_56;
		WeightsStore7[57] <= Wgt_7_57;
		WeightsStore7[58] <= Wgt_7_58;
		WeightsStore7[59] <= Wgt_7_59;
		WeightsStore7[60] <= Wgt_7_60;
		WeightsStore7[61] <= Wgt_7_61;
		WeightsStore7[62] <= Wgt_7_62;
		WeightsStore7[63] <= Wgt_7_63;
		WeightsStore7[64] <= Wgt_7_64;
		WeightsStore7[65] <= Wgt_7_65;
		WeightsStore7[66] <= Wgt_7_66;
		WeightsStore7[67] <= Wgt_7_67;
		WeightsStore7[68] <= Wgt_7_68;
		WeightsStore7[69] <= Wgt_7_69;
		WeightsStore7[70] <= Wgt_7_70;
		WeightsStore7[71] <= Wgt_7_71;
		WeightsStore7[72] <= Wgt_7_72;
		WeightsStore7[73] <= Wgt_7_73;
		WeightsStore7[74] <= Wgt_7_74;
		WeightsStore7[75] <= Wgt_7_75;
		WeightsStore7[76] <= Wgt_7_76;
		WeightsStore7[77] <= Wgt_7_77;
		WeightsStore7[78] <= Wgt_7_78;
		WeightsStore7[79] <= Wgt_7_79;
		WeightsStore7[80] <= Wgt_7_80;
		WeightsStore7[81] <= Wgt_7_81;
		WeightsStore7[82] <= Wgt_7_82;
		WeightsStore7[83] <= Wgt_7_83;
		WeightsStore7[84] <= Wgt_7_84;
		WeightsStore7[85] <= Wgt_7_85;
		WeightsStore7[86] <= Wgt_7_86;
		WeightsStore7[87] <= Wgt_7_87;
		WeightsStore7[88] <= Wgt_7_88;
		WeightsStore7[89] <= Wgt_7_89;
		WeightsStore7[90] <= Wgt_7_90;
		WeightsStore7[91] <= Wgt_7_91;
		WeightsStore7[92] <= Wgt_7_92;
		WeightsStore7[93] <= Wgt_7_93;
		WeightsStore7[94] <= Wgt_7_94;
		WeightsStore7[95] <= Wgt_7_95;
		WeightsStore7[96] <= Wgt_7_96;
		WeightsStore7[97] <= Wgt_7_97;
		WeightsStore7[98] <= Wgt_7_98;
		WeightsStore7[99] <= Wgt_7_99;
		WeightsStore7[100] <= Wgt_7_100;
		WeightsStore7[101] <= Wgt_7_101;
		WeightsStore7[102] <= Wgt_7_102;
		WeightsStore7[103] <= Wgt_7_103;
		WeightsStore7[104] <= Wgt_7_104;
		WeightsStore7[105] <= Wgt_7_105;
		WeightsStore7[106] <= Wgt_7_106;
		WeightsStore7[107] <= Wgt_7_107;
		WeightsStore7[108] <= Wgt_7_108;
		WeightsStore7[109] <= Wgt_7_109;
		WeightsStore7[110] <= Wgt_7_110;
		WeightsStore7[111] <= Wgt_7_111;
		WeightsStore7[112] <= Wgt_7_112;
		WeightsStore7[113] <= Wgt_7_113;
		WeightsStore7[114] <= Wgt_7_114;
		WeightsStore7[115] <= Wgt_7_115;
		WeightsStore7[116] <= Wgt_7_116;
		WeightsStore7[117] <= Wgt_7_117;
		WeightsStore7[118] <= Wgt_7_118;
		WeightsStore7[119] <= Wgt_7_119;
		WeightsStore7[120] <= Wgt_7_120;
		WeightsStore7[121] <= Wgt_7_121;
		WeightsStore7[122] <= Wgt_7_122;
		WeightsStore7[123] <= Wgt_7_123;
		WeightsStore7[124] <= Wgt_7_124;
		WeightsStore7[125] <= Wgt_7_125;
		WeightsStore7[126] <= Wgt_7_126;
		WeightsStore7[127] <= Wgt_7_127;
		WeightsStore7[128] <= Wgt_7_128;
		WeightsStore7[129] <= Wgt_7_129;
		WeightsStore7[130] <= Wgt_7_130;
		WeightsStore7[131] <= Wgt_7_131;
		WeightsStore7[132] <= Wgt_7_132;
		WeightsStore7[133] <= Wgt_7_133;
		WeightsStore7[134] <= Wgt_7_134;
		WeightsStore7[135] <= Wgt_7_135;
		WeightsStore7[136] <= Wgt_7_136;
		WeightsStore7[137] <= Wgt_7_137;
		WeightsStore7[138] <= Wgt_7_138;
		WeightsStore7[139] <= Wgt_7_139;
		WeightsStore7[140] <= Wgt_7_140;
		WeightsStore7[141] <= Wgt_7_141;
		WeightsStore7[142] <= Wgt_7_142;
		WeightsStore7[143] <= Wgt_7_143;
		WeightsStore7[144] <= Wgt_7_144;
		WeightsStore7[145] <= Wgt_7_145;
		WeightsStore7[146] <= Wgt_7_146;
		WeightsStore7[147] <= Wgt_7_147;
		WeightsStore7[148] <= Wgt_7_148;
		WeightsStore7[149] <= Wgt_7_149;
		WeightsStore7[150] <= Wgt_7_150;
		WeightsStore7[151] <= Wgt_7_151;
		WeightsStore7[152] <= Wgt_7_152;
		WeightsStore7[153] <= Wgt_7_153;
		WeightsStore7[154] <= Wgt_7_154;
		WeightsStore7[155] <= Wgt_7_155;
		WeightsStore7[156] <= Wgt_7_156;
		WeightsStore7[157] <= Wgt_7_157;
		WeightsStore7[158] <= Wgt_7_158;
		WeightsStore7[159] <= Wgt_7_159;
		WeightsStore7[160] <= Wgt_7_160;
		WeightsStore7[161] <= Wgt_7_161;
		WeightsStore7[162] <= Wgt_7_162;
		WeightsStore7[163] <= Wgt_7_163;
		WeightsStore7[164] <= Wgt_7_164;
		WeightsStore7[165] <= Wgt_7_165;
		WeightsStore7[166] <= Wgt_7_166;
		WeightsStore7[167] <= Wgt_7_167;
		WeightsStore7[168] <= Wgt_7_168;
		WeightsStore7[169] <= Wgt_7_169;
		WeightsStore7[170] <= Wgt_7_170;
		WeightsStore7[171] <= Wgt_7_171;
		WeightsStore7[172] <= Wgt_7_172;
		WeightsStore7[173] <= Wgt_7_173;
		WeightsStore7[174] <= Wgt_7_174;
		WeightsStore7[175] <= Wgt_7_175;
		WeightsStore7[176] <= Wgt_7_176;
		WeightsStore7[177] <= Wgt_7_177;
		WeightsStore7[178] <= Wgt_7_178;
		WeightsStore7[179] <= Wgt_7_179;
		WeightsStore7[180] <= Wgt_7_180;
		WeightsStore7[181] <= Wgt_7_181;
		WeightsStore7[182] <= Wgt_7_182;
		WeightsStore7[183] <= Wgt_7_183;
		WeightsStore7[184] <= Wgt_7_184;
		WeightsStore7[185] <= Wgt_7_185;
		WeightsStore7[186] <= Wgt_7_186;
		WeightsStore7[187] <= Wgt_7_187;
		WeightsStore7[188] <= Wgt_7_188;
		WeightsStore7[189] <= Wgt_7_189;
		WeightsStore7[190] <= Wgt_7_190;
		WeightsStore7[191] <= Wgt_7_191;
		WeightsStore7[192] <= Wgt_7_192;
		WeightsStore7[193] <= Wgt_7_193;
		WeightsStore7[194] <= Wgt_7_194;
		WeightsStore7[195] <= Wgt_7_195;
		WeightsStore7[196] <= Wgt_7_196;
		WeightsStore7[197] <= Wgt_7_197;
		WeightsStore7[198] <= Wgt_7_198;
		WeightsStore7[199] <= Wgt_7_199;
		WeightsStore7[200] <= Wgt_7_200;
		WeightsStore7[201] <= Wgt_7_201;
		WeightsStore7[202] <= Wgt_7_202;
		WeightsStore7[203] <= Wgt_7_203;
		WeightsStore7[204] <= Wgt_7_204;
		WeightsStore7[205] <= Wgt_7_205;
		WeightsStore7[206] <= Wgt_7_206;
		WeightsStore7[207] <= Wgt_7_207;
		WeightsStore7[208] <= Wgt_7_208;
		WeightsStore7[209] <= Wgt_7_209;
		WeightsStore7[210] <= Wgt_7_210;
		WeightsStore7[211] <= Wgt_7_211;
		WeightsStore7[212] <= Wgt_7_212;
		WeightsStore7[213] <= Wgt_7_213;
		WeightsStore7[214] <= Wgt_7_214;
		WeightsStore7[215] <= Wgt_7_215;
		WeightsStore7[216] <= Wgt_7_216;
		WeightsStore7[217] <= Wgt_7_217;
		WeightsStore7[218] <= Wgt_7_218;
		WeightsStore7[219] <= Wgt_7_219;
		WeightsStore7[220] <= Wgt_7_220;
		WeightsStore7[221] <= Wgt_7_221;
		WeightsStore7[222] <= Wgt_7_222;
		WeightsStore7[223] <= Wgt_7_223;
		WeightsStore7[224] <= Wgt_7_224;
		WeightsStore7[225] <= Wgt_7_225;
		WeightsStore7[226] <= Wgt_7_226;
		WeightsStore7[227] <= Wgt_7_227;
		WeightsStore7[228] <= Wgt_7_228;
		WeightsStore7[229] <= Wgt_7_229;
		WeightsStore7[230] <= Wgt_7_230;
		WeightsStore7[231] <= Wgt_7_231;
		WeightsStore7[232] <= Wgt_7_232;
		WeightsStore7[233] <= Wgt_7_233;
		WeightsStore7[234] <= Wgt_7_234;
		WeightsStore7[235] <= Wgt_7_235;
		WeightsStore7[236] <= Wgt_7_236;
		WeightsStore7[237] <= Wgt_7_237;
		WeightsStore7[238] <= Wgt_7_238;
		WeightsStore7[239] <= Wgt_7_239;
		WeightsStore7[240] <= Wgt_7_240;
		WeightsStore7[241] <= Wgt_7_241;
		WeightsStore7[242] <= Wgt_7_242;
		WeightsStore7[243] <= Wgt_7_243;
		WeightsStore7[244] <= Wgt_7_244;
		WeightsStore7[245] <= Wgt_7_245;
		WeightsStore7[246] <= Wgt_7_246;
		WeightsStore7[247] <= Wgt_7_247;
		WeightsStore7[248] <= Wgt_7_248;
		WeightsStore7[249] <= Wgt_7_249;
		WeightsStore7[250] <= Wgt_7_250;
		WeightsStore7[251] <= Wgt_7_251;
		WeightsStore7[252] <= Wgt_7_252;
		WeightsStore7[253] <= Wgt_7_253;
		WeightsStore7[254] <= Wgt_7_254;
		WeightsStore7[255] <= Wgt_7_255;
		WeightsStore7[256] <= Wgt_7_256;
		WeightsStore7[257] <= Wgt_7_257;
		WeightsStore7[258] <= Wgt_7_258;
		WeightsStore7[259] <= Wgt_7_259;
		WeightsStore7[260] <= Wgt_7_260;
		WeightsStore7[261] <= Wgt_7_261;
		WeightsStore7[262] <= Wgt_7_262;
		WeightsStore7[263] <= Wgt_7_263;
		WeightsStore7[264] <= Wgt_7_264;
		WeightsStore7[265] <= Wgt_7_265;
		WeightsStore7[266] <= Wgt_7_266;
		WeightsStore7[267] <= Wgt_7_267;
		WeightsStore7[268] <= Wgt_7_268;
		WeightsStore7[269] <= Wgt_7_269;
		WeightsStore7[270] <= Wgt_7_270;
		WeightsStore7[271] <= Wgt_7_271;
		WeightsStore7[272] <= Wgt_7_272;
		WeightsStore7[273] <= Wgt_7_273;
		WeightsStore7[274] <= Wgt_7_274;
		WeightsStore7[275] <= Wgt_7_275;
		WeightsStore7[276] <= Wgt_7_276;
		WeightsStore7[277] <= Wgt_7_277;
		WeightsStore7[278] <= Wgt_7_278;
		WeightsStore7[279] <= Wgt_7_279;
		WeightsStore7[280] <= Wgt_7_280;
		WeightsStore7[281] <= Wgt_7_281;
		WeightsStore7[282] <= Wgt_7_282;
		WeightsStore7[283] <= Wgt_7_283;
		WeightsStore7[284] <= Wgt_7_284;
		WeightsStore7[285] <= Wgt_7_285;
		WeightsStore7[286] <= Wgt_7_286;
		WeightsStore7[287] <= Wgt_7_287;
		WeightsStore7[288] <= Wgt_7_288;
		WeightsStore7[289] <= Wgt_7_289;
		WeightsStore7[290] <= Wgt_7_290;
		WeightsStore7[291] <= Wgt_7_291;
		WeightsStore7[292] <= Wgt_7_292;
		WeightsStore7[293] <= Wgt_7_293;
		WeightsStore7[294] <= Wgt_7_294;
		WeightsStore7[295] <= Wgt_7_295;
		WeightsStore7[296] <= Wgt_7_296;
		WeightsStore7[297] <= Wgt_7_297;
		WeightsStore7[298] <= Wgt_7_298;
		WeightsStore7[299] <= Wgt_7_299;
		WeightsStore7[300] <= Wgt_7_300;
		WeightsStore7[301] <= Wgt_7_301;
		WeightsStore7[302] <= Wgt_7_302;
		WeightsStore7[303] <= Wgt_7_303;
		WeightsStore7[304] <= Wgt_7_304;
		WeightsStore7[305] <= Wgt_7_305;
		WeightsStore7[306] <= Wgt_7_306;
		WeightsStore7[307] <= Wgt_7_307;
		WeightsStore7[308] <= Wgt_7_308;
		WeightsStore7[309] <= Wgt_7_309;
		WeightsStore7[310] <= Wgt_7_310;
		WeightsStore7[311] <= Wgt_7_311;
		WeightsStore7[312] <= Wgt_7_312;
		WeightsStore7[313] <= Wgt_7_313;
		WeightsStore7[314] <= Wgt_7_314;
		WeightsStore7[315] <= Wgt_7_315;
		WeightsStore7[316] <= Wgt_7_316;
		WeightsStore7[317] <= Wgt_7_317;
		WeightsStore7[318] <= Wgt_7_318;
		WeightsStore7[319] <= Wgt_7_319;
		WeightsStore7[320] <= Wgt_7_320;
		WeightsStore7[321] <= Wgt_7_321;
		WeightsStore7[322] <= Wgt_7_322;
		WeightsStore7[323] <= Wgt_7_323;
		WeightsStore7[324] <= Wgt_7_324;
		WeightsStore7[325] <= Wgt_7_325;
		WeightsStore7[326] <= Wgt_7_326;
		WeightsStore7[327] <= Wgt_7_327;
		WeightsStore7[328] <= Wgt_7_328;
		WeightsStore7[329] <= Wgt_7_329;
		WeightsStore7[330] <= Wgt_7_330;
		WeightsStore7[331] <= Wgt_7_331;
		WeightsStore7[332] <= Wgt_7_332;
		WeightsStore7[333] <= Wgt_7_333;
		WeightsStore7[334] <= Wgt_7_334;
		WeightsStore7[335] <= Wgt_7_335;
		WeightsStore7[336] <= Wgt_7_336;
		WeightsStore7[337] <= Wgt_7_337;
		WeightsStore7[338] <= Wgt_7_338;
		WeightsStore7[339] <= Wgt_7_339;
		WeightsStore7[340] <= Wgt_7_340;
		WeightsStore7[341] <= Wgt_7_341;
		WeightsStore7[342] <= Wgt_7_342;
		WeightsStore7[343] <= Wgt_7_343;
		WeightsStore7[344] <= Wgt_7_344;
		WeightsStore7[345] <= Wgt_7_345;
		WeightsStore7[346] <= Wgt_7_346;
		WeightsStore7[347] <= Wgt_7_347;
		WeightsStore7[348] <= Wgt_7_348;
		WeightsStore7[349] <= Wgt_7_349;
		WeightsStore7[350] <= Wgt_7_350;
		WeightsStore7[351] <= Wgt_7_351;
		WeightsStore7[352] <= Wgt_7_352;
		WeightsStore7[353] <= Wgt_7_353;
		WeightsStore7[354] <= Wgt_7_354;
		WeightsStore7[355] <= Wgt_7_355;
		WeightsStore7[356] <= Wgt_7_356;
		WeightsStore7[357] <= Wgt_7_357;
		WeightsStore7[358] <= Wgt_7_358;
		WeightsStore7[359] <= Wgt_7_359;
		WeightsStore7[360] <= Wgt_7_360;
		WeightsStore7[361] <= Wgt_7_361;
		WeightsStore7[362] <= Wgt_7_362;
		WeightsStore7[363] <= Wgt_7_363;
		WeightsStore7[364] <= Wgt_7_364;
		WeightsStore7[365] <= Wgt_7_365;
		WeightsStore7[366] <= Wgt_7_366;
		WeightsStore7[367] <= Wgt_7_367;
		WeightsStore7[368] <= Wgt_7_368;
		WeightsStore7[369] <= Wgt_7_369;
		WeightsStore7[370] <= Wgt_7_370;
		WeightsStore7[371] <= Wgt_7_371;
		WeightsStore7[372] <= Wgt_7_372;
		WeightsStore7[373] <= Wgt_7_373;
		WeightsStore7[374] <= Wgt_7_374;
		WeightsStore7[375] <= Wgt_7_375;
		WeightsStore7[376] <= Wgt_7_376;
		WeightsStore7[377] <= Wgt_7_377;
		WeightsStore7[378] <= Wgt_7_378;
		WeightsStore7[379] <= Wgt_7_379;
		WeightsStore7[380] <= Wgt_7_380;
		WeightsStore7[381] <= Wgt_7_381;
		WeightsStore7[382] <= Wgt_7_382;
		WeightsStore7[383] <= Wgt_7_383;
		WeightsStore7[384] <= Wgt_7_384;
		WeightsStore7[385] <= Wgt_7_385;
		WeightsStore7[386] <= Wgt_7_386;
		WeightsStore7[387] <= Wgt_7_387;
		WeightsStore7[388] <= Wgt_7_388;
		WeightsStore7[389] <= Wgt_7_389;
		WeightsStore7[390] <= Wgt_7_390;
		WeightsStore7[391] <= Wgt_7_391;
		WeightsStore7[392] <= Wgt_7_392;
		WeightsStore7[393] <= Wgt_7_393;
		WeightsStore7[394] <= Wgt_7_394;
		WeightsStore7[395] <= Wgt_7_395;
		WeightsStore7[396] <= Wgt_7_396;
		WeightsStore7[397] <= Wgt_7_397;
		WeightsStore7[398] <= Wgt_7_398;
		WeightsStore7[399] <= Wgt_7_399;
		WeightsStore7[400] <= Wgt_7_400;
		WeightsStore7[401] <= Wgt_7_401;
		WeightsStore7[402] <= Wgt_7_402;
		WeightsStore7[403] <= Wgt_7_403;
		WeightsStore7[404] <= Wgt_7_404;
		WeightsStore7[405] <= Wgt_7_405;
		WeightsStore7[406] <= Wgt_7_406;
		WeightsStore7[407] <= Wgt_7_407;
		WeightsStore7[408] <= Wgt_7_408;
		WeightsStore7[409] <= Wgt_7_409;
		WeightsStore7[410] <= Wgt_7_410;
		WeightsStore7[411] <= Wgt_7_411;
		WeightsStore7[412] <= Wgt_7_412;
		WeightsStore7[413] <= Wgt_7_413;
		WeightsStore7[414] <= Wgt_7_414;
		WeightsStore7[415] <= Wgt_7_415;
		WeightsStore7[416] <= Wgt_7_416;
		WeightsStore7[417] <= Wgt_7_417;
		WeightsStore7[418] <= Wgt_7_418;
		WeightsStore7[419] <= Wgt_7_419;
		WeightsStore7[420] <= Wgt_7_420;
		WeightsStore7[421] <= Wgt_7_421;
		WeightsStore7[422] <= Wgt_7_422;
		WeightsStore7[423] <= Wgt_7_423;
		WeightsStore7[424] <= Wgt_7_424;
		WeightsStore7[425] <= Wgt_7_425;
		WeightsStore7[426] <= Wgt_7_426;
		WeightsStore7[427] <= Wgt_7_427;
		WeightsStore7[428] <= Wgt_7_428;
		WeightsStore7[429] <= Wgt_7_429;
		WeightsStore7[430] <= Wgt_7_430;
		WeightsStore7[431] <= Wgt_7_431;
		WeightsStore7[432] <= Wgt_7_432;
		WeightsStore7[433] <= Wgt_7_433;
		WeightsStore7[434] <= Wgt_7_434;
		WeightsStore7[435] <= Wgt_7_435;
		WeightsStore7[436] <= Wgt_7_436;
		WeightsStore7[437] <= Wgt_7_437;
		WeightsStore7[438] <= Wgt_7_438;
		WeightsStore7[439] <= Wgt_7_439;
		WeightsStore7[440] <= Wgt_7_440;
		WeightsStore7[441] <= Wgt_7_441;
		WeightsStore7[442] <= Wgt_7_442;
		WeightsStore7[443] <= Wgt_7_443;
		WeightsStore7[444] <= Wgt_7_444;
		WeightsStore7[445] <= Wgt_7_445;
		WeightsStore7[446] <= Wgt_7_446;
		WeightsStore7[447] <= Wgt_7_447;
		WeightsStore7[448] <= Wgt_7_448;
		WeightsStore7[449] <= Wgt_7_449;
		WeightsStore7[450] <= Wgt_7_450;
		WeightsStore7[451] <= Wgt_7_451;
		WeightsStore7[452] <= Wgt_7_452;
		WeightsStore7[453] <= Wgt_7_453;
		WeightsStore7[454] <= Wgt_7_454;
		WeightsStore7[455] <= Wgt_7_455;
		WeightsStore7[456] <= Wgt_7_456;
		WeightsStore7[457] <= Wgt_7_457;
		WeightsStore7[458] <= Wgt_7_458;
		WeightsStore7[459] <= Wgt_7_459;
		WeightsStore7[460] <= Wgt_7_460;
		WeightsStore7[461] <= Wgt_7_461;
		WeightsStore7[462] <= Wgt_7_462;
		WeightsStore7[463] <= Wgt_7_463;
		WeightsStore7[464] <= Wgt_7_464;
		WeightsStore7[465] <= Wgt_7_465;
		WeightsStore7[466] <= Wgt_7_466;
		WeightsStore7[467] <= Wgt_7_467;
		WeightsStore7[468] <= Wgt_7_468;
		WeightsStore7[469] <= Wgt_7_469;
		WeightsStore7[470] <= Wgt_7_470;
		WeightsStore7[471] <= Wgt_7_471;
		WeightsStore7[472] <= Wgt_7_472;
		WeightsStore7[473] <= Wgt_7_473;
		WeightsStore7[474] <= Wgt_7_474;
		WeightsStore7[475] <= Wgt_7_475;
		WeightsStore7[476] <= Wgt_7_476;
		WeightsStore7[477] <= Wgt_7_477;
		WeightsStore7[478] <= Wgt_7_478;
		WeightsStore7[479] <= Wgt_7_479;
		WeightsStore7[480] <= Wgt_7_480;
		WeightsStore7[481] <= Wgt_7_481;
		WeightsStore7[482] <= Wgt_7_482;
		WeightsStore7[483] <= Wgt_7_483;
		WeightsStore7[484] <= Wgt_7_484;
		WeightsStore7[485] <= Wgt_7_485;
		WeightsStore7[486] <= Wgt_7_486;
		WeightsStore7[487] <= Wgt_7_487;
		WeightsStore7[488] <= Wgt_7_488;
		WeightsStore7[489] <= Wgt_7_489;
		WeightsStore7[490] <= Wgt_7_490;
		WeightsStore7[491] <= Wgt_7_491;
		WeightsStore7[492] <= Wgt_7_492;
		WeightsStore7[493] <= Wgt_7_493;
		WeightsStore7[494] <= Wgt_7_494;
		WeightsStore7[495] <= Wgt_7_495;
		WeightsStore7[496] <= Wgt_7_496;
		WeightsStore7[497] <= Wgt_7_497;
		WeightsStore7[498] <= Wgt_7_498;
		WeightsStore7[499] <= Wgt_7_499;
		WeightsStore7[500] <= Wgt_7_500;
		WeightsStore7[501] <= Wgt_7_501;
		WeightsStore7[502] <= Wgt_7_502;
		WeightsStore7[503] <= Wgt_7_503;
		WeightsStore7[504] <= Wgt_7_504;
		WeightsStore7[505] <= Wgt_7_505;
		WeightsStore7[506] <= Wgt_7_506;
		WeightsStore7[507] <= Wgt_7_507;
		WeightsStore7[508] <= Wgt_7_508;
		WeightsStore7[509] <= Wgt_7_509;
		WeightsStore7[510] <= Wgt_7_510;
		WeightsStore7[511] <= Wgt_7_511;
		WeightsStore7[512] <= Wgt_7_512;
		WeightsStore7[513] <= Wgt_7_513;
		WeightsStore7[514] <= Wgt_7_514;
		WeightsStore7[515] <= Wgt_7_515;
		WeightsStore7[516] <= Wgt_7_516;
		WeightsStore7[517] <= Wgt_7_517;
		WeightsStore7[518] <= Wgt_7_518;
		WeightsStore7[519] <= Wgt_7_519;
		WeightsStore7[520] <= Wgt_7_520;
		WeightsStore7[521] <= Wgt_7_521;
		WeightsStore7[522] <= Wgt_7_522;
		WeightsStore7[523] <= Wgt_7_523;
		WeightsStore7[524] <= Wgt_7_524;
		WeightsStore7[525] <= Wgt_7_525;
		WeightsStore7[526] <= Wgt_7_526;
		WeightsStore7[527] <= Wgt_7_527;
		WeightsStore7[528] <= Wgt_7_528;
		WeightsStore7[529] <= Wgt_7_529;
		WeightsStore7[530] <= Wgt_7_530;
		WeightsStore7[531] <= Wgt_7_531;
		WeightsStore7[532] <= Wgt_7_532;
		WeightsStore7[533] <= Wgt_7_533;
		WeightsStore7[534] <= Wgt_7_534;
		WeightsStore7[535] <= Wgt_7_535;
		WeightsStore7[536] <= Wgt_7_536;
		WeightsStore7[537] <= Wgt_7_537;
		WeightsStore7[538] <= Wgt_7_538;
		WeightsStore7[539] <= Wgt_7_539;
		WeightsStore7[540] <= Wgt_7_540;
		WeightsStore7[541] <= Wgt_7_541;
		WeightsStore7[542] <= Wgt_7_542;
		WeightsStore7[543] <= Wgt_7_543;
		WeightsStore7[544] <= Wgt_7_544;
		WeightsStore7[545] <= Wgt_7_545;
		WeightsStore7[546] <= Wgt_7_546;
		WeightsStore7[547] <= Wgt_7_547;
		WeightsStore7[548] <= Wgt_7_548;
		WeightsStore7[549] <= Wgt_7_549;
		WeightsStore7[550] <= Wgt_7_550;
		WeightsStore7[551] <= Wgt_7_551;
		WeightsStore7[552] <= Wgt_7_552;
		WeightsStore7[553] <= Wgt_7_553;
		WeightsStore7[554] <= Wgt_7_554;
		WeightsStore7[555] <= Wgt_7_555;
		WeightsStore7[556] <= Wgt_7_556;
		WeightsStore7[557] <= Wgt_7_557;
		WeightsStore7[558] <= Wgt_7_558;
		WeightsStore7[559] <= Wgt_7_559;
		WeightsStore7[560] <= Wgt_7_560;
		WeightsStore7[561] <= Wgt_7_561;
		WeightsStore7[562] <= Wgt_7_562;
		WeightsStore7[563] <= Wgt_7_563;
		WeightsStore7[564] <= Wgt_7_564;
		WeightsStore7[565] <= Wgt_7_565;
		WeightsStore7[566] <= Wgt_7_566;
		WeightsStore7[567] <= Wgt_7_567;
		WeightsStore7[568] <= Wgt_7_568;
		WeightsStore7[569] <= Wgt_7_569;
		WeightsStore7[570] <= Wgt_7_570;
		WeightsStore7[571] <= Wgt_7_571;
		WeightsStore7[572] <= Wgt_7_572;
		WeightsStore7[573] <= Wgt_7_573;
		WeightsStore7[574] <= Wgt_7_574;
		WeightsStore7[575] <= Wgt_7_575;
		WeightsStore7[576] <= Wgt_7_576;
		WeightsStore7[577] <= Wgt_7_577;
		WeightsStore7[578] <= Wgt_7_578;
		WeightsStore7[579] <= Wgt_7_579;
		WeightsStore7[580] <= Wgt_7_580;
		WeightsStore7[581] <= Wgt_7_581;
		WeightsStore7[582] <= Wgt_7_582;
		WeightsStore7[583] <= Wgt_7_583;
		WeightsStore7[584] <= Wgt_7_584;
		WeightsStore7[585] <= Wgt_7_585;
		WeightsStore7[586] <= Wgt_7_586;
		WeightsStore7[587] <= Wgt_7_587;
		WeightsStore7[588] <= Wgt_7_588;
		WeightsStore7[589] <= Wgt_7_589;
		WeightsStore7[590] <= Wgt_7_590;
		WeightsStore7[591] <= Wgt_7_591;
		WeightsStore7[592] <= Wgt_7_592;
		WeightsStore7[593] <= Wgt_7_593;
		WeightsStore7[594] <= Wgt_7_594;
		WeightsStore7[595] <= Wgt_7_595;
		WeightsStore7[596] <= Wgt_7_596;
		WeightsStore7[597] <= Wgt_7_597;
		WeightsStore7[598] <= Wgt_7_598;
		WeightsStore7[599] <= Wgt_7_599;
		WeightsStore7[600] <= Wgt_7_600;
		WeightsStore7[601] <= Wgt_7_601;
		WeightsStore7[602] <= Wgt_7_602;
		WeightsStore7[603] <= Wgt_7_603;
		WeightsStore7[604] <= Wgt_7_604;
		WeightsStore7[605] <= Wgt_7_605;
		WeightsStore7[606] <= Wgt_7_606;
		WeightsStore7[607] <= Wgt_7_607;
		WeightsStore7[608] <= Wgt_7_608;
		WeightsStore7[609] <= Wgt_7_609;
		WeightsStore7[610] <= Wgt_7_610;
		WeightsStore7[611] <= Wgt_7_611;
		WeightsStore7[612] <= Wgt_7_612;
		WeightsStore7[613] <= Wgt_7_613;
		WeightsStore7[614] <= Wgt_7_614;
		WeightsStore7[615] <= Wgt_7_615;
		WeightsStore7[616] <= Wgt_7_616;
		WeightsStore7[617] <= Wgt_7_617;
		WeightsStore7[618] <= Wgt_7_618;
		WeightsStore7[619] <= Wgt_7_619;
		WeightsStore7[620] <= Wgt_7_620;
		WeightsStore7[621] <= Wgt_7_621;
		WeightsStore7[622] <= Wgt_7_622;
		WeightsStore7[623] <= Wgt_7_623;
		WeightsStore7[624] <= Wgt_7_624;
		WeightsStore7[625] <= Wgt_7_625;
		WeightsStore7[626] <= Wgt_7_626;
		WeightsStore7[627] <= Wgt_7_627;
		WeightsStore7[628] <= Wgt_7_628;
		WeightsStore7[629] <= Wgt_7_629;
		WeightsStore7[630] <= Wgt_7_630;
		WeightsStore7[631] <= Wgt_7_631;
		WeightsStore7[632] <= Wgt_7_632;
		WeightsStore7[633] <= Wgt_7_633;
		WeightsStore7[634] <= Wgt_7_634;
		WeightsStore7[635] <= Wgt_7_635;
		WeightsStore7[636] <= Wgt_7_636;
		WeightsStore7[637] <= Wgt_7_637;
		WeightsStore7[638] <= Wgt_7_638;
		WeightsStore7[639] <= Wgt_7_639;
		WeightsStore7[640] <= Wgt_7_640;
		WeightsStore7[641] <= Wgt_7_641;
		WeightsStore7[642] <= Wgt_7_642;
		WeightsStore7[643] <= Wgt_7_643;
		WeightsStore7[644] <= Wgt_7_644;
		WeightsStore7[645] <= Wgt_7_645;
		WeightsStore7[646] <= Wgt_7_646;
		WeightsStore7[647] <= Wgt_7_647;
		WeightsStore7[648] <= Wgt_7_648;
		WeightsStore7[649] <= Wgt_7_649;
		WeightsStore7[650] <= Wgt_7_650;
		WeightsStore7[651] <= Wgt_7_651;
		WeightsStore7[652] <= Wgt_7_652;
		WeightsStore7[653] <= Wgt_7_653;
		WeightsStore7[654] <= Wgt_7_654;
		WeightsStore7[655] <= Wgt_7_655;
		WeightsStore7[656] <= Wgt_7_656;
		WeightsStore7[657] <= Wgt_7_657;
		WeightsStore7[658] <= Wgt_7_658;
		WeightsStore7[659] <= Wgt_7_659;
		WeightsStore7[660] <= Wgt_7_660;
		WeightsStore7[661] <= Wgt_7_661;
		WeightsStore7[662] <= Wgt_7_662;
		WeightsStore7[663] <= Wgt_7_663;
		WeightsStore7[664] <= Wgt_7_664;
		WeightsStore7[665] <= Wgt_7_665;
		WeightsStore7[666] <= Wgt_7_666;
		WeightsStore7[667] <= Wgt_7_667;
		WeightsStore7[668] <= Wgt_7_668;
		WeightsStore7[669] <= Wgt_7_669;
		WeightsStore7[670] <= Wgt_7_670;
		WeightsStore7[671] <= Wgt_7_671;
		WeightsStore7[672] <= Wgt_7_672;
		WeightsStore7[673] <= Wgt_7_673;
		WeightsStore7[674] <= Wgt_7_674;
		WeightsStore7[675] <= Wgt_7_675;
		WeightsStore7[676] <= Wgt_7_676;
		WeightsStore7[677] <= Wgt_7_677;
		WeightsStore7[678] <= Wgt_7_678;
		WeightsStore7[679] <= Wgt_7_679;
		WeightsStore7[680] <= Wgt_7_680;
		WeightsStore7[681] <= Wgt_7_681;
		WeightsStore7[682] <= Wgt_7_682;
		WeightsStore7[683] <= Wgt_7_683;
		WeightsStore7[684] <= Wgt_7_684;
		WeightsStore7[685] <= Wgt_7_685;
		WeightsStore7[686] <= Wgt_7_686;
		WeightsStore7[687] <= Wgt_7_687;
		WeightsStore7[688] <= Wgt_7_688;
		WeightsStore7[689] <= Wgt_7_689;
		WeightsStore7[690] <= Wgt_7_690;
		WeightsStore7[691] <= Wgt_7_691;
		WeightsStore7[692] <= Wgt_7_692;
		WeightsStore7[693] <= Wgt_7_693;
		WeightsStore7[694] <= Wgt_7_694;
		WeightsStore7[695] <= Wgt_7_695;
		WeightsStore7[696] <= Wgt_7_696;
		WeightsStore7[697] <= Wgt_7_697;
		WeightsStore7[698] <= Wgt_7_698;
		WeightsStore7[699] <= Wgt_7_699;
		WeightsStore7[700] <= Wgt_7_700;
		WeightsStore7[701] <= Wgt_7_701;
		WeightsStore7[702] <= Wgt_7_702;
		WeightsStore7[703] <= Wgt_7_703;
		WeightsStore7[704] <= Wgt_7_704;
		WeightsStore7[705] <= Wgt_7_705;
		WeightsStore7[706] <= Wgt_7_706;
		WeightsStore7[707] <= Wgt_7_707;
		WeightsStore7[708] <= Wgt_7_708;
		WeightsStore7[709] <= Wgt_7_709;
		WeightsStore7[710] <= Wgt_7_710;
		WeightsStore7[711] <= Wgt_7_711;
		WeightsStore7[712] <= Wgt_7_712;
		WeightsStore7[713] <= Wgt_7_713;
		WeightsStore7[714] <= Wgt_7_714;
		WeightsStore7[715] <= Wgt_7_715;
		WeightsStore7[716] <= Wgt_7_716;
		WeightsStore7[717] <= Wgt_7_717;
		WeightsStore7[718] <= Wgt_7_718;
		WeightsStore7[719] <= Wgt_7_719;
		WeightsStore7[720] <= Wgt_7_720;
		WeightsStore7[721] <= Wgt_7_721;
		WeightsStore7[722] <= Wgt_7_722;
		WeightsStore7[723] <= Wgt_7_723;
		WeightsStore7[724] <= Wgt_7_724;
		WeightsStore7[725] <= Wgt_7_725;
		WeightsStore7[726] <= Wgt_7_726;
		WeightsStore7[727] <= Wgt_7_727;
		WeightsStore7[728] <= Wgt_7_728;
		WeightsStore7[729] <= Wgt_7_729;
		WeightsStore7[730] <= Wgt_7_730;
		WeightsStore7[731] <= Wgt_7_731;
		WeightsStore7[732] <= Wgt_7_732;
		WeightsStore7[733] <= Wgt_7_733;
		WeightsStore7[734] <= Wgt_7_734;
		WeightsStore7[735] <= Wgt_7_735;
		WeightsStore7[736] <= Wgt_7_736;
		WeightsStore7[737] <= Wgt_7_737;
		WeightsStore7[738] <= Wgt_7_738;
		WeightsStore7[739] <= Wgt_7_739;
		WeightsStore7[740] <= Wgt_7_740;
		WeightsStore7[741] <= Wgt_7_741;
		WeightsStore7[742] <= Wgt_7_742;
		WeightsStore7[743] <= Wgt_7_743;
		WeightsStore7[744] <= Wgt_7_744;
		WeightsStore7[745] <= Wgt_7_745;
		WeightsStore7[746] <= Wgt_7_746;
		WeightsStore7[747] <= Wgt_7_747;
		WeightsStore7[748] <= Wgt_7_748;
		WeightsStore7[749] <= Wgt_7_749;
		WeightsStore7[750] <= Wgt_7_750;
		WeightsStore7[751] <= Wgt_7_751;
		WeightsStore7[752] <= Wgt_7_752;
		WeightsStore7[753] <= Wgt_7_753;
		WeightsStore7[754] <= Wgt_7_754;
		WeightsStore7[755] <= Wgt_7_755;
		WeightsStore7[756] <= Wgt_7_756;
		WeightsStore7[757] <= Wgt_7_757;
		WeightsStore7[758] <= Wgt_7_758;
		WeightsStore7[759] <= Wgt_7_759;
		WeightsStore7[760] <= Wgt_7_760;
		WeightsStore7[761] <= Wgt_7_761;
		WeightsStore7[762] <= Wgt_7_762;
		WeightsStore7[763] <= Wgt_7_763;
		WeightsStore7[764] <= Wgt_7_764;
		WeightsStore7[765] <= Wgt_7_765;
		WeightsStore7[766] <= Wgt_7_766;
		WeightsStore7[767] <= Wgt_7_767;
		WeightsStore7[768] <= Wgt_7_768;
		WeightsStore7[769] <= Wgt_7_769;
		WeightsStore7[770] <= Wgt_7_770;
		WeightsStore7[771] <= Wgt_7_771;
		WeightsStore7[772] <= Wgt_7_772;
		WeightsStore7[773] <= Wgt_7_773;
		WeightsStore7[774] <= Wgt_7_774;
		WeightsStore7[775] <= Wgt_7_775;
		WeightsStore7[776] <= Wgt_7_776;
		WeightsStore7[777] <= Wgt_7_777;
		WeightsStore7[778] <= Wgt_7_778;
		WeightsStore7[779] <= Wgt_7_779;
		WeightsStore7[780] <= Wgt_7_780;
		WeightsStore7[781] <= Wgt_7_781;
		WeightsStore7[782] <= Wgt_7_782;
		WeightsStore7[783] <= Wgt_7_783;
		WeightsStore7[784] <= Wgt_7_784;
		WeightsStore8[0] <= Wgt_8_0;
		WeightsStore8[1] <= Wgt_8_1;
		WeightsStore8[2] <= Wgt_8_2;
		WeightsStore8[3] <= Wgt_8_3;
		WeightsStore8[4] <= Wgt_8_4;
		WeightsStore8[5] <= Wgt_8_5;
		WeightsStore8[6] <= Wgt_8_6;
		WeightsStore8[7] <= Wgt_8_7;
		WeightsStore8[8] <= Wgt_8_8;
		WeightsStore8[9] <= Wgt_8_9;
		WeightsStore8[10] <= Wgt_8_10;
		WeightsStore8[11] <= Wgt_8_11;
		WeightsStore8[12] <= Wgt_8_12;
		WeightsStore8[13] <= Wgt_8_13;
		WeightsStore8[14] <= Wgt_8_14;
		WeightsStore8[15] <= Wgt_8_15;
		WeightsStore8[16] <= Wgt_8_16;
		WeightsStore8[17] <= Wgt_8_17;
		WeightsStore8[18] <= Wgt_8_18;
		WeightsStore8[19] <= Wgt_8_19;
		WeightsStore8[20] <= Wgt_8_20;
		WeightsStore8[21] <= Wgt_8_21;
		WeightsStore8[22] <= Wgt_8_22;
		WeightsStore8[23] <= Wgt_8_23;
		WeightsStore8[24] <= Wgt_8_24;
		WeightsStore8[25] <= Wgt_8_25;
		WeightsStore8[26] <= Wgt_8_26;
		WeightsStore8[27] <= Wgt_8_27;
		WeightsStore8[28] <= Wgt_8_28;
		WeightsStore8[29] <= Wgt_8_29;
		WeightsStore8[30] <= Wgt_8_30;
		WeightsStore8[31] <= Wgt_8_31;
		WeightsStore8[32] <= Wgt_8_32;
		WeightsStore8[33] <= Wgt_8_33;
		WeightsStore8[34] <= Wgt_8_34;
		WeightsStore8[35] <= Wgt_8_35;
		WeightsStore8[36] <= Wgt_8_36;
		WeightsStore8[37] <= Wgt_8_37;
		WeightsStore8[38] <= Wgt_8_38;
		WeightsStore8[39] <= Wgt_8_39;
		WeightsStore8[40] <= Wgt_8_40;
		WeightsStore8[41] <= Wgt_8_41;
		WeightsStore8[42] <= Wgt_8_42;
		WeightsStore8[43] <= Wgt_8_43;
		WeightsStore8[44] <= Wgt_8_44;
		WeightsStore8[45] <= Wgt_8_45;
		WeightsStore8[46] <= Wgt_8_46;
		WeightsStore8[47] <= Wgt_8_47;
		WeightsStore8[48] <= Wgt_8_48;
		WeightsStore8[49] <= Wgt_8_49;
		WeightsStore8[50] <= Wgt_8_50;
		WeightsStore8[51] <= Wgt_8_51;
		WeightsStore8[52] <= Wgt_8_52;
		WeightsStore8[53] <= Wgt_8_53;
		WeightsStore8[54] <= Wgt_8_54;
		WeightsStore8[55] <= Wgt_8_55;
		WeightsStore8[56] <= Wgt_8_56;
		WeightsStore8[57] <= Wgt_8_57;
		WeightsStore8[58] <= Wgt_8_58;
		WeightsStore8[59] <= Wgt_8_59;
		WeightsStore8[60] <= Wgt_8_60;
		WeightsStore8[61] <= Wgt_8_61;
		WeightsStore8[62] <= Wgt_8_62;
		WeightsStore8[63] <= Wgt_8_63;
		WeightsStore8[64] <= Wgt_8_64;
		WeightsStore8[65] <= Wgt_8_65;
		WeightsStore8[66] <= Wgt_8_66;
		WeightsStore8[67] <= Wgt_8_67;
		WeightsStore8[68] <= Wgt_8_68;
		WeightsStore8[69] <= Wgt_8_69;
		WeightsStore8[70] <= Wgt_8_70;
		WeightsStore8[71] <= Wgt_8_71;
		WeightsStore8[72] <= Wgt_8_72;
		WeightsStore8[73] <= Wgt_8_73;
		WeightsStore8[74] <= Wgt_8_74;
		WeightsStore8[75] <= Wgt_8_75;
		WeightsStore8[76] <= Wgt_8_76;
		WeightsStore8[77] <= Wgt_8_77;
		WeightsStore8[78] <= Wgt_8_78;
		WeightsStore8[79] <= Wgt_8_79;
		WeightsStore8[80] <= Wgt_8_80;
		WeightsStore8[81] <= Wgt_8_81;
		WeightsStore8[82] <= Wgt_8_82;
		WeightsStore8[83] <= Wgt_8_83;
		WeightsStore8[84] <= Wgt_8_84;
		WeightsStore8[85] <= Wgt_8_85;
		WeightsStore8[86] <= Wgt_8_86;
		WeightsStore8[87] <= Wgt_8_87;
		WeightsStore8[88] <= Wgt_8_88;
		WeightsStore8[89] <= Wgt_8_89;
		WeightsStore8[90] <= Wgt_8_90;
		WeightsStore8[91] <= Wgt_8_91;
		WeightsStore8[92] <= Wgt_8_92;
		WeightsStore8[93] <= Wgt_8_93;
		WeightsStore8[94] <= Wgt_8_94;
		WeightsStore8[95] <= Wgt_8_95;
		WeightsStore8[96] <= Wgt_8_96;
		WeightsStore8[97] <= Wgt_8_97;
		WeightsStore8[98] <= Wgt_8_98;
		WeightsStore8[99] <= Wgt_8_99;
		WeightsStore8[100] <= Wgt_8_100;
		WeightsStore8[101] <= Wgt_8_101;
		WeightsStore8[102] <= Wgt_8_102;
		WeightsStore8[103] <= Wgt_8_103;
		WeightsStore8[104] <= Wgt_8_104;
		WeightsStore8[105] <= Wgt_8_105;
		WeightsStore8[106] <= Wgt_8_106;
		WeightsStore8[107] <= Wgt_8_107;
		WeightsStore8[108] <= Wgt_8_108;
		WeightsStore8[109] <= Wgt_8_109;
		WeightsStore8[110] <= Wgt_8_110;
		WeightsStore8[111] <= Wgt_8_111;
		WeightsStore8[112] <= Wgt_8_112;
		WeightsStore8[113] <= Wgt_8_113;
		WeightsStore8[114] <= Wgt_8_114;
		WeightsStore8[115] <= Wgt_8_115;
		WeightsStore8[116] <= Wgt_8_116;
		WeightsStore8[117] <= Wgt_8_117;
		WeightsStore8[118] <= Wgt_8_118;
		WeightsStore8[119] <= Wgt_8_119;
		WeightsStore8[120] <= Wgt_8_120;
		WeightsStore8[121] <= Wgt_8_121;
		WeightsStore8[122] <= Wgt_8_122;
		WeightsStore8[123] <= Wgt_8_123;
		WeightsStore8[124] <= Wgt_8_124;
		WeightsStore8[125] <= Wgt_8_125;
		WeightsStore8[126] <= Wgt_8_126;
		WeightsStore8[127] <= Wgt_8_127;
		WeightsStore8[128] <= Wgt_8_128;
		WeightsStore8[129] <= Wgt_8_129;
		WeightsStore8[130] <= Wgt_8_130;
		WeightsStore8[131] <= Wgt_8_131;
		WeightsStore8[132] <= Wgt_8_132;
		WeightsStore8[133] <= Wgt_8_133;
		WeightsStore8[134] <= Wgt_8_134;
		WeightsStore8[135] <= Wgt_8_135;
		WeightsStore8[136] <= Wgt_8_136;
		WeightsStore8[137] <= Wgt_8_137;
		WeightsStore8[138] <= Wgt_8_138;
		WeightsStore8[139] <= Wgt_8_139;
		WeightsStore8[140] <= Wgt_8_140;
		WeightsStore8[141] <= Wgt_8_141;
		WeightsStore8[142] <= Wgt_8_142;
		WeightsStore8[143] <= Wgt_8_143;
		WeightsStore8[144] <= Wgt_8_144;
		WeightsStore8[145] <= Wgt_8_145;
		WeightsStore8[146] <= Wgt_8_146;
		WeightsStore8[147] <= Wgt_8_147;
		WeightsStore8[148] <= Wgt_8_148;
		WeightsStore8[149] <= Wgt_8_149;
		WeightsStore8[150] <= Wgt_8_150;
		WeightsStore8[151] <= Wgt_8_151;
		WeightsStore8[152] <= Wgt_8_152;
		WeightsStore8[153] <= Wgt_8_153;
		WeightsStore8[154] <= Wgt_8_154;
		WeightsStore8[155] <= Wgt_8_155;
		WeightsStore8[156] <= Wgt_8_156;
		WeightsStore8[157] <= Wgt_8_157;
		WeightsStore8[158] <= Wgt_8_158;
		WeightsStore8[159] <= Wgt_8_159;
		WeightsStore8[160] <= Wgt_8_160;
		WeightsStore8[161] <= Wgt_8_161;
		WeightsStore8[162] <= Wgt_8_162;
		WeightsStore8[163] <= Wgt_8_163;
		WeightsStore8[164] <= Wgt_8_164;
		WeightsStore8[165] <= Wgt_8_165;
		WeightsStore8[166] <= Wgt_8_166;
		WeightsStore8[167] <= Wgt_8_167;
		WeightsStore8[168] <= Wgt_8_168;
		WeightsStore8[169] <= Wgt_8_169;
		WeightsStore8[170] <= Wgt_8_170;
		WeightsStore8[171] <= Wgt_8_171;
		WeightsStore8[172] <= Wgt_8_172;
		WeightsStore8[173] <= Wgt_8_173;
		WeightsStore8[174] <= Wgt_8_174;
		WeightsStore8[175] <= Wgt_8_175;
		WeightsStore8[176] <= Wgt_8_176;
		WeightsStore8[177] <= Wgt_8_177;
		WeightsStore8[178] <= Wgt_8_178;
		WeightsStore8[179] <= Wgt_8_179;
		WeightsStore8[180] <= Wgt_8_180;
		WeightsStore8[181] <= Wgt_8_181;
		WeightsStore8[182] <= Wgt_8_182;
		WeightsStore8[183] <= Wgt_8_183;
		WeightsStore8[184] <= Wgt_8_184;
		WeightsStore8[185] <= Wgt_8_185;
		WeightsStore8[186] <= Wgt_8_186;
		WeightsStore8[187] <= Wgt_8_187;
		WeightsStore8[188] <= Wgt_8_188;
		WeightsStore8[189] <= Wgt_8_189;
		WeightsStore8[190] <= Wgt_8_190;
		WeightsStore8[191] <= Wgt_8_191;
		WeightsStore8[192] <= Wgt_8_192;
		WeightsStore8[193] <= Wgt_8_193;
		WeightsStore8[194] <= Wgt_8_194;
		WeightsStore8[195] <= Wgt_8_195;
		WeightsStore8[196] <= Wgt_8_196;
		WeightsStore8[197] <= Wgt_8_197;
		WeightsStore8[198] <= Wgt_8_198;
		WeightsStore8[199] <= Wgt_8_199;
		WeightsStore8[200] <= Wgt_8_200;
		WeightsStore8[201] <= Wgt_8_201;
		WeightsStore8[202] <= Wgt_8_202;
		WeightsStore8[203] <= Wgt_8_203;
		WeightsStore8[204] <= Wgt_8_204;
		WeightsStore8[205] <= Wgt_8_205;
		WeightsStore8[206] <= Wgt_8_206;
		WeightsStore8[207] <= Wgt_8_207;
		WeightsStore8[208] <= Wgt_8_208;
		WeightsStore8[209] <= Wgt_8_209;
		WeightsStore8[210] <= Wgt_8_210;
		WeightsStore8[211] <= Wgt_8_211;
		WeightsStore8[212] <= Wgt_8_212;
		WeightsStore8[213] <= Wgt_8_213;
		WeightsStore8[214] <= Wgt_8_214;
		WeightsStore8[215] <= Wgt_8_215;
		WeightsStore8[216] <= Wgt_8_216;
		WeightsStore8[217] <= Wgt_8_217;
		WeightsStore8[218] <= Wgt_8_218;
		WeightsStore8[219] <= Wgt_8_219;
		WeightsStore8[220] <= Wgt_8_220;
		WeightsStore8[221] <= Wgt_8_221;
		WeightsStore8[222] <= Wgt_8_222;
		WeightsStore8[223] <= Wgt_8_223;
		WeightsStore8[224] <= Wgt_8_224;
		WeightsStore8[225] <= Wgt_8_225;
		WeightsStore8[226] <= Wgt_8_226;
		WeightsStore8[227] <= Wgt_8_227;
		WeightsStore8[228] <= Wgt_8_228;
		WeightsStore8[229] <= Wgt_8_229;
		WeightsStore8[230] <= Wgt_8_230;
		WeightsStore8[231] <= Wgt_8_231;
		WeightsStore8[232] <= Wgt_8_232;
		WeightsStore8[233] <= Wgt_8_233;
		WeightsStore8[234] <= Wgt_8_234;
		WeightsStore8[235] <= Wgt_8_235;
		WeightsStore8[236] <= Wgt_8_236;
		WeightsStore8[237] <= Wgt_8_237;
		WeightsStore8[238] <= Wgt_8_238;
		WeightsStore8[239] <= Wgt_8_239;
		WeightsStore8[240] <= Wgt_8_240;
		WeightsStore8[241] <= Wgt_8_241;
		WeightsStore8[242] <= Wgt_8_242;
		WeightsStore8[243] <= Wgt_8_243;
		WeightsStore8[244] <= Wgt_8_244;
		WeightsStore8[245] <= Wgt_8_245;
		WeightsStore8[246] <= Wgt_8_246;
		WeightsStore8[247] <= Wgt_8_247;
		WeightsStore8[248] <= Wgt_8_248;
		WeightsStore8[249] <= Wgt_8_249;
		WeightsStore8[250] <= Wgt_8_250;
		WeightsStore8[251] <= Wgt_8_251;
		WeightsStore8[252] <= Wgt_8_252;
		WeightsStore8[253] <= Wgt_8_253;
		WeightsStore8[254] <= Wgt_8_254;
		WeightsStore8[255] <= Wgt_8_255;
		WeightsStore8[256] <= Wgt_8_256;
		WeightsStore8[257] <= Wgt_8_257;
		WeightsStore8[258] <= Wgt_8_258;
		WeightsStore8[259] <= Wgt_8_259;
		WeightsStore8[260] <= Wgt_8_260;
		WeightsStore8[261] <= Wgt_8_261;
		WeightsStore8[262] <= Wgt_8_262;
		WeightsStore8[263] <= Wgt_8_263;
		WeightsStore8[264] <= Wgt_8_264;
		WeightsStore8[265] <= Wgt_8_265;
		WeightsStore8[266] <= Wgt_8_266;
		WeightsStore8[267] <= Wgt_8_267;
		WeightsStore8[268] <= Wgt_8_268;
		WeightsStore8[269] <= Wgt_8_269;
		WeightsStore8[270] <= Wgt_8_270;
		WeightsStore8[271] <= Wgt_8_271;
		WeightsStore8[272] <= Wgt_8_272;
		WeightsStore8[273] <= Wgt_8_273;
		WeightsStore8[274] <= Wgt_8_274;
		WeightsStore8[275] <= Wgt_8_275;
		WeightsStore8[276] <= Wgt_8_276;
		WeightsStore8[277] <= Wgt_8_277;
		WeightsStore8[278] <= Wgt_8_278;
		WeightsStore8[279] <= Wgt_8_279;
		WeightsStore8[280] <= Wgt_8_280;
		WeightsStore8[281] <= Wgt_8_281;
		WeightsStore8[282] <= Wgt_8_282;
		WeightsStore8[283] <= Wgt_8_283;
		WeightsStore8[284] <= Wgt_8_284;
		WeightsStore8[285] <= Wgt_8_285;
		WeightsStore8[286] <= Wgt_8_286;
		WeightsStore8[287] <= Wgt_8_287;
		WeightsStore8[288] <= Wgt_8_288;
		WeightsStore8[289] <= Wgt_8_289;
		WeightsStore8[290] <= Wgt_8_290;
		WeightsStore8[291] <= Wgt_8_291;
		WeightsStore8[292] <= Wgt_8_292;
		WeightsStore8[293] <= Wgt_8_293;
		WeightsStore8[294] <= Wgt_8_294;
		WeightsStore8[295] <= Wgt_8_295;
		WeightsStore8[296] <= Wgt_8_296;
		WeightsStore8[297] <= Wgt_8_297;
		WeightsStore8[298] <= Wgt_8_298;
		WeightsStore8[299] <= Wgt_8_299;
		WeightsStore8[300] <= Wgt_8_300;
		WeightsStore8[301] <= Wgt_8_301;
		WeightsStore8[302] <= Wgt_8_302;
		WeightsStore8[303] <= Wgt_8_303;
		WeightsStore8[304] <= Wgt_8_304;
		WeightsStore8[305] <= Wgt_8_305;
		WeightsStore8[306] <= Wgt_8_306;
		WeightsStore8[307] <= Wgt_8_307;
		WeightsStore8[308] <= Wgt_8_308;
		WeightsStore8[309] <= Wgt_8_309;
		WeightsStore8[310] <= Wgt_8_310;
		WeightsStore8[311] <= Wgt_8_311;
		WeightsStore8[312] <= Wgt_8_312;
		WeightsStore8[313] <= Wgt_8_313;
		WeightsStore8[314] <= Wgt_8_314;
		WeightsStore8[315] <= Wgt_8_315;
		WeightsStore8[316] <= Wgt_8_316;
		WeightsStore8[317] <= Wgt_8_317;
		WeightsStore8[318] <= Wgt_8_318;
		WeightsStore8[319] <= Wgt_8_319;
		WeightsStore8[320] <= Wgt_8_320;
		WeightsStore8[321] <= Wgt_8_321;
		WeightsStore8[322] <= Wgt_8_322;
		WeightsStore8[323] <= Wgt_8_323;
		WeightsStore8[324] <= Wgt_8_324;
		WeightsStore8[325] <= Wgt_8_325;
		WeightsStore8[326] <= Wgt_8_326;
		WeightsStore8[327] <= Wgt_8_327;
		WeightsStore8[328] <= Wgt_8_328;
		WeightsStore8[329] <= Wgt_8_329;
		WeightsStore8[330] <= Wgt_8_330;
		WeightsStore8[331] <= Wgt_8_331;
		WeightsStore8[332] <= Wgt_8_332;
		WeightsStore8[333] <= Wgt_8_333;
		WeightsStore8[334] <= Wgt_8_334;
		WeightsStore8[335] <= Wgt_8_335;
		WeightsStore8[336] <= Wgt_8_336;
		WeightsStore8[337] <= Wgt_8_337;
		WeightsStore8[338] <= Wgt_8_338;
		WeightsStore8[339] <= Wgt_8_339;
		WeightsStore8[340] <= Wgt_8_340;
		WeightsStore8[341] <= Wgt_8_341;
		WeightsStore8[342] <= Wgt_8_342;
		WeightsStore8[343] <= Wgt_8_343;
		WeightsStore8[344] <= Wgt_8_344;
		WeightsStore8[345] <= Wgt_8_345;
		WeightsStore8[346] <= Wgt_8_346;
		WeightsStore8[347] <= Wgt_8_347;
		WeightsStore8[348] <= Wgt_8_348;
		WeightsStore8[349] <= Wgt_8_349;
		WeightsStore8[350] <= Wgt_8_350;
		WeightsStore8[351] <= Wgt_8_351;
		WeightsStore8[352] <= Wgt_8_352;
		WeightsStore8[353] <= Wgt_8_353;
		WeightsStore8[354] <= Wgt_8_354;
		WeightsStore8[355] <= Wgt_8_355;
		WeightsStore8[356] <= Wgt_8_356;
		WeightsStore8[357] <= Wgt_8_357;
		WeightsStore8[358] <= Wgt_8_358;
		WeightsStore8[359] <= Wgt_8_359;
		WeightsStore8[360] <= Wgt_8_360;
		WeightsStore8[361] <= Wgt_8_361;
		WeightsStore8[362] <= Wgt_8_362;
		WeightsStore8[363] <= Wgt_8_363;
		WeightsStore8[364] <= Wgt_8_364;
		WeightsStore8[365] <= Wgt_8_365;
		WeightsStore8[366] <= Wgt_8_366;
		WeightsStore8[367] <= Wgt_8_367;
		WeightsStore8[368] <= Wgt_8_368;
		WeightsStore8[369] <= Wgt_8_369;
		WeightsStore8[370] <= Wgt_8_370;
		WeightsStore8[371] <= Wgt_8_371;
		WeightsStore8[372] <= Wgt_8_372;
		WeightsStore8[373] <= Wgt_8_373;
		WeightsStore8[374] <= Wgt_8_374;
		WeightsStore8[375] <= Wgt_8_375;
		WeightsStore8[376] <= Wgt_8_376;
		WeightsStore8[377] <= Wgt_8_377;
		WeightsStore8[378] <= Wgt_8_378;
		WeightsStore8[379] <= Wgt_8_379;
		WeightsStore8[380] <= Wgt_8_380;
		WeightsStore8[381] <= Wgt_8_381;
		WeightsStore8[382] <= Wgt_8_382;
		WeightsStore8[383] <= Wgt_8_383;
		WeightsStore8[384] <= Wgt_8_384;
		WeightsStore8[385] <= Wgt_8_385;
		WeightsStore8[386] <= Wgt_8_386;
		WeightsStore8[387] <= Wgt_8_387;
		WeightsStore8[388] <= Wgt_8_388;
		WeightsStore8[389] <= Wgt_8_389;
		WeightsStore8[390] <= Wgt_8_390;
		WeightsStore8[391] <= Wgt_8_391;
		WeightsStore8[392] <= Wgt_8_392;
		WeightsStore8[393] <= Wgt_8_393;
		WeightsStore8[394] <= Wgt_8_394;
		WeightsStore8[395] <= Wgt_8_395;
		WeightsStore8[396] <= Wgt_8_396;
		WeightsStore8[397] <= Wgt_8_397;
		WeightsStore8[398] <= Wgt_8_398;
		WeightsStore8[399] <= Wgt_8_399;
		WeightsStore8[400] <= Wgt_8_400;
		WeightsStore8[401] <= Wgt_8_401;
		WeightsStore8[402] <= Wgt_8_402;
		WeightsStore8[403] <= Wgt_8_403;
		WeightsStore8[404] <= Wgt_8_404;
		WeightsStore8[405] <= Wgt_8_405;
		WeightsStore8[406] <= Wgt_8_406;
		WeightsStore8[407] <= Wgt_8_407;
		WeightsStore8[408] <= Wgt_8_408;
		WeightsStore8[409] <= Wgt_8_409;
		WeightsStore8[410] <= Wgt_8_410;
		WeightsStore8[411] <= Wgt_8_411;
		WeightsStore8[412] <= Wgt_8_412;
		WeightsStore8[413] <= Wgt_8_413;
		WeightsStore8[414] <= Wgt_8_414;
		WeightsStore8[415] <= Wgt_8_415;
		WeightsStore8[416] <= Wgt_8_416;
		WeightsStore8[417] <= Wgt_8_417;
		WeightsStore8[418] <= Wgt_8_418;
		WeightsStore8[419] <= Wgt_8_419;
		WeightsStore8[420] <= Wgt_8_420;
		WeightsStore8[421] <= Wgt_8_421;
		WeightsStore8[422] <= Wgt_8_422;
		WeightsStore8[423] <= Wgt_8_423;
		WeightsStore8[424] <= Wgt_8_424;
		WeightsStore8[425] <= Wgt_8_425;
		WeightsStore8[426] <= Wgt_8_426;
		WeightsStore8[427] <= Wgt_8_427;
		WeightsStore8[428] <= Wgt_8_428;
		WeightsStore8[429] <= Wgt_8_429;
		WeightsStore8[430] <= Wgt_8_430;
		WeightsStore8[431] <= Wgt_8_431;
		WeightsStore8[432] <= Wgt_8_432;
		WeightsStore8[433] <= Wgt_8_433;
		WeightsStore8[434] <= Wgt_8_434;
		WeightsStore8[435] <= Wgt_8_435;
		WeightsStore8[436] <= Wgt_8_436;
		WeightsStore8[437] <= Wgt_8_437;
		WeightsStore8[438] <= Wgt_8_438;
		WeightsStore8[439] <= Wgt_8_439;
		WeightsStore8[440] <= Wgt_8_440;
		WeightsStore8[441] <= Wgt_8_441;
		WeightsStore8[442] <= Wgt_8_442;
		WeightsStore8[443] <= Wgt_8_443;
		WeightsStore8[444] <= Wgt_8_444;
		WeightsStore8[445] <= Wgt_8_445;
		WeightsStore8[446] <= Wgt_8_446;
		WeightsStore8[447] <= Wgt_8_447;
		WeightsStore8[448] <= Wgt_8_448;
		WeightsStore8[449] <= Wgt_8_449;
		WeightsStore8[450] <= Wgt_8_450;
		WeightsStore8[451] <= Wgt_8_451;
		WeightsStore8[452] <= Wgt_8_452;
		WeightsStore8[453] <= Wgt_8_453;
		WeightsStore8[454] <= Wgt_8_454;
		WeightsStore8[455] <= Wgt_8_455;
		WeightsStore8[456] <= Wgt_8_456;
		WeightsStore8[457] <= Wgt_8_457;
		WeightsStore8[458] <= Wgt_8_458;
		WeightsStore8[459] <= Wgt_8_459;
		WeightsStore8[460] <= Wgt_8_460;
		WeightsStore8[461] <= Wgt_8_461;
		WeightsStore8[462] <= Wgt_8_462;
		WeightsStore8[463] <= Wgt_8_463;
		WeightsStore8[464] <= Wgt_8_464;
		WeightsStore8[465] <= Wgt_8_465;
		WeightsStore8[466] <= Wgt_8_466;
		WeightsStore8[467] <= Wgt_8_467;
		WeightsStore8[468] <= Wgt_8_468;
		WeightsStore8[469] <= Wgt_8_469;
		WeightsStore8[470] <= Wgt_8_470;
		WeightsStore8[471] <= Wgt_8_471;
		WeightsStore8[472] <= Wgt_8_472;
		WeightsStore8[473] <= Wgt_8_473;
		WeightsStore8[474] <= Wgt_8_474;
		WeightsStore8[475] <= Wgt_8_475;
		WeightsStore8[476] <= Wgt_8_476;
		WeightsStore8[477] <= Wgt_8_477;
		WeightsStore8[478] <= Wgt_8_478;
		WeightsStore8[479] <= Wgt_8_479;
		WeightsStore8[480] <= Wgt_8_480;
		WeightsStore8[481] <= Wgt_8_481;
		WeightsStore8[482] <= Wgt_8_482;
		WeightsStore8[483] <= Wgt_8_483;
		WeightsStore8[484] <= Wgt_8_484;
		WeightsStore8[485] <= Wgt_8_485;
		WeightsStore8[486] <= Wgt_8_486;
		WeightsStore8[487] <= Wgt_8_487;
		WeightsStore8[488] <= Wgt_8_488;
		WeightsStore8[489] <= Wgt_8_489;
		WeightsStore8[490] <= Wgt_8_490;
		WeightsStore8[491] <= Wgt_8_491;
		WeightsStore8[492] <= Wgt_8_492;
		WeightsStore8[493] <= Wgt_8_493;
		WeightsStore8[494] <= Wgt_8_494;
		WeightsStore8[495] <= Wgt_8_495;
		WeightsStore8[496] <= Wgt_8_496;
		WeightsStore8[497] <= Wgt_8_497;
		WeightsStore8[498] <= Wgt_8_498;
		WeightsStore8[499] <= Wgt_8_499;
		WeightsStore8[500] <= Wgt_8_500;
		WeightsStore8[501] <= Wgt_8_501;
		WeightsStore8[502] <= Wgt_8_502;
		WeightsStore8[503] <= Wgt_8_503;
		WeightsStore8[504] <= Wgt_8_504;
		WeightsStore8[505] <= Wgt_8_505;
		WeightsStore8[506] <= Wgt_8_506;
		WeightsStore8[507] <= Wgt_8_507;
		WeightsStore8[508] <= Wgt_8_508;
		WeightsStore8[509] <= Wgt_8_509;
		WeightsStore8[510] <= Wgt_8_510;
		WeightsStore8[511] <= Wgt_8_511;
		WeightsStore8[512] <= Wgt_8_512;
		WeightsStore8[513] <= Wgt_8_513;
		WeightsStore8[514] <= Wgt_8_514;
		WeightsStore8[515] <= Wgt_8_515;
		WeightsStore8[516] <= Wgt_8_516;
		WeightsStore8[517] <= Wgt_8_517;
		WeightsStore8[518] <= Wgt_8_518;
		WeightsStore8[519] <= Wgt_8_519;
		WeightsStore8[520] <= Wgt_8_520;
		WeightsStore8[521] <= Wgt_8_521;
		WeightsStore8[522] <= Wgt_8_522;
		WeightsStore8[523] <= Wgt_8_523;
		WeightsStore8[524] <= Wgt_8_524;
		WeightsStore8[525] <= Wgt_8_525;
		WeightsStore8[526] <= Wgt_8_526;
		WeightsStore8[527] <= Wgt_8_527;
		WeightsStore8[528] <= Wgt_8_528;
		WeightsStore8[529] <= Wgt_8_529;
		WeightsStore8[530] <= Wgt_8_530;
		WeightsStore8[531] <= Wgt_8_531;
		WeightsStore8[532] <= Wgt_8_532;
		WeightsStore8[533] <= Wgt_8_533;
		WeightsStore8[534] <= Wgt_8_534;
		WeightsStore8[535] <= Wgt_8_535;
		WeightsStore8[536] <= Wgt_8_536;
		WeightsStore8[537] <= Wgt_8_537;
		WeightsStore8[538] <= Wgt_8_538;
		WeightsStore8[539] <= Wgt_8_539;
		WeightsStore8[540] <= Wgt_8_540;
		WeightsStore8[541] <= Wgt_8_541;
		WeightsStore8[542] <= Wgt_8_542;
		WeightsStore8[543] <= Wgt_8_543;
		WeightsStore8[544] <= Wgt_8_544;
		WeightsStore8[545] <= Wgt_8_545;
		WeightsStore8[546] <= Wgt_8_546;
		WeightsStore8[547] <= Wgt_8_547;
		WeightsStore8[548] <= Wgt_8_548;
		WeightsStore8[549] <= Wgt_8_549;
		WeightsStore8[550] <= Wgt_8_550;
		WeightsStore8[551] <= Wgt_8_551;
		WeightsStore8[552] <= Wgt_8_552;
		WeightsStore8[553] <= Wgt_8_553;
		WeightsStore8[554] <= Wgt_8_554;
		WeightsStore8[555] <= Wgt_8_555;
		WeightsStore8[556] <= Wgt_8_556;
		WeightsStore8[557] <= Wgt_8_557;
		WeightsStore8[558] <= Wgt_8_558;
		WeightsStore8[559] <= Wgt_8_559;
		WeightsStore8[560] <= Wgt_8_560;
		WeightsStore8[561] <= Wgt_8_561;
		WeightsStore8[562] <= Wgt_8_562;
		WeightsStore8[563] <= Wgt_8_563;
		WeightsStore8[564] <= Wgt_8_564;
		WeightsStore8[565] <= Wgt_8_565;
		WeightsStore8[566] <= Wgt_8_566;
		WeightsStore8[567] <= Wgt_8_567;
		WeightsStore8[568] <= Wgt_8_568;
		WeightsStore8[569] <= Wgt_8_569;
		WeightsStore8[570] <= Wgt_8_570;
		WeightsStore8[571] <= Wgt_8_571;
		WeightsStore8[572] <= Wgt_8_572;
		WeightsStore8[573] <= Wgt_8_573;
		WeightsStore8[574] <= Wgt_8_574;
		WeightsStore8[575] <= Wgt_8_575;
		WeightsStore8[576] <= Wgt_8_576;
		WeightsStore8[577] <= Wgt_8_577;
		WeightsStore8[578] <= Wgt_8_578;
		WeightsStore8[579] <= Wgt_8_579;
		WeightsStore8[580] <= Wgt_8_580;
		WeightsStore8[581] <= Wgt_8_581;
		WeightsStore8[582] <= Wgt_8_582;
		WeightsStore8[583] <= Wgt_8_583;
		WeightsStore8[584] <= Wgt_8_584;
		WeightsStore8[585] <= Wgt_8_585;
		WeightsStore8[586] <= Wgt_8_586;
		WeightsStore8[587] <= Wgt_8_587;
		WeightsStore8[588] <= Wgt_8_588;
		WeightsStore8[589] <= Wgt_8_589;
		WeightsStore8[590] <= Wgt_8_590;
		WeightsStore8[591] <= Wgt_8_591;
		WeightsStore8[592] <= Wgt_8_592;
		WeightsStore8[593] <= Wgt_8_593;
		WeightsStore8[594] <= Wgt_8_594;
		WeightsStore8[595] <= Wgt_8_595;
		WeightsStore8[596] <= Wgt_8_596;
		WeightsStore8[597] <= Wgt_8_597;
		WeightsStore8[598] <= Wgt_8_598;
		WeightsStore8[599] <= Wgt_8_599;
		WeightsStore8[600] <= Wgt_8_600;
		WeightsStore8[601] <= Wgt_8_601;
		WeightsStore8[602] <= Wgt_8_602;
		WeightsStore8[603] <= Wgt_8_603;
		WeightsStore8[604] <= Wgt_8_604;
		WeightsStore8[605] <= Wgt_8_605;
		WeightsStore8[606] <= Wgt_8_606;
		WeightsStore8[607] <= Wgt_8_607;
		WeightsStore8[608] <= Wgt_8_608;
		WeightsStore8[609] <= Wgt_8_609;
		WeightsStore8[610] <= Wgt_8_610;
		WeightsStore8[611] <= Wgt_8_611;
		WeightsStore8[612] <= Wgt_8_612;
		WeightsStore8[613] <= Wgt_8_613;
		WeightsStore8[614] <= Wgt_8_614;
		WeightsStore8[615] <= Wgt_8_615;
		WeightsStore8[616] <= Wgt_8_616;
		WeightsStore8[617] <= Wgt_8_617;
		WeightsStore8[618] <= Wgt_8_618;
		WeightsStore8[619] <= Wgt_8_619;
		WeightsStore8[620] <= Wgt_8_620;
		WeightsStore8[621] <= Wgt_8_621;
		WeightsStore8[622] <= Wgt_8_622;
		WeightsStore8[623] <= Wgt_8_623;
		WeightsStore8[624] <= Wgt_8_624;
		WeightsStore8[625] <= Wgt_8_625;
		WeightsStore8[626] <= Wgt_8_626;
		WeightsStore8[627] <= Wgt_8_627;
		WeightsStore8[628] <= Wgt_8_628;
		WeightsStore8[629] <= Wgt_8_629;
		WeightsStore8[630] <= Wgt_8_630;
		WeightsStore8[631] <= Wgt_8_631;
		WeightsStore8[632] <= Wgt_8_632;
		WeightsStore8[633] <= Wgt_8_633;
		WeightsStore8[634] <= Wgt_8_634;
		WeightsStore8[635] <= Wgt_8_635;
		WeightsStore8[636] <= Wgt_8_636;
		WeightsStore8[637] <= Wgt_8_637;
		WeightsStore8[638] <= Wgt_8_638;
		WeightsStore8[639] <= Wgt_8_639;
		WeightsStore8[640] <= Wgt_8_640;
		WeightsStore8[641] <= Wgt_8_641;
		WeightsStore8[642] <= Wgt_8_642;
		WeightsStore8[643] <= Wgt_8_643;
		WeightsStore8[644] <= Wgt_8_644;
		WeightsStore8[645] <= Wgt_8_645;
		WeightsStore8[646] <= Wgt_8_646;
		WeightsStore8[647] <= Wgt_8_647;
		WeightsStore8[648] <= Wgt_8_648;
		WeightsStore8[649] <= Wgt_8_649;
		WeightsStore8[650] <= Wgt_8_650;
		WeightsStore8[651] <= Wgt_8_651;
		WeightsStore8[652] <= Wgt_8_652;
		WeightsStore8[653] <= Wgt_8_653;
		WeightsStore8[654] <= Wgt_8_654;
		WeightsStore8[655] <= Wgt_8_655;
		WeightsStore8[656] <= Wgt_8_656;
		WeightsStore8[657] <= Wgt_8_657;
		WeightsStore8[658] <= Wgt_8_658;
		WeightsStore8[659] <= Wgt_8_659;
		WeightsStore8[660] <= Wgt_8_660;
		WeightsStore8[661] <= Wgt_8_661;
		WeightsStore8[662] <= Wgt_8_662;
		WeightsStore8[663] <= Wgt_8_663;
		WeightsStore8[664] <= Wgt_8_664;
		WeightsStore8[665] <= Wgt_8_665;
		WeightsStore8[666] <= Wgt_8_666;
		WeightsStore8[667] <= Wgt_8_667;
		WeightsStore8[668] <= Wgt_8_668;
		WeightsStore8[669] <= Wgt_8_669;
		WeightsStore8[670] <= Wgt_8_670;
		WeightsStore8[671] <= Wgt_8_671;
		WeightsStore8[672] <= Wgt_8_672;
		WeightsStore8[673] <= Wgt_8_673;
		WeightsStore8[674] <= Wgt_8_674;
		WeightsStore8[675] <= Wgt_8_675;
		WeightsStore8[676] <= Wgt_8_676;
		WeightsStore8[677] <= Wgt_8_677;
		WeightsStore8[678] <= Wgt_8_678;
		WeightsStore8[679] <= Wgt_8_679;
		WeightsStore8[680] <= Wgt_8_680;
		WeightsStore8[681] <= Wgt_8_681;
		WeightsStore8[682] <= Wgt_8_682;
		WeightsStore8[683] <= Wgt_8_683;
		WeightsStore8[684] <= Wgt_8_684;
		WeightsStore8[685] <= Wgt_8_685;
		WeightsStore8[686] <= Wgt_8_686;
		WeightsStore8[687] <= Wgt_8_687;
		WeightsStore8[688] <= Wgt_8_688;
		WeightsStore8[689] <= Wgt_8_689;
		WeightsStore8[690] <= Wgt_8_690;
		WeightsStore8[691] <= Wgt_8_691;
		WeightsStore8[692] <= Wgt_8_692;
		WeightsStore8[693] <= Wgt_8_693;
		WeightsStore8[694] <= Wgt_8_694;
		WeightsStore8[695] <= Wgt_8_695;
		WeightsStore8[696] <= Wgt_8_696;
		WeightsStore8[697] <= Wgt_8_697;
		WeightsStore8[698] <= Wgt_8_698;
		WeightsStore8[699] <= Wgt_8_699;
		WeightsStore8[700] <= Wgt_8_700;
		WeightsStore8[701] <= Wgt_8_701;
		WeightsStore8[702] <= Wgt_8_702;
		WeightsStore8[703] <= Wgt_8_703;
		WeightsStore8[704] <= Wgt_8_704;
		WeightsStore8[705] <= Wgt_8_705;
		WeightsStore8[706] <= Wgt_8_706;
		WeightsStore8[707] <= Wgt_8_707;
		WeightsStore8[708] <= Wgt_8_708;
		WeightsStore8[709] <= Wgt_8_709;
		WeightsStore8[710] <= Wgt_8_710;
		WeightsStore8[711] <= Wgt_8_711;
		WeightsStore8[712] <= Wgt_8_712;
		WeightsStore8[713] <= Wgt_8_713;
		WeightsStore8[714] <= Wgt_8_714;
		WeightsStore8[715] <= Wgt_8_715;
		WeightsStore8[716] <= Wgt_8_716;
		WeightsStore8[717] <= Wgt_8_717;
		WeightsStore8[718] <= Wgt_8_718;
		WeightsStore8[719] <= Wgt_8_719;
		WeightsStore8[720] <= Wgt_8_720;
		WeightsStore8[721] <= Wgt_8_721;
		WeightsStore8[722] <= Wgt_8_722;
		WeightsStore8[723] <= Wgt_8_723;
		WeightsStore8[724] <= Wgt_8_724;
		WeightsStore8[725] <= Wgt_8_725;
		WeightsStore8[726] <= Wgt_8_726;
		WeightsStore8[727] <= Wgt_8_727;
		WeightsStore8[728] <= Wgt_8_728;
		WeightsStore8[729] <= Wgt_8_729;
		WeightsStore8[730] <= Wgt_8_730;
		WeightsStore8[731] <= Wgt_8_731;
		WeightsStore8[732] <= Wgt_8_732;
		WeightsStore8[733] <= Wgt_8_733;
		WeightsStore8[734] <= Wgt_8_734;
		WeightsStore8[735] <= Wgt_8_735;
		WeightsStore8[736] <= Wgt_8_736;
		WeightsStore8[737] <= Wgt_8_737;
		WeightsStore8[738] <= Wgt_8_738;
		WeightsStore8[739] <= Wgt_8_739;
		WeightsStore8[740] <= Wgt_8_740;
		WeightsStore8[741] <= Wgt_8_741;
		WeightsStore8[742] <= Wgt_8_742;
		WeightsStore8[743] <= Wgt_8_743;
		WeightsStore8[744] <= Wgt_8_744;
		WeightsStore8[745] <= Wgt_8_745;
		WeightsStore8[746] <= Wgt_8_746;
		WeightsStore8[747] <= Wgt_8_747;
		WeightsStore8[748] <= Wgt_8_748;
		WeightsStore8[749] <= Wgt_8_749;
		WeightsStore8[750] <= Wgt_8_750;
		WeightsStore8[751] <= Wgt_8_751;
		WeightsStore8[752] <= Wgt_8_752;
		WeightsStore8[753] <= Wgt_8_753;
		WeightsStore8[754] <= Wgt_8_754;
		WeightsStore8[755] <= Wgt_8_755;
		WeightsStore8[756] <= Wgt_8_756;
		WeightsStore8[757] <= Wgt_8_757;
		WeightsStore8[758] <= Wgt_8_758;
		WeightsStore8[759] <= Wgt_8_759;
		WeightsStore8[760] <= Wgt_8_760;
		WeightsStore8[761] <= Wgt_8_761;
		WeightsStore8[762] <= Wgt_8_762;
		WeightsStore8[763] <= Wgt_8_763;
		WeightsStore8[764] <= Wgt_8_764;
		WeightsStore8[765] <= Wgt_8_765;
		WeightsStore8[766] <= Wgt_8_766;
		WeightsStore8[767] <= Wgt_8_767;
		WeightsStore8[768] <= Wgt_8_768;
		WeightsStore8[769] <= Wgt_8_769;
		WeightsStore8[770] <= Wgt_8_770;
		WeightsStore8[771] <= Wgt_8_771;
		WeightsStore8[772] <= Wgt_8_772;
		WeightsStore8[773] <= Wgt_8_773;
		WeightsStore8[774] <= Wgt_8_774;
		WeightsStore8[775] <= Wgt_8_775;
		WeightsStore8[776] <= Wgt_8_776;
		WeightsStore8[777] <= Wgt_8_777;
		WeightsStore8[778] <= Wgt_8_778;
		WeightsStore8[779] <= Wgt_8_779;
		WeightsStore8[780] <= Wgt_8_780;
		WeightsStore8[781] <= Wgt_8_781;
		WeightsStore8[782] <= Wgt_8_782;
		WeightsStore8[783] <= Wgt_8_783;
		WeightsStore8[784] <= Wgt_8_784;
		WeightsStore9[0] <= Wgt_9_0;
		WeightsStore9[1] <= Wgt_9_1;
		WeightsStore9[2] <= Wgt_9_2;
		WeightsStore9[3] <= Wgt_9_3;
		WeightsStore9[4] <= Wgt_9_4;
		WeightsStore9[5] <= Wgt_9_5;
		WeightsStore9[6] <= Wgt_9_6;
		WeightsStore9[7] <= Wgt_9_7;
		WeightsStore9[8] <= Wgt_9_8;
		WeightsStore9[9] <= Wgt_9_9;
		WeightsStore9[10] <= Wgt_9_10;
		WeightsStore9[11] <= Wgt_9_11;
		WeightsStore9[12] <= Wgt_9_12;
		WeightsStore9[13] <= Wgt_9_13;
		WeightsStore9[14] <= Wgt_9_14;
		WeightsStore9[15] <= Wgt_9_15;
		WeightsStore9[16] <= Wgt_9_16;
		WeightsStore9[17] <= Wgt_9_17;
		WeightsStore9[18] <= Wgt_9_18;
		WeightsStore9[19] <= Wgt_9_19;
		WeightsStore9[20] <= Wgt_9_20;
		WeightsStore9[21] <= Wgt_9_21;
		WeightsStore9[22] <= Wgt_9_22;
		WeightsStore9[23] <= Wgt_9_23;
		WeightsStore9[24] <= Wgt_9_24;
		WeightsStore9[25] <= Wgt_9_25;
		WeightsStore9[26] <= Wgt_9_26;
		WeightsStore9[27] <= Wgt_9_27;
		WeightsStore9[28] <= Wgt_9_28;
		WeightsStore9[29] <= Wgt_9_29;
		WeightsStore9[30] <= Wgt_9_30;
		WeightsStore9[31] <= Wgt_9_31;
		WeightsStore9[32] <= Wgt_9_32;
		WeightsStore9[33] <= Wgt_9_33;
		WeightsStore9[34] <= Wgt_9_34;
		WeightsStore9[35] <= Wgt_9_35;
		WeightsStore9[36] <= Wgt_9_36;
		WeightsStore9[37] <= Wgt_9_37;
		WeightsStore9[38] <= Wgt_9_38;
		WeightsStore9[39] <= Wgt_9_39;
		WeightsStore9[40] <= Wgt_9_40;
		WeightsStore9[41] <= Wgt_9_41;
		WeightsStore9[42] <= Wgt_9_42;
		WeightsStore9[43] <= Wgt_9_43;
		WeightsStore9[44] <= Wgt_9_44;
		WeightsStore9[45] <= Wgt_9_45;
		WeightsStore9[46] <= Wgt_9_46;
		WeightsStore9[47] <= Wgt_9_47;
		WeightsStore9[48] <= Wgt_9_48;
		WeightsStore9[49] <= Wgt_9_49;
		WeightsStore9[50] <= Wgt_9_50;
		WeightsStore9[51] <= Wgt_9_51;
		WeightsStore9[52] <= Wgt_9_52;
		WeightsStore9[53] <= Wgt_9_53;
		WeightsStore9[54] <= Wgt_9_54;
		WeightsStore9[55] <= Wgt_9_55;
		WeightsStore9[56] <= Wgt_9_56;
		WeightsStore9[57] <= Wgt_9_57;
		WeightsStore9[58] <= Wgt_9_58;
		WeightsStore9[59] <= Wgt_9_59;
		WeightsStore9[60] <= Wgt_9_60;
		WeightsStore9[61] <= Wgt_9_61;
		WeightsStore9[62] <= Wgt_9_62;
		WeightsStore9[63] <= Wgt_9_63;
		WeightsStore9[64] <= Wgt_9_64;
		WeightsStore9[65] <= Wgt_9_65;
		WeightsStore9[66] <= Wgt_9_66;
		WeightsStore9[67] <= Wgt_9_67;
		WeightsStore9[68] <= Wgt_9_68;
		WeightsStore9[69] <= Wgt_9_69;
		WeightsStore9[70] <= Wgt_9_70;
		WeightsStore9[71] <= Wgt_9_71;
		WeightsStore9[72] <= Wgt_9_72;
		WeightsStore9[73] <= Wgt_9_73;
		WeightsStore9[74] <= Wgt_9_74;
		WeightsStore9[75] <= Wgt_9_75;
		WeightsStore9[76] <= Wgt_9_76;
		WeightsStore9[77] <= Wgt_9_77;
		WeightsStore9[78] <= Wgt_9_78;
		WeightsStore9[79] <= Wgt_9_79;
		WeightsStore9[80] <= Wgt_9_80;
		WeightsStore9[81] <= Wgt_9_81;
		WeightsStore9[82] <= Wgt_9_82;
		WeightsStore9[83] <= Wgt_9_83;
		WeightsStore9[84] <= Wgt_9_84;
		WeightsStore9[85] <= Wgt_9_85;
		WeightsStore9[86] <= Wgt_9_86;
		WeightsStore9[87] <= Wgt_9_87;
		WeightsStore9[88] <= Wgt_9_88;
		WeightsStore9[89] <= Wgt_9_89;
		WeightsStore9[90] <= Wgt_9_90;
		WeightsStore9[91] <= Wgt_9_91;
		WeightsStore9[92] <= Wgt_9_92;
		WeightsStore9[93] <= Wgt_9_93;
		WeightsStore9[94] <= Wgt_9_94;
		WeightsStore9[95] <= Wgt_9_95;
		WeightsStore9[96] <= Wgt_9_96;
		WeightsStore9[97] <= Wgt_9_97;
		WeightsStore9[98] <= Wgt_9_98;
		WeightsStore9[99] <= Wgt_9_99;
		WeightsStore9[100] <= Wgt_9_100;
		WeightsStore9[101] <= Wgt_9_101;
		WeightsStore9[102] <= Wgt_9_102;
		WeightsStore9[103] <= Wgt_9_103;
		WeightsStore9[104] <= Wgt_9_104;
		WeightsStore9[105] <= Wgt_9_105;
		WeightsStore9[106] <= Wgt_9_106;
		WeightsStore9[107] <= Wgt_9_107;
		WeightsStore9[108] <= Wgt_9_108;
		WeightsStore9[109] <= Wgt_9_109;
		WeightsStore9[110] <= Wgt_9_110;
		WeightsStore9[111] <= Wgt_9_111;
		WeightsStore9[112] <= Wgt_9_112;
		WeightsStore9[113] <= Wgt_9_113;
		WeightsStore9[114] <= Wgt_9_114;
		WeightsStore9[115] <= Wgt_9_115;
		WeightsStore9[116] <= Wgt_9_116;
		WeightsStore9[117] <= Wgt_9_117;
		WeightsStore9[118] <= Wgt_9_118;
		WeightsStore9[119] <= Wgt_9_119;
		WeightsStore9[120] <= Wgt_9_120;
		WeightsStore9[121] <= Wgt_9_121;
		WeightsStore9[122] <= Wgt_9_122;
		WeightsStore9[123] <= Wgt_9_123;
		WeightsStore9[124] <= Wgt_9_124;
		WeightsStore9[125] <= Wgt_9_125;
		WeightsStore9[126] <= Wgt_9_126;
		WeightsStore9[127] <= Wgt_9_127;
		WeightsStore9[128] <= Wgt_9_128;
		WeightsStore9[129] <= Wgt_9_129;
		WeightsStore9[130] <= Wgt_9_130;
		WeightsStore9[131] <= Wgt_9_131;
		WeightsStore9[132] <= Wgt_9_132;
		WeightsStore9[133] <= Wgt_9_133;
		WeightsStore9[134] <= Wgt_9_134;
		WeightsStore9[135] <= Wgt_9_135;
		WeightsStore9[136] <= Wgt_9_136;
		WeightsStore9[137] <= Wgt_9_137;
		WeightsStore9[138] <= Wgt_9_138;
		WeightsStore9[139] <= Wgt_9_139;
		WeightsStore9[140] <= Wgt_9_140;
		WeightsStore9[141] <= Wgt_9_141;
		WeightsStore9[142] <= Wgt_9_142;
		WeightsStore9[143] <= Wgt_9_143;
		WeightsStore9[144] <= Wgt_9_144;
		WeightsStore9[145] <= Wgt_9_145;
		WeightsStore9[146] <= Wgt_9_146;
		WeightsStore9[147] <= Wgt_9_147;
		WeightsStore9[148] <= Wgt_9_148;
		WeightsStore9[149] <= Wgt_9_149;
		WeightsStore9[150] <= Wgt_9_150;
		WeightsStore9[151] <= Wgt_9_151;
		WeightsStore9[152] <= Wgt_9_152;
		WeightsStore9[153] <= Wgt_9_153;
		WeightsStore9[154] <= Wgt_9_154;
		WeightsStore9[155] <= Wgt_9_155;
		WeightsStore9[156] <= Wgt_9_156;
		WeightsStore9[157] <= Wgt_9_157;
		WeightsStore9[158] <= Wgt_9_158;
		WeightsStore9[159] <= Wgt_9_159;
		WeightsStore9[160] <= Wgt_9_160;
		WeightsStore9[161] <= Wgt_9_161;
		WeightsStore9[162] <= Wgt_9_162;
		WeightsStore9[163] <= Wgt_9_163;
		WeightsStore9[164] <= Wgt_9_164;
		WeightsStore9[165] <= Wgt_9_165;
		WeightsStore9[166] <= Wgt_9_166;
		WeightsStore9[167] <= Wgt_9_167;
		WeightsStore9[168] <= Wgt_9_168;
		WeightsStore9[169] <= Wgt_9_169;
		WeightsStore9[170] <= Wgt_9_170;
		WeightsStore9[171] <= Wgt_9_171;
		WeightsStore9[172] <= Wgt_9_172;
		WeightsStore9[173] <= Wgt_9_173;
		WeightsStore9[174] <= Wgt_9_174;
		WeightsStore9[175] <= Wgt_9_175;
		WeightsStore9[176] <= Wgt_9_176;
		WeightsStore9[177] <= Wgt_9_177;
		WeightsStore9[178] <= Wgt_9_178;
		WeightsStore9[179] <= Wgt_9_179;
		WeightsStore9[180] <= Wgt_9_180;
		WeightsStore9[181] <= Wgt_9_181;
		WeightsStore9[182] <= Wgt_9_182;
		WeightsStore9[183] <= Wgt_9_183;
		WeightsStore9[184] <= Wgt_9_184;
		WeightsStore9[185] <= Wgt_9_185;
		WeightsStore9[186] <= Wgt_9_186;
		WeightsStore9[187] <= Wgt_9_187;
		WeightsStore9[188] <= Wgt_9_188;
		WeightsStore9[189] <= Wgt_9_189;
		WeightsStore9[190] <= Wgt_9_190;
		WeightsStore9[191] <= Wgt_9_191;
		WeightsStore9[192] <= Wgt_9_192;
		WeightsStore9[193] <= Wgt_9_193;
		WeightsStore9[194] <= Wgt_9_194;
		WeightsStore9[195] <= Wgt_9_195;
		WeightsStore9[196] <= Wgt_9_196;
		WeightsStore9[197] <= Wgt_9_197;
		WeightsStore9[198] <= Wgt_9_198;
		WeightsStore9[199] <= Wgt_9_199;
		WeightsStore9[200] <= Wgt_9_200;
		WeightsStore9[201] <= Wgt_9_201;
		WeightsStore9[202] <= Wgt_9_202;
		WeightsStore9[203] <= Wgt_9_203;
		WeightsStore9[204] <= Wgt_9_204;
		WeightsStore9[205] <= Wgt_9_205;
		WeightsStore9[206] <= Wgt_9_206;
		WeightsStore9[207] <= Wgt_9_207;
		WeightsStore9[208] <= Wgt_9_208;
		WeightsStore9[209] <= Wgt_9_209;
		WeightsStore9[210] <= Wgt_9_210;
		WeightsStore9[211] <= Wgt_9_211;
		WeightsStore9[212] <= Wgt_9_212;
		WeightsStore9[213] <= Wgt_9_213;
		WeightsStore9[214] <= Wgt_9_214;
		WeightsStore9[215] <= Wgt_9_215;
		WeightsStore9[216] <= Wgt_9_216;
		WeightsStore9[217] <= Wgt_9_217;
		WeightsStore9[218] <= Wgt_9_218;
		WeightsStore9[219] <= Wgt_9_219;
		WeightsStore9[220] <= Wgt_9_220;
		WeightsStore9[221] <= Wgt_9_221;
		WeightsStore9[222] <= Wgt_9_222;
		WeightsStore9[223] <= Wgt_9_223;
		WeightsStore9[224] <= Wgt_9_224;
		WeightsStore9[225] <= Wgt_9_225;
		WeightsStore9[226] <= Wgt_9_226;
		WeightsStore9[227] <= Wgt_9_227;
		WeightsStore9[228] <= Wgt_9_228;
		WeightsStore9[229] <= Wgt_9_229;
		WeightsStore9[230] <= Wgt_9_230;
		WeightsStore9[231] <= Wgt_9_231;
		WeightsStore9[232] <= Wgt_9_232;
		WeightsStore9[233] <= Wgt_9_233;
		WeightsStore9[234] <= Wgt_9_234;
		WeightsStore9[235] <= Wgt_9_235;
		WeightsStore9[236] <= Wgt_9_236;
		WeightsStore9[237] <= Wgt_9_237;
		WeightsStore9[238] <= Wgt_9_238;
		WeightsStore9[239] <= Wgt_9_239;
		WeightsStore9[240] <= Wgt_9_240;
		WeightsStore9[241] <= Wgt_9_241;
		WeightsStore9[242] <= Wgt_9_242;
		WeightsStore9[243] <= Wgt_9_243;
		WeightsStore9[244] <= Wgt_9_244;
		WeightsStore9[245] <= Wgt_9_245;
		WeightsStore9[246] <= Wgt_9_246;
		WeightsStore9[247] <= Wgt_9_247;
		WeightsStore9[248] <= Wgt_9_248;
		WeightsStore9[249] <= Wgt_9_249;
		WeightsStore9[250] <= Wgt_9_250;
		WeightsStore9[251] <= Wgt_9_251;
		WeightsStore9[252] <= Wgt_9_252;
		WeightsStore9[253] <= Wgt_9_253;
		WeightsStore9[254] <= Wgt_9_254;
		WeightsStore9[255] <= Wgt_9_255;
		WeightsStore9[256] <= Wgt_9_256;
		WeightsStore9[257] <= Wgt_9_257;
		WeightsStore9[258] <= Wgt_9_258;
		WeightsStore9[259] <= Wgt_9_259;
		WeightsStore9[260] <= Wgt_9_260;
		WeightsStore9[261] <= Wgt_9_261;
		WeightsStore9[262] <= Wgt_9_262;
		WeightsStore9[263] <= Wgt_9_263;
		WeightsStore9[264] <= Wgt_9_264;
		WeightsStore9[265] <= Wgt_9_265;
		WeightsStore9[266] <= Wgt_9_266;
		WeightsStore9[267] <= Wgt_9_267;
		WeightsStore9[268] <= Wgt_9_268;
		WeightsStore9[269] <= Wgt_9_269;
		WeightsStore9[270] <= Wgt_9_270;
		WeightsStore9[271] <= Wgt_9_271;
		WeightsStore9[272] <= Wgt_9_272;
		WeightsStore9[273] <= Wgt_9_273;
		WeightsStore9[274] <= Wgt_9_274;
		WeightsStore9[275] <= Wgt_9_275;
		WeightsStore9[276] <= Wgt_9_276;
		WeightsStore9[277] <= Wgt_9_277;
		WeightsStore9[278] <= Wgt_9_278;
		WeightsStore9[279] <= Wgt_9_279;
		WeightsStore9[280] <= Wgt_9_280;
		WeightsStore9[281] <= Wgt_9_281;
		WeightsStore9[282] <= Wgt_9_282;
		WeightsStore9[283] <= Wgt_9_283;
		WeightsStore9[284] <= Wgt_9_284;
		WeightsStore9[285] <= Wgt_9_285;
		WeightsStore9[286] <= Wgt_9_286;
		WeightsStore9[287] <= Wgt_9_287;
		WeightsStore9[288] <= Wgt_9_288;
		WeightsStore9[289] <= Wgt_9_289;
		WeightsStore9[290] <= Wgt_9_290;
		WeightsStore9[291] <= Wgt_9_291;
		WeightsStore9[292] <= Wgt_9_292;
		WeightsStore9[293] <= Wgt_9_293;
		WeightsStore9[294] <= Wgt_9_294;
		WeightsStore9[295] <= Wgt_9_295;
		WeightsStore9[296] <= Wgt_9_296;
		WeightsStore9[297] <= Wgt_9_297;
		WeightsStore9[298] <= Wgt_9_298;
		WeightsStore9[299] <= Wgt_9_299;
		WeightsStore9[300] <= Wgt_9_300;
		WeightsStore9[301] <= Wgt_9_301;
		WeightsStore9[302] <= Wgt_9_302;
		WeightsStore9[303] <= Wgt_9_303;
		WeightsStore9[304] <= Wgt_9_304;
		WeightsStore9[305] <= Wgt_9_305;
		WeightsStore9[306] <= Wgt_9_306;
		WeightsStore9[307] <= Wgt_9_307;
		WeightsStore9[308] <= Wgt_9_308;
		WeightsStore9[309] <= Wgt_9_309;
		WeightsStore9[310] <= Wgt_9_310;
		WeightsStore9[311] <= Wgt_9_311;
		WeightsStore9[312] <= Wgt_9_312;
		WeightsStore9[313] <= Wgt_9_313;
		WeightsStore9[314] <= Wgt_9_314;
		WeightsStore9[315] <= Wgt_9_315;
		WeightsStore9[316] <= Wgt_9_316;
		WeightsStore9[317] <= Wgt_9_317;
		WeightsStore9[318] <= Wgt_9_318;
		WeightsStore9[319] <= Wgt_9_319;
		WeightsStore9[320] <= Wgt_9_320;
		WeightsStore9[321] <= Wgt_9_321;
		WeightsStore9[322] <= Wgt_9_322;
		WeightsStore9[323] <= Wgt_9_323;
		WeightsStore9[324] <= Wgt_9_324;
		WeightsStore9[325] <= Wgt_9_325;
		WeightsStore9[326] <= Wgt_9_326;
		WeightsStore9[327] <= Wgt_9_327;
		WeightsStore9[328] <= Wgt_9_328;
		WeightsStore9[329] <= Wgt_9_329;
		WeightsStore9[330] <= Wgt_9_330;
		WeightsStore9[331] <= Wgt_9_331;
		WeightsStore9[332] <= Wgt_9_332;
		WeightsStore9[333] <= Wgt_9_333;
		WeightsStore9[334] <= Wgt_9_334;
		WeightsStore9[335] <= Wgt_9_335;
		WeightsStore9[336] <= Wgt_9_336;
		WeightsStore9[337] <= Wgt_9_337;
		WeightsStore9[338] <= Wgt_9_338;
		WeightsStore9[339] <= Wgt_9_339;
		WeightsStore9[340] <= Wgt_9_340;
		WeightsStore9[341] <= Wgt_9_341;
		WeightsStore9[342] <= Wgt_9_342;
		WeightsStore9[343] <= Wgt_9_343;
		WeightsStore9[344] <= Wgt_9_344;
		WeightsStore9[345] <= Wgt_9_345;
		WeightsStore9[346] <= Wgt_9_346;
		WeightsStore9[347] <= Wgt_9_347;
		WeightsStore9[348] <= Wgt_9_348;
		WeightsStore9[349] <= Wgt_9_349;
		WeightsStore9[350] <= Wgt_9_350;
		WeightsStore9[351] <= Wgt_9_351;
		WeightsStore9[352] <= Wgt_9_352;
		WeightsStore9[353] <= Wgt_9_353;
		WeightsStore9[354] <= Wgt_9_354;
		WeightsStore9[355] <= Wgt_9_355;
		WeightsStore9[356] <= Wgt_9_356;
		WeightsStore9[357] <= Wgt_9_357;
		WeightsStore9[358] <= Wgt_9_358;
		WeightsStore9[359] <= Wgt_9_359;
		WeightsStore9[360] <= Wgt_9_360;
		WeightsStore9[361] <= Wgt_9_361;
		WeightsStore9[362] <= Wgt_9_362;
		WeightsStore9[363] <= Wgt_9_363;
		WeightsStore9[364] <= Wgt_9_364;
		WeightsStore9[365] <= Wgt_9_365;
		WeightsStore9[366] <= Wgt_9_366;
		WeightsStore9[367] <= Wgt_9_367;
		WeightsStore9[368] <= Wgt_9_368;
		WeightsStore9[369] <= Wgt_9_369;
		WeightsStore9[370] <= Wgt_9_370;
		WeightsStore9[371] <= Wgt_9_371;
		WeightsStore9[372] <= Wgt_9_372;
		WeightsStore9[373] <= Wgt_9_373;
		WeightsStore9[374] <= Wgt_9_374;
		WeightsStore9[375] <= Wgt_9_375;
		WeightsStore9[376] <= Wgt_9_376;
		WeightsStore9[377] <= Wgt_9_377;
		WeightsStore9[378] <= Wgt_9_378;
		WeightsStore9[379] <= Wgt_9_379;
		WeightsStore9[380] <= Wgt_9_380;
		WeightsStore9[381] <= Wgt_9_381;
		WeightsStore9[382] <= Wgt_9_382;
		WeightsStore9[383] <= Wgt_9_383;
		WeightsStore9[384] <= Wgt_9_384;
		WeightsStore9[385] <= Wgt_9_385;
		WeightsStore9[386] <= Wgt_9_386;
		WeightsStore9[387] <= Wgt_9_387;
		WeightsStore9[388] <= Wgt_9_388;
		WeightsStore9[389] <= Wgt_9_389;
		WeightsStore9[390] <= Wgt_9_390;
		WeightsStore9[391] <= Wgt_9_391;
		WeightsStore9[392] <= Wgt_9_392;
		WeightsStore9[393] <= Wgt_9_393;
		WeightsStore9[394] <= Wgt_9_394;
		WeightsStore9[395] <= Wgt_9_395;
		WeightsStore9[396] <= Wgt_9_396;
		WeightsStore9[397] <= Wgt_9_397;
		WeightsStore9[398] <= Wgt_9_398;
		WeightsStore9[399] <= Wgt_9_399;
		WeightsStore9[400] <= Wgt_9_400;
		WeightsStore9[401] <= Wgt_9_401;
		WeightsStore9[402] <= Wgt_9_402;
		WeightsStore9[403] <= Wgt_9_403;
		WeightsStore9[404] <= Wgt_9_404;
		WeightsStore9[405] <= Wgt_9_405;
		WeightsStore9[406] <= Wgt_9_406;
		WeightsStore9[407] <= Wgt_9_407;
		WeightsStore9[408] <= Wgt_9_408;
		WeightsStore9[409] <= Wgt_9_409;
		WeightsStore9[410] <= Wgt_9_410;
		WeightsStore9[411] <= Wgt_9_411;
		WeightsStore9[412] <= Wgt_9_412;
		WeightsStore9[413] <= Wgt_9_413;
		WeightsStore9[414] <= Wgt_9_414;
		WeightsStore9[415] <= Wgt_9_415;
		WeightsStore9[416] <= Wgt_9_416;
		WeightsStore9[417] <= Wgt_9_417;
		WeightsStore9[418] <= Wgt_9_418;
		WeightsStore9[419] <= Wgt_9_419;
		WeightsStore9[420] <= Wgt_9_420;
		WeightsStore9[421] <= Wgt_9_421;
		WeightsStore9[422] <= Wgt_9_422;
		WeightsStore9[423] <= Wgt_9_423;
		WeightsStore9[424] <= Wgt_9_424;
		WeightsStore9[425] <= Wgt_9_425;
		WeightsStore9[426] <= Wgt_9_426;
		WeightsStore9[427] <= Wgt_9_427;
		WeightsStore9[428] <= Wgt_9_428;
		WeightsStore9[429] <= Wgt_9_429;
		WeightsStore9[430] <= Wgt_9_430;
		WeightsStore9[431] <= Wgt_9_431;
		WeightsStore9[432] <= Wgt_9_432;
		WeightsStore9[433] <= Wgt_9_433;
		WeightsStore9[434] <= Wgt_9_434;
		WeightsStore9[435] <= Wgt_9_435;
		WeightsStore9[436] <= Wgt_9_436;
		WeightsStore9[437] <= Wgt_9_437;
		WeightsStore9[438] <= Wgt_9_438;
		WeightsStore9[439] <= Wgt_9_439;
		WeightsStore9[440] <= Wgt_9_440;
		WeightsStore9[441] <= Wgt_9_441;
		WeightsStore9[442] <= Wgt_9_442;
		WeightsStore9[443] <= Wgt_9_443;
		WeightsStore9[444] <= Wgt_9_444;
		WeightsStore9[445] <= Wgt_9_445;
		WeightsStore9[446] <= Wgt_9_446;
		WeightsStore9[447] <= Wgt_9_447;
		WeightsStore9[448] <= Wgt_9_448;
		WeightsStore9[449] <= Wgt_9_449;
		WeightsStore9[450] <= Wgt_9_450;
		WeightsStore9[451] <= Wgt_9_451;
		WeightsStore9[452] <= Wgt_9_452;
		WeightsStore9[453] <= Wgt_9_453;
		WeightsStore9[454] <= Wgt_9_454;
		WeightsStore9[455] <= Wgt_9_455;
		WeightsStore9[456] <= Wgt_9_456;
		WeightsStore9[457] <= Wgt_9_457;
		WeightsStore9[458] <= Wgt_9_458;
		WeightsStore9[459] <= Wgt_9_459;
		WeightsStore9[460] <= Wgt_9_460;
		WeightsStore9[461] <= Wgt_9_461;
		WeightsStore9[462] <= Wgt_9_462;
		WeightsStore9[463] <= Wgt_9_463;
		WeightsStore9[464] <= Wgt_9_464;
		WeightsStore9[465] <= Wgt_9_465;
		WeightsStore9[466] <= Wgt_9_466;
		WeightsStore9[467] <= Wgt_9_467;
		WeightsStore9[468] <= Wgt_9_468;
		WeightsStore9[469] <= Wgt_9_469;
		WeightsStore9[470] <= Wgt_9_470;
		WeightsStore9[471] <= Wgt_9_471;
		WeightsStore9[472] <= Wgt_9_472;
		WeightsStore9[473] <= Wgt_9_473;
		WeightsStore9[474] <= Wgt_9_474;
		WeightsStore9[475] <= Wgt_9_475;
		WeightsStore9[476] <= Wgt_9_476;
		WeightsStore9[477] <= Wgt_9_477;
		WeightsStore9[478] <= Wgt_9_478;
		WeightsStore9[479] <= Wgt_9_479;
		WeightsStore9[480] <= Wgt_9_480;
		WeightsStore9[481] <= Wgt_9_481;
		WeightsStore9[482] <= Wgt_9_482;
		WeightsStore9[483] <= Wgt_9_483;
		WeightsStore9[484] <= Wgt_9_484;
		WeightsStore9[485] <= Wgt_9_485;
		WeightsStore9[486] <= Wgt_9_486;
		WeightsStore9[487] <= Wgt_9_487;
		WeightsStore9[488] <= Wgt_9_488;
		WeightsStore9[489] <= Wgt_9_489;
		WeightsStore9[490] <= Wgt_9_490;
		WeightsStore9[491] <= Wgt_9_491;
		WeightsStore9[492] <= Wgt_9_492;
		WeightsStore9[493] <= Wgt_9_493;
		WeightsStore9[494] <= Wgt_9_494;
		WeightsStore9[495] <= Wgt_9_495;
		WeightsStore9[496] <= Wgt_9_496;
		WeightsStore9[497] <= Wgt_9_497;
		WeightsStore9[498] <= Wgt_9_498;
		WeightsStore9[499] <= Wgt_9_499;
		WeightsStore9[500] <= Wgt_9_500;
		WeightsStore9[501] <= Wgt_9_501;
		WeightsStore9[502] <= Wgt_9_502;
		WeightsStore9[503] <= Wgt_9_503;
		WeightsStore9[504] <= Wgt_9_504;
		WeightsStore9[505] <= Wgt_9_505;
		WeightsStore9[506] <= Wgt_9_506;
		WeightsStore9[507] <= Wgt_9_507;
		WeightsStore9[508] <= Wgt_9_508;
		WeightsStore9[509] <= Wgt_9_509;
		WeightsStore9[510] <= Wgt_9_510;
		WeightsStore9[511] <= Wgt_9_511;
		WeightsStore9[512] <= Wgt_9_512;
		WeightsStore9[513] <= Wgt_9_513;
		WeightsStore9[514] <= Wgt_9_514;
		WeightsStore9[515] <= Wgt_9_515;
		WeightsStore9[516] <= Wgt_9_516;
		WeightsStore9[517] <= Wgt_9_517;
		WeightsStore9[518] <= Wgt_9_518;
		WeightsStore9[519] <= Wgt_9_519;
		WeightsStore9[520] <= Wgt_9_520;
		WeightsStore9[521] <= Wgt_9_521;
		WeightsStore9[522] <= Wgt_9_522;
		WeightsStore9[523] <= Wgt_9_523;
		WeightsStore9[524] <= Wgt_9_524;
		WeightsStore9[525] <= Wgt_9_525;
		WeightsStore9[526] <= Wgt_9_526;
		WeightsStore9[527] <= Wgt_9_527;
		WeightsStore9[528] <= Wgt_9_528;
		WeightsStore9[529] <= Wgt_9_529;
		WeightsStore9[530] <= Wgt_9_530;
		WeightsStore9[531] <= Wgt_9_531;
		WeightsStore9[532] <= Wgt_9_532;
		WeightsStore9[533] <= Wgt_9_533;
		WeightsStore9[534] <= Wgt_9_534;
		WeightsStore9[535] <= Wgt_9_535;
		WeightsStore9[536] <= Wgt_9_536;
		WeightsStore9[537] <= Wgt_9_537;
		WeightsStore9[538] <= Wgt_9_538;
		WeightsStore9[539] <= Wgt_9_539;
		WeightsStore9[540] <= Wgt_9_540;
		WeightsStore9[541] <= Wgt_9_541;
		WeightsStore9[542] <= Wgt_9_542;
		WeightsStore9[543] <= Wgt_9_543;
		WeightsStore9[544] <= Wgt_9_544;
		WeightsStore9[545] <= Wgt_9_545;
		WeightsStore9[546] <= Wgt_9_546;
		WeightsStore9[547] <= Wgt_9_547;
		WeightsStore9[548] <= Wgt_9_548;
		WeightsStore9[549] <= Wgt_9_549;
		WeightsStore9[550] <= Wgt_9_550;
		WeightsStore9[551] <= Wgt_9_551;
		WeightsStore9[552] <= Wgt_9_552;
		WeightsStore9[553] <= Wgt_9_553;
		WeightsStore9[554] <= Wgt_9_554;
		WeightsStore9[555] <= Wgt_9_555;
		WeightsStore9[556] <= Wgt_9_556;
		WeightsStore9[557] <= Wgt_9_557;
		WeightsStore9[558] <= Wgt_9_558;
		WeightsStore9[559] <= Wgt_9_559;
		WeightsStore9[560] <= Wgt_9_560;
		WeightsStore9[561] <= Wgt_9_561;
		WeightsStore9[562] <= Wgt_9_562;
		WeightsStore9[563] <= Wgt_9_563;
		WeightsStore9[564] <= Wgt_9_564;
		WeightsStore9[565] <= Wgt_9_565;
		WeightsStore9[566] <= Wgt_9_566;
		WeightsStore9[567] <= Wgt_9_567;
		WeightsStore9[568] <= Wgt_9_568;
		WeightsStore9[569] <= Wgt_9_569;
		WeightsStore9[570] <= Wgt_9_570;
		WeightsStore9[571] <= Wgt_9_571;
		WeightsStore9[572] <= Wgt_9_572;
		WeightsStore9[573] <= Wgt_9_573;
		WeightsStore9[574] <= Wgt_9_574;
		WeightsStore9[575] <= Wgt_9_575;
		WeightsStore9[576] <= Wgt_9_576;
		WeightsStore9[577] <= Wgt_9_577;
		WeightsStore9[578] <= Wgt_9_578;
		WeightsStore9[579] <= Wgt_9_579;
		WeightsStore9[580] <= Wgt_9_580;
		WeightsStore9[581] <= Wgt_9_581;
		WeightsStore9[582] <= Wgt_9_582;
		WeightsStore9[583] <= Wgt_9_583;
		WeightsStore9[584] <= Wgt_9_584;
		WeightsStore9[585] <= Wgt_9_585;
		WeightsStore9[586] <= Wgt_9_586;
		WeightsStore9[587] <= Wgt_9_587;
		WeightsStore9[588] <= Wgt_9_588;
		WeightsStore9[589] <= Wgt_9_589;
		WeightsStore9[590] <= Wgt_9_590;
		WeightsStore9[591] <= Wgt_9_591;
		WeightsStore9[592] <= Wgt_9_592;
		WeightsStore9[593] <= Wgt_9_593;
		WeightsStore9[594] <= Wgt_9_594;
		WeightsStore9[595] <= Wgt_9_595;
		WeightsStore9[596] <= Wgt_9_596;
		WeightsStore9[597] <= Wgt_9_597;
		WeightsStore9[598] <= Wgt_9_598;
		WeightsStore9[599] <= Wgt_9_599;
		WeightsStore9[600] <= Wgt_9_600;
		WeightsStore9[601] <= Wgt_9_601;
		WeightsStore9[602] <= Wgt_9_602;
		WeightsStore9[603] <= Wgt_9_603;
		WeightsStore9[604] <= Wgt_9_604;
		WeightsStore9[605] <= Wgt_9_605;
		WeightsStore9[606] <= Wgt_9_606;
		WeightsStore9[607] <= Wgt_9_607;
		WeightsStore9[608] <= Wgt_9_608;
		WeightsStore9[609] <= Wgt_9_609;
		WeightsStore9[610] <= Wgt_9_610;
		WeightsStore9[611] <= Wgt_9_611;
		WeightsStore9[612] <= Wgt_9_612;
		WeightsStore9[613] <= Wgt_9_613;
		WeightsStore9[614] <= Wgt_9_614;
		WeightsStore9[615] <= Wgt_9_615;
		WeightsStore9[616] <= Wgt_9_616;
		WeightsStore9[617] <= Wgt_9_617;
		WeightsStore9[618] <= Wgt_9_618;
		WeightsStore9[619] <= Wgt_9_619;
		WeightsStore9[620] <= Wgt_9_620;
		WeightsStore9[621] <= Wgt_9_621;
		WeightsStore9[622] <= Wgt_9_622;
		WeightsStore9[623] <= Wgt_9_623;
		WeightsStore9[624] <= Wgt_9_624;
		WeightsStore9[625] <= Wgt_9_625;
		WeightsStore9[626] <= Wgt_9_626;
		WeightsStore9[627] <= Wgt_9_627;
		WeightsStore9[628] <= Wgt_9_628;
		WeightsStore9[629] <= Wgt_9_629;
		WeightsStore9[630] <= Wgt_9_630;
		WeightsStore9[631] <= Wgt_9_631;
		WeightsStore9[632] <= Wgt_9_632;
		WeightsStore9[633] <= Wgt_9_633;
		WeightsStore9[634] <= Wgt_9_634;
		WeightsStore9[635] <= Wgt_9_635;
		WeightsStore9[636] <= Wgt_9_636;
		WeightsStore9[637] <= Wgt_9_637;
		WeightsStore9[638] <= Wgt_9_638;
		WeightsStore9[639] <= Wgt_9_639;
		WeightsStore9[640] <= Wgt_9_640;
		WeightsStore9[641] <= Wgt_9_641;
		WeightsStore9[642] <= Wgt_9_642;
		WeightsStore9[643] <= Wgt_9_643;
		WeightsStore9[644] <= Wgt_9_644;
		WeightsStore9[645] <= Wgt_9_645;
		WeightsStore9[646] <= Wgt_9_646;
		WeightsStore9[647] <= Wgt_9_647;
		WeightsStore9[648] <= Wgt_9_648;
		WeightsStore9[649] <= Wgt_9_649;
		WeightsStore9[650] <= Wgt_9_650;
		WeightsStore9[651] <= Wgt_9_651;
		WeightsStore9[652] <= Wgt_9_652;
		WeightsStore9[653] <= Wgt_9_653;
		WeightsStore9[654] <= Wgt_9_654;
		WeightsStore9[655] <= Wgt_9_655;
		WeightsStore9[656] <= Wgt_9_656;
		WeightsStore9[657] <= Wgt_9_657;
		WeightsStore9[658] <= Wgt_9_658;
		WeightsStore9[659] <= Wgt_9_659;
		WeightsStore9[660] <= Wgt_9_660;
		WeightsStore9[661] <= Wgt_9_661;
		WeightsStore9[662] <= Wgt_9_662;
		WeightsStore9[663] <= Wgt_9_663;
		WeightsStore9[664] <= Wgt_9_664;
		WeightsStore9[665] <= Wgt_9_665;
		WeightsStore9[666] <= Wgt_9_666;
		WeightsStore9[667] <= Wgt_9_667;
		WeightsStore9[668] <= Wgt_9_668;
		WeightsStore9[669] <= Wgt_9_669;
		WeightsStore9[670] <= Wgt_9_670;
		WeightsStore9[671] <= Wgt_9_671;
		WeightsStore9[672] <= Wgt_9_672;
		WeightsStore9[673] <= Wgt_9_673;
		WeightsStore9[674] <= Wgt_9_674;
		WeightsStore9[675] <= Wgt_9_675;
		WeightsStore9[676] <= Wgt_9_676;
		WeightsStore9[677] <= Wgt_9_677;
		WeightsStore9[678] <= Wgt_9_678;
		WeightsStore9[679] <= Wgt_9_679;
		WeightsStore9[680] <= Wgt_9_680;
		WeightsStore9[681] <= Wgt_9_681;
		WeightsStore9[682] <= Wgt_9_682;
		WeightsStore9[683] <= Wgt_9_683;
		WeightsStore9[684] <= Wgt_9_684;
		WeightsStore9[685] <= Wgt_9_685;
		WeightsStore9[686] <= Wgt_9_686;
		WeightsStore9[687] <= Wgt_9_687;
		WeightsStore9[688] <= Wgt_9_688;
		WeightsStore9[689] <= Wgt_9_689;
		WeightsStore9[690] <= Wgt_9_690;
		WeightsStore9[691] <= Wgt_9_691;
		WeightsStore9[692] <= Wgt_9_692;
		WeightsStore9[693] <= Wgt_9_693;
		WeightsStore9[694] <= Wgt_9_694;
		WeightsStore9[695] <= Wgt_9_695;
		WeightsStore9[696] <= Wgt_9_696;
		WeightsStore9[697] <= Wgt_9_697;
		WeightsStore9[698] <= Wgt_9_698;
		WeightsStore9[699] <= Wgt_9_699;
		WeightsStore9[700] <= Wgt_9_700;
		WeightsStore9[701] <= Wgt_9_701;
		WeightsStore9[702] <= Wgt_9_702;
		WeightsStore9[703] <= Wgt_9_703;
		WeightsStore9[704] <= Wgt_9_704;
		WeightsStore9[705] <= Wgt_9_705;
		WeightsStore9[706] <= Wgt_9_706;
		WeightsStore9[707] <= Wgt_9_707;
		WeightsStore9[708] <= Wgt_9_708;
		WeightsStore9[709] <= Wgt_9_709;
		WeightsStore9[710] <= Wgt_9_710;
		WeightsStore9[711] <= Wgt_9_711;
		WeightsStore9[712] <= Wgt_9_712;
		WeightsStore9[713] <= Wgt_9_713;
		WeightsStore9[714] <= Wgt_9_714;
		WeightsStore9[715] <= Wgt_9_715;
		WeightsStore9[716] <= Wgt_9_716;
		WeightsStore9[717] <= Wgt_9_717;
		WeightsStore9[718] <= Wgt_9_718;
		WeightsStore9[719] <= Wgt_9_719;
		WeightsStore9[720] <= Wgt_9_720;
		WeightsStore9[721] <= Wgt_9_721;
		WeightsStore9[722] <= Wgt_9_722;
		WeightsStore9[723] <= Wgt_9_723;
		WeightsStore9[724] <= Wgt_9_724;
		WeightsStore9[725] <= Wgt_9_725;
		WeightsStore9[726] <= Wgt_9_726;
		WeightsStore9[727] <= Wgt_9_727;
		WeightsStore9[728] <= Wgt_9_728;
		WeightsStore9[729] <= Wgt_9_729;
		WeightsStore9[730] <= Wgt_9_730;
		WeightsStore9[731] <= Wgt_9_731;
		WeightsStore9[732] <= Wgt_9_732;
		WeightsStore9[733] <= Wgt_9_733;
		WeightsStore9[734] <= Wgt_9_734;
		WeightsStore9[735] <= Wgt_9_735;
		WeightsStore9[736] <= Wgt_9_736;
		WeightsStore9[737] <= Wgt_9_737;
		WeightsStore9[738] <= Wgt_9_738;
		WeightsStore9[739] <= Wgt_9_739;
		WeightsStore9[740] <= Wgt_9_740;
		WeightsStore9[741] <= Wgt_9_741;
		WeightsStore9[742] <= Wgt_9_742;
		WeightsStore9[743] <= Wgt_9_743;
		WeightsStore9[744] <= Wgt_9_744;
		WeightsStore9[745] <= Wgt_9_745;
		WeightsStore9[746] <= Wgt_9_746;
		WeightsStore9[747] <= Wgt_9_747;
		WeightsStore9[748] <= Wgt_9_748;
		WeightsStore9[749] <= Wgt_9_749;
		WeightsStore9[750] <= Wgt_9_750;
		WeightsStore9[751] <= Wgt_9_751;
		WeightsStore9[752] <= Wgt_9_752;
		WeightsStore9[753] <= Wgt_9_753;
		WeightsStore9[754] <= Wgt_9_754;
		WeightsStore9[755] <= Wgt_9_755;
		WeightsStore9[756] <= Wgt_9_756;
		WeightsStore9[757] <= Wgt_9_757;
		WeightsStore9[758] <= Wgt_9_758;
		WeightsStore9[759] <= Wgt_9_759;
		WeightsStore9[760] <= Wgt_9_760;
		WeightsStore9[761] <= Wgt_9_761;
		WeightsStore9[762] <= Wgt_9_762;
		WeightsStore9[763] <= Wgt_9_763;
		WeightsStore9[764] <= Wgt_9_764;
		WeightsStore9[765] <= Wgt_9_765;
		WeightsStore9[766] <= Wgt_9_766;
		WeightsStore9[767] <= Wgt_9_767;
		WeightsStore9[768] <= Wgt_9_768;
		WeightsStore9[769] <= Wgt_9_769;
		WeightsStore9[770] <= Wgt_9_770;
		WeightsStore9[771] <= Wgt_9_771;
		WeightsStore9[772] <= Wgt_9_772;
		WeightsStore9[773] <= Wgt_9_773;
		WeightsStore9[774] <= Wgt_9_774;
		WeightsStore9[775] <= Wgt_9_775;
		WeightsStore9[776] <= Wgt_9_776;
		WeightsStore9[777] <= Wgt_9_777;
		WeightsStore9[778] <= Wgt_9_778;
		WeightsStore9[779] <= Wgt_9_779;
		WeightsStore9[780] <= Wgt_9_780;
		WeightsStore9[781] <= Wgt_9_781;
		WeightsStore9[782] <= Wgt_9_782;
		WeightsStore9[783] <= Wgt_9_783;
		WeightsStore9[784] <= Wgt_9_784;
	end else begin
		internalReset = 1'b1;
		switchCounter <= switchCounter + 32'd1;
		if(switchCounter == 32'd0)begin
		end else if(switchCounter == 32'd6)begin
			PixelsStore[0] <= PixelsStore[28];
			PixelsStore[1] <= PixelsStore[29];
			PixelsStore[2] <= PixelsStore[30];
			PixelsStore[3] <= PixelsStore[31];
			PixelsStore[4] <= PixelsStore[32];
			PixelsStore[5] <= PixelsStore[33];
			PixelsStore[6] <= PixelsStore[34];
			PixelsStore[7] <= PixelsStore[35];
			PixelsStore[8] <= PixelsStore[36];
			PixelsStore[9] <= PixelsStore[37];
			PixelsStore[10] <= PixelsStore[38];
			PixelsStore[11] <= PixelsStore[39];
			PixelsStore[12] <= PixelsStore[40];
			PixelsStore[13] <= PixelsStore[41];
			PixelsStore[14] <= PixelsStore[42];
			PixelsStore[15] <= PixelsStore[43];
			PixelsStore[16] <= PixelsStore[44];
			PixelsStore[17] <= PixelsStore[45];
			PixelsStore[18] <= PixelsStore[46];
			PixelsStore[19] <= PixelsStore[47];
			PixelsStore[20] <= PixelsStore[48];
			PixelsStore[21] <= PixelsStore[49];
			PixelsStore[22] <= PixelsStore[50];
			PixelsStore[23] <= PixelsStore[51];
			PixelsStore[24] <= PixelsStore[52];
			PixelsStore[25] <= PixelsStore[53];
			PixelsStore[26] <= PixelsStore[54];
			PixelsStore[27] <= PixelsStore[55];
			WeightsStore0[0] <= WeightsStore0[28];
			WeightsStore0[1] <= WeightsStore0[29];
			WeightsStore0[2] <= WeightsStore0[30];
			WeightsStore0[3] <= WeightsStore0[31];
			WeightsStore0[4] <= WeightsStore0[32];
			WeightsStore0[5] <= WeightsStore0[33];
			WeightsStore0[6] <= WeightsStore0[34];
			WeightsStore0[7] <= WeightsStore0[35];
			WeightsStore0[8] <= WeightsStore0[36];
			WeightsStore0[9] <= WeightsStore0[37];
			WeightsStore0[10] <= WeightsStore0[38];
			WeightsStore0[11] <= WeightsStore0[39];
			WeightsStore0[12] <= WeightsStore0[40];
			WeightsStore0[13] <= WeightsStore0[41];
			WeightsStore0[14] <= WeightsStore0[42];
			WeightsStore0[15] <= WeightsStore0[43];
			WeightsStore0[16] <= WeightsStore0[44];
			WeightsStore0[17] <= WeightsStore0[45];
			WeightsStore0[18] <= WeightsStore0[46];
			WeightsStore0[19] <= WeightsStore0[47];
			WeightsStore0[20] <= WeightsStore0[48];
			WeightsStore0[21] <= WeightsStore0[49];
			WeightsStore0[22] <= WeightsStore0[50];
			WeightsStore0[23] <= WeightsStore0[51];
			WeightsStore0[24] <= WeightsStore0[52];
			WeightsStore0[25] <= WeightsStore0[53];
			WeightsStore0[26] <= WeightsStore0[54];
			WeightsStore0[27] <= WeightsStore0[55];
			WeightsStore1[0] <= WeightsStore1[28];
			WeightsStore1[1] <= WeightsStore1[29];
			WeightsStore1[2] <= WeightsStore1[30];
			WeightsStore1[3] <= WeightsStore1[31];
			WeightsStore1[4] <= WeightsStore1[32];
			WeightsStore1[5] <= WeightsStore1[33];
			WeightsStore1[6] <= WeightsStore1[34];
			WeightsStore1[7] <= WeightsStore1[35];
			WeightsStore1[8] <= WeightsStore1[36];
			WeightsStore1[9] <= WeightsStore1[37];
			WeightsStore1[10] <= WeightsStore1[38];
			WeightsStore1[11] <= WeightsStore1[39];
			WeightsStore1[12] <= WeightsStore1[40];
			WeightsStore1[13] <= WeightsStore1[41];
			WeightsStore1[14] <= WeightsStore1[42];
			WeightsStore1[15] <= WeightsStore1[43];
			WeightsStore1[16] <= WeightsStore1[44];
			WeightsStore1[17] <= WeightsStore1[45];
			WeightsStore1[18] <= WeightsStore1[46];
			WeightsStore1[19] <= WeightsStore1[47];
			WeightsStore1[20] <= WeightsStore1[48];
			WeightsStore1[21] <= WeightsStore1[49];
			WeightsStore1[22] <= WeightsStore1[50];
			WeightsStore1[23] <= WeightsStore1[51];
			WeightsStore1[24] <= WeightsStore1[52];
			WeightsStore1[25] <= WeightsStore1[53];
			WeightsStore1[26] <= WeightsStore1[54];
			WeightsStore1[27] <= WeightsStore1[55];
			WeightsStore2[0] <= WeightsStore2[28];
			WeightsStore2[1] <= WeightsStore2[29];
			WeightsStore2[2] <= WeightsStore2[30];
			WeightsStore2[3] <= WeightsStore2[31];
			WeightsStore2[4] <= WeightsStore2[32];
			WeightsStore2[5] <= WeightsStore2[33];
			WeightsStore2[6] <= WeightsStore2[34];
			WeightsStore2[7] <= WeightsStore2[35];
			WeightsStore2[8] <= WeightsStore2[36];
			WeightsStore2[9] <= WeightsStore2[37];
			WeightsStore2[10] <= WeightsStore2[38];
			WeightsStore2[11] <= WeightsStore2[39];
			WeightsStore2[12] <= WeightsStore2[40];
			WeightsStore2[13] <= WeightsStore2[41];
			WeightsStore2[14] <= WeightsStore2[42];
			WeightsStore2[15] <= WeightsStore2[43];
			WeightsStore2[16] <= WeightsStore2[44];
			WeightsStore2[17] <= WeightsStore2[45];
			WeightsStore2[18] <= WeightsStore2[46];
			WeightsStore2[19] <= WeightsStore2[47];
			WeightsStore2[20] <= WeightsStore2[48];
			WeightsStore2[21] <= WeightsStore2[49];
			WeightsStore2[22] <= WeightsStore2[50];
			WeightsStore2[23] <= WeightsStore2[51];
			WeightsStore2[24] <= WeightsStore2[52];
			WeightsStore2[25] <= WeightsStore2[53];
			WeightsStore2[26] <= WeightsStore2[54];
			WeightsStore2[27] <= WeightsStore2[55];
			WeightsStore3[0] <= WeightsStore3[28];
			WeightsStore3[1] <= WeightsStore3[29];
			WeightsStore3[2] <= WeightsStore3[30];
			WeightsStore3[3] <= WeightsStore3[31];
			WeightsStore3[4] <= WeightsStore3[32];
			WeightsStore3[5] <= WeightsStore3[33];
			WeightsStore3[6] <= WeightsStore3[34];
			WeightsStore3[7] <= WeightsStore3[35];
			WeightsStore3[8] <= WeightsStore3[36];
			WeightsStore3[9] <= WeightsStore3[37];
			WeightsStore3[10] <= WeightsStore3[38];
			WeightsStore3[11] <= WeightsStore3[39];
			WeightsStore3[12] <= WeightsStore3[40];
			WeightsStore3[13] <= WeightsStore3[41];
			WeightsStore3[14] <= WeightsStore3[42];
			WeightsStore3[15] <= WeightsStore3[43];
			WeightsStore3[16] <= WeightsStore3[44];
			WeightsStore3[17] <= WeightsStore3[45];
			WeightsStore3[18] <= WeightsStore3[46];
			WeightsStore3[19] <= WeightsStore3[47];
			WeightsStore3[20] <= WeightsStore3[48];
			WeightsStore3[21] <= WeightsStore3[49];
			WeightsStore3[22] <= WeightsStore3[50];
			WeightsStore3[23] <= WeightsStore3[51];
			WeightsStore3[24] <= WeightsStore3[52];
			WeightsStore3[25] <= WeightsStore3[53];
			WeightsStore3[26] <= WeightsStore3[54];
			WeightsStore3[27] <= WeightsStore3[55];
			WeightsStore4[0] <= WeightsStore4[28];
			WeightsStore4[1] <= WeightsStore4[29];
			WeightsStore4[2] <= WeightsStore4[30];
			WeightsStore4[3] <= WeightsStore4[31];
			WeightsStore4[4] <= WeightsStore4[32];
			WeightsStore4[5] <= WeightsStore4[33];
			WeightsStore4[6] <= WeightsStore4[34];
			WeightsStore4[7] <= WeightsStore4[35];
			WeightsStore4[8] <= WeightsStore4[36];
			WeightsStore4[9] <= WeightsStore4[37];
			WeightsStore4[10] <= WeightsStore4[38];
			WeightsStore4[11] <= WeightsStore4[39];
			WeightsStore4[12] <= WeightsStore4[40];
			WeightsStore4[13] <= WeightsStore4[41];
			WeightsStore4[14] <= WeightsStore4[42];
			WeightsStore4[15] <= WeightsStore4[43];
			WeightsStore4[16] <= WeightsStore4[44];
			WeightsStore4[17] <= WeightsStore4[45];
			WeightsStore4[18] <= WeightsStore4[46];
			WeightsStore4[19] <= WeightsStore4[47];
			WeightsStore4[20] <= WeightsStore4[48];
			WeightsStore4[21] <= WeightsStore4[49];
			WeightsStore4[22] <= WeightsStore4[50];
			WeightsStore4[23] <= WeightsStore4[51];
			WeightsStore4[24] <= WeightsStore4[52];
			WeightsStore4[25] <= WeightsStore4[53];
			WeightsStore4[26] <= WeightsStore4[54];
			WeightsStore4[27] <= WeightsStore4[55];
			WeightsStore5[0] <= WeightsStore5[28];
			WeightsStore5[1] <= WeightsStore5[29];
			WeightsStore5[2] <= WeightsStore5[30];
			WeightsStore5[3] <= WeightsStore5[31];
			WeightsStore5[4] <= WeightsStore5[32];
			WeightsStore5[5] <= WeightsStore5[33];
			WeightsStore5[6] <= WeightsStore5[34];
			WeightsStore5[7] <= WeightsStore5[35];
			WeightsStore5[8] <= WeightsStore5[36];
			WeightsStore5[9] <= WeightsStore5[37];
			WeightsStore5[10] <= WeightsStore5[38];
			WeightsStore5[11] <= WeightsStore5[39];
			WeightsStore5[12] <= WeightsStore5[40];
			WeightsStore5[13] <= WeightsStore5[41];
			WeightsStore5[14] <= WeightsStore5[42];
			WeightsStore5[15] <= WeightsStore5[43];
			WeightsStore5[16] <= WeightsStore5[44];
			WeightsStore5[17] <= WeightsStore5[45];
			WeightsStore5[18] <= WeightsStore5[46];
			WeightsStore5[19] <= WeightsStore5[47];
			WeightsStore5[20] <= WeightsStore5[48];
			WeightsStore5[21] <= WeightsStore5[49];
			WeightsStore5[22] <= WeightsStore5[50];
			WeightsStore5[23] <= WeightsStore5[51];
			WeightsStore5[24] <= WeightsStore5[52];
			WeightsStore5[25] <= WeightsStore5[53];
			WeightsStore5[26] <= WeightsStore5[54];
			WeightsStore5[27] <= WeightsStore5[55];
			WeightsStore6[0] <= WeightsStore6[28];
			WeightsStore6[1] <= WeightsStore6[29];
			WeightsStore6[2] <= WeightsStore6[30];
			WeightsStore6[3] <= WeightsStore6[31];
			WeightsStore6[4] <= WeightsStore6[32];
			WeightsStore6[5] <= WeightsStore6[33];
			WeightsStore6[6] <= WeightsStore6[34];
			WeightsStore6[7] <= WeightsStore6[35];
			WeightsStore6[8] <= WeightsStore6[36];
			WeightsStore6[9] <= WeightsStore6[37];
			WeightsStore6[10] <= WeightsStore6[38];
			WeightsStore6[11] <= WeightsStore6[39];
			WeightsStore6[12] <= WeightsStore6[40];
			WeightsStore6[13] <= WeightsStore6[41];
			WeightsStore6[14] <= WeightsStore6[42];
			WeightsStore6[15] <= WeightsStore6[43];
			WeightsStore6[16] <= WeightsStore6[44];
			WeightsStore6[17] <= WeightsStore6[45];
			WeightsStore6[18] <= WeightsStore6[46];
			WeightsStore6[19] <= WeightsStore6[47];
			WeightsStore6[20] <= WeightsStore6[48];
			WeightsStore6[21] <= WeightsStore6[49];
			WeightsStore6[22] <= WeightsStore6[50];
			WeightsStore6[23] <= WeightsStore6[51];
			WeightsStore6[24] <= WeightsStore6[52];
			WeightsStore6[25] <= WeightsStore6[53];
			WeightsStore6[26] <= WeightsStore6[54];
			WeightsStore6[27] <= WeightsStore6[55];
			WeightsStore7[0] <= WeightsStore7[28];
			WeightsStore7[1] <= WeightsStore7[29];
			WeightsStore7[2] <= WeightsStore7[30];
			WeightsStore7[3] <= WeightsStore7[31];
			WeightsStore7[4] <= WeightsStore7[32];
			WeightsStore7[5] <= WeightsStore7[33];
			WeightsStore7[6] <= WeightsStore7[34];
			WeightsStore7[7] <= WeightsStore7[35];
			WeightsStore7[8] <= WeightsStore7[36];
			WeightsStore7[9] <= WeightsStore7[37];
			WeightsStore7[10] <= WeightsStore7[38];
			WeightsStore7[11] <= WeightsStore7[39];
			WeightsStore7[12] <= WeightsStore7[40];
			WeightsStore7[13] <= WeightsStore7[41];
			WeightsStore7[14] <= WeightsStore7[42];
			WeightsStore7[15] <= WeightsStore7[43];
			WeightsStore7[16] <= WeightsStore7[44];
			WeightsStore7[17] <= WeightsStore7[45];
			WeightsStore7[18] <= WeightsStore7[46];
			WeightsStore7[19] <= WeightsStore7[47];
			WeightsStore7[20] <= WeightsStore7[48];
			WeightsStore7[21] <= WeightsStore7[49];
			WeightsStore7[22] <= WeightsStore7[50];
			WeightsStore7[23] <= WeightsStore7[51];
			WeightsStore7[24] <= WeightsStore7[52];
			WeightsStore7[25] <= WeightsStore7[53];
			WeightsStore7[26] <= WeightsStore7[54];
			WeightsStore7[27] <= WeightsStore7[55];
			WeightsStore8[0] <= WeightsStore8[28];
			WeightsStore8[1] <= WeightsStore8[29];
			WeightsStore8[2] <= WeightsStore8[30];
			WeightsStore8[3] <= WeightsStore8[31];
			WeightsStore8[4] <= WeightsStore8[32];
			WeightsStore8[5] <= WeightsStore8[33];
			WeightsStore8[6] <= WeightsStore8[34];
			WeightsStore8[7] <= WeightsStore8[35];
			WeightsStore8[8] <= WeightsStore8[36];
			WeightsStore8[9] <= WeightsStore8[37];
			WeightsStore8[10] <= WeightsStore8[38];
			WeightsStore8[11] <= WeightsStore8[39];
			WeightsStore8[12] <= WeightsStore8[40];
			WeightsStore8[13] <= WeightsStore8[41];
			WeightsStore8[14] <= WeightsStore8[42];
			WeightsStore8[15] <= WeightsStore8[43];
			WeightsStore8[16] <= WeightsStore8[44];
			WeightsStore8[17] <= WeightsStore8[45];
			WeightsStore8[18] <= WeightsStore8[46];
			WeightsStore8[19] <= WeightsStore8[47];
			WeightsStore8[20] <= WeightsStore8[48];
			WeightsStore8[21] <= WeightsStore8[49];
			WeightsStore8[22] <= WeightsStore8[50];
			WeightsStore8[23] <= WeightsStore8[51];
			WeightsStore8[24] <= WeightsStore8[52];
			WeightsStore8[25] <= WeightsStore8[53];
			WeightsStore8[26] <= WeightsStore8[54];
			WeightsStore8[27] <= WeightsStore8[55];
			WeightsStore9[0] <= WeightsStore9[28];
			WeightsStore9[1] <= WeightsStore9[29];
			WeightsStore9[2] <= WeightsStore9[30];
			WeightsStore9[3] <= WeightsStore9[31];
			WeightsStore9[4] <= WeightsStore9[32];
			WeightsStore9[5] <= WeightsStore9[33];
			WeightsStore9[6] <= WeightsStore9[34];
			WeightsStore9[7] <= WeightsStore9[35];
			WeightsStore9[8] <= WeightsStore9[36];
			WeightsStore9[9] <= WeightsStore9[37];
			WeightsStore9[10] <= WeightsStore9[38];
			WeightsStore9[11] <= WeightsStore9[39];
			WeightsStore9[12] <= WeightsStore9[40];
			WeightsStore9[13] <= WeightsStore9[41];
			WeightsStore9[14] <= WeightsStore9[42];
			WeightsStore9[15] <= WeightsStore9[43];
			WeightsStore9[16] <= WeightsStore9[44];
			WeightsStore9[17] <= WeightsStore9[45];
			WeightsStore9[18] <= WeightsStore9[46];
			WeightsStore9[19] <= WeightsStore9[47];
			WeightsStore9[20] <= WeightsStore9[48];
			WeightsStore9[21] <= WeightsStore9[49];
			WeightsStore9[22] <= WeightsStore9[50];
			WeightsStore9[23] <= WeightsStore9[51];
			WeightsStore9[24] <= WeightsStore9[52];
			WeightsStore9[25] <= WeightsStore9[53];
			WeightsStore9[26] <= WeightsStore9[54];
			WeightsStore9[27] <= WeightsStore9[55];
		end else if(switchCounter == 32'd13)begin
			PixelsStore[0] <= PixelsStore[56];
			PixelsStore[1] <= PixelsStore[57];
			PixelsStore[2] <= PixelsStore[58];
			PixelsStore[3] <= PixelsStore[59];
			PixelsStore[4] <= PixelsStore[60];
			PixelsStore[5] <= PixelsStore[61];
			PixelsStore[6] <= PixelsStore[62];
			PixelsStore[7] <= PixelsStore[63];
			PixelsStore[8] <= PixelsStore[64];
			PixelsStore[9] <= PixelsStore[65];
			PixelsStore[10] <= PixelsStore[66];
			PixelsStore[11] <= PixelsStore[67];
			PixelsStore[12] <= PixelsStore[68];
			PixelsStore[13] <= PixelsStore[69];
			PixelsStore[14] <= PixelsStore[70];
			PixelsStore[15] <= PixelsStore[71];
			PixelsStore[16] <= PixelsStore[72];
			PixelsStore[17] <= PixelsStore[73];
			PixelsStore[18] <= PixelsStore[74];
			PixelsStore[19] <= PixelsStore[75];
			PixelsStore[20] <= PixelsStore[76];
			PixelsStore[21] <= PixelsStore[77];
			PixelsStore[22] <= PixelsStore[78];
			PixelsStore[23] <= PixelsStore[79];
			PixelsStore[24] <= PixelsStore[80];
			PixelsStore[25] <= PixelsStore[81];
			PixelsStore[26] <= PixelsStore[82];
			PixelsStore[27] <= PixelsStore[83];
			WeightsStore0[0] <= WeightsStore0[56];
			WeightsStore0[1] <= WeightsStore0[57];
			WeightsStore0[2] <= WeightsStore0[58];
			WeightsStore0[3] <= WeightsStore0[59];
			WeightsStore0[4] <= WeightsStore0[60];
			WeightsStore0[5] <= WeightsStore0[61];
			WeightsStore0[6] <= WeightsStore0[62];
			WeightsStore0[7] <= WeightsStore0[63];
			WeightsStore0[8] <= WeightsStore0[64];
			WeightsStore0[9] <= WeightsStore0[65];
			WeightsStore0[10] <= WeightsStore0[66];
			WeightsStore0[11] <= WeightsStore0[67];
			WeightsStore0[12] <= WeightsStore0[68];
			WeightsStore0[13] <= WeightsStore0[69];
			WeightsStore0[14] <= WeightsStore0[70];
			WeightsStore0[15] <= WeightsStore0[71];
			WeightsStore0[16] <= WeightsStore0[72];
			WeightsStore0[17] <= WeightsStore0[73];
			WeightsStore0[18] <= WeightsStore0[74];
			WeightsStore0[19] <= WeightsStore0[75];
			WeightsStore0[20] <= WeightsStore0[76];
			WeightsStore0[21] <= WeightsStore0[77];
			WeightsStore0[22] <= WeightsStore0[78];
			WeightsStore0[23] <= WeightsStore0[79];
			WeightsStore0[24] <= WeightsStore0[80];
			WeightsStore0[25] <= WeightsStore0[81];
			WeightsStore0[26] <= WeightsStore0[82];
			WeightsStore0[27] <= WeightsStore0[83];
			WeightsStore1[0] <= WeightsStore1[56];
			WeightsStore1[1] <= WeightsStore1[57];
			WeightsStore1[2] <= WeightsStore1[58];
			WeightsStore1[3] <= WeightsStore1[59];
			WeightsStore1[4] <= WeightsStore1[60];
			WeightsStore1[5] <= WeightsStore1[61];
			WeightsStore1[6] <= WeightsStore1[62];
			WeightsStore1[7] <= WeightsStore1[63];
			WeightsStore1[8] <= WeightsStore1[64];
			WeightsStore1[9] <= WeightsStore1[65];
			WeightsStore1[10] <= WeightsStore1[66];
			WeightsStore1[11] <= WeightsStore1[67];
			WeightsStore1[12] <= WeightsStore1[68];
			WeightsStore1[13] <= WeightsStore1[69];
			WeightsStore1[14] <= WeightsStore1[70];
			WeightsStore1[15] <= WeightsStore1[71];
			WeightsStore1[16] <= WeightsStore1[72];
			WeightsStore1[17] <= WeightsStore1[73];
			WeightsStore1[18] <= WeightsStore1[74];
			WeightsStore1[19] <= WeightsStore1[75];
			WeightsStore1[20] <= WeightsStore1[76];
			WeightsStore1[21] <= WeightsStore1[77];
			WeightsStore1[22] <= WeightsStore1[78];
			WeightsStore1[23] <= WeightsStore1[79];
			WeightsStore1[24] <= WeightsStore1[80];
			WeightsStore1[25] <= WeightsStore1[81];
			WeightsStore1[26] <= WeightsStore1[82];
			WeightsStore1[27] <= WeightsStore1[83];
			WeightsStore2[0] <= WeightsStore2[56];
			WeightsStore2[1] <= WeightsStore2[57];
			WeightsStore2[2] <= WeightsStore2[58];
			WeightsStore2[3] <= WeightsStore2[59];
			WeightsStore2[4] <= WeightsStore2[60];
			WeightsStore2[5] <= WeightsStore2[61];
			WeightsStore2[6] <= WeightsStore2[62];
			WeightsStore2[7] <= WeightsStore2[63];
			WeightsStore2[8] <= WeightsStore2[64];
			WeightsStore2[9] <= WeightsStore2[65];
			WeightsStore2[10] <= WeightsStore2[66];
			WeightsStore2[11] <= WeightsStore2[67];
			WeightsStore2[12] <= WeightsStore2[68];
			WeightsStore2[13] <= WeightsStore2[69];
			WeightsStore2[14] <= WeightsStore2[70];
			WeightsStore2[15] <= WeightsStore2[71];
			WeightsStore2[16] <= WeightsStore2[72];
			WeightsStore2[17] <= WeightsStore2[73];
			WeightsStore2[18] <= WeightsStore2[74];
			WeightsStore2[19] <= WeightsStore2[75];
			WeightsStore2[20] <= WeightsStore2[76];
			WeightsStore2[21] <= WeightsStore2[77];
			WeightsStore2[22] <= WeightsStore2[78];
			WeightsStore2[23] <= WeightsStore2[79];
			WeightsStore2[24] <= WeightsStore2[80];
			WeightsStore2[25] <= WeightsStore2[81];
			WeightsStore2[26] <= WeightsStore2[82];
			WeightsStore2[27] <= WeightsStore2[83];
			WeightsStore3[0] <= WeightsStore3[56];
			WeightsStore3[1] <= WeightsStore3[57];
			WeightsStore3[2] <= WeightsStore3[58];
			WeightsStore3[3] <= WeightsStore3[59];
			WeightsStore3[4] <= WeightsStore3[60];
			WeightsStore3[5] <= WeightsStore3[61];
			WeightsStore3[6] <= WeightsStore3[62];
			WeightsStore3[7] <= WeightsStore3[63];
			WeightsStore3[8] <= WeightsStore3[64];
			WeightsStore3[9] <= WeightsStore3[65];
			WeightsStore3[10] <= WeightsStore3[66];
			WeightsStore3[11] <= WeightsStore3[67];
			WeightsStore3[12] <= WeightsStore3[68];
			WeightsStore3[13] <= WeightsStore3[69];
			WeightsStore3[14] <= WeightsStore3[70];
			WeightsStore3[15] <= WeightsStore3[71];
			WeightsStore3[16] <= WeightsStore3[72];
			WeightsStore3[17] <= WeightsStore3[73];
			WeightsStore3[18] <= WeightsStore3[74];
			WeightsStore3[19] <= WeightsStore3[75];
			WeightsStore3[20] <= WeightsStore3[76];
			WeightsStore3[21] <= WeightsStore3[77];
			WeightsStore3[22] <= WeightsStore3[78];
			WeightsStore3[23] <= WeightsStore3[79];
			WeightsStore3[24] <= WeightsStore3[80];
			WeightsStore3[25] <= WeightsStore3[81];
			WeightsStore3[26] <= WeightsStore3[82];
			WeightsStore3[27] <= WeightsStore3[83];
			WeightsStore4[0] <= WeightsStore4[56];
			WeightsStore4[1] <= WeightsStore4[57];
			WeightsStore4[2] <= WeightsStore4[58];
			WeightsStore4[3] <= WeightsStore4[59];
			WeightsStore4[4] <= WeightsStore4[60];
			WeightsStore4[5] <= WeightsStore4[61];
			WeightsStore4[6] <= WeightsStore4[62];
			WeightsStore4[7] <= WeightsStore4[63];
			WeightsStore4[8] <= WeightsStore4[64];
			WeightsStore4[9] <= WeightsStore4[65];
			WeightsStore4[10] <= WeightsStore4[66];
			WeightsStore4[11] <= WeightsStore4[67];
			WeightsStore4[12] <= WeightsStore4[68];
			WeightsStore4[13] <= WeightsStore4[69];
			WeightsStore4[14] <= WeightsStore4[70];
			WeightsStore4[15] <= WeightsStore4[71];
			WeightsStore4[16] <= WeightsStore4[72];
			WeightsStore4[17] <= WeightsStore4[73];
			WeightsStore4[18] <= WeightsStore4[74];
			WeightsStore4[19] <= WeightsStore4[75];
			WeightsStore4[20] <= WeightsStore4[76];
			WeightsStore4[21] <= WeightsStore4[77];
			WeightsStore4[22] <= WeightsStore4[78];
			WeightsStore4[23] <= WeightsStore4[79];
			WeightsStore4[24] <= WeightsStore4[80];
			WeightsStore4[25] <= WeightsStore4[81];
			WeightsStore4[26] <= WeightsStore4[82];
			WeightsStore4[27] <= WeightsStore4[83];
			WeightsStore5[0] <= WeightsStore5[56];
			WeightsStore5[1] <= WeightsStore5[57];
			WeightsStore5[2] <= WeightsStore5[58];
			WeightsStore5[3] <= WeightsStore5[59];
			WeightsStore5[4] <= WeightsStore5[60];
			WeightsStore5[5] <= WeightsStore5[61];
			WeightsStore5[6] <= WeightsStore5[62];
			WeightsStore5[7] <= WeightsStore5[63];
			WeightsStore5[8] <= WeightsStore5[64];
			WeightsStore5[9] <= WeightsStore5[65];
			WeightsStore5[10] <= WeightsStore5[66];
			WeightsStore5[11] <= WeightsStore5[67];
			WeightsStore5[12] <= WeightsStore5[68];
			WeightsStore5[13] <= WeightsStore5[69];
			WeightsStore5[14] <= WeightsStore5[70];
			WeightsStore5[15] <= WeightsStore5[71];
			WeightsStore5[16] <= WeightsStore5[72];
			WeightsStore5[17] <= WeightsStore5[73];
			WeightsStore5[18] <= WeightsStore5[74];
			WeightsStore5[19] <= WeightsStore5[75];
			WeightsStore5[20] <= WeightsStore5[76];
			WeightsStore5[21] <= WeightsStore5[77];
			WeightsStore5[22] <= WeightsStore5[78];
			WeightsStore5[23] <= WeightsStore5[79];
			WeightsStore5[24] <= WeightsStore5[80];
			WeightsStore5[25] <= WeightsStore5[81];
			WeightsStore5[26] <= WeightsStore5[82];
			WeightsStore5[27] <= WeightsStore5[83];
			WeightsStore6[0] <= WeightsStore6[56];
			WeightsStore6[1] <= WeightsStore6[57];
			WeightsStore6[2] <= WeightsStore6[58];
			WeightsStore6[3] <= WeightsStore6[59];
			WeightsStore6[4] <= WeightsStore6[60];
			WeightsStore6[5] <= WeightsStore6[61];
			WeightsStore6[6] <= WeightsStore6[62];
			WeightsStore6[7] <= WeightsStore6[63];
			WeightsStore6[8] <= WeightsStore6[64];
			WeightsStore6[9] <= WeightsStore6[65];
			WeightsStore6[10] <= WeightsStore6[66];
			WeightsStore6[11] <= WeightsStore6[67];
			WeightsStore6[12] <= WeightsStore6[68];
			WeightsStore6[13] <= WeightsStore6[69];
			WeightsStore6[14] <= WeightsStore6[70];
			WeightsStore6[15] <= WeightsStore6[71];
			WeightsStore6[16] <= WeightsStore6[72];
			WeightsStore6[17] <= WeightsStore6[73];
			WeightsStore6[18] <= WeightsStore6[74];
			WeightsStore6[19] <= WeightsStore6[75];
			WeightsStore6[20] <= WeightsStore6[76];
			WeightsStore6[21] <= WeightsStore6[77];
			WeightsStore6[22] <= WeightsStore6[78];
			WeightsStore6[23] <= WeightsStore6[79];
			WeightsStore6[24] <= WeightsStore6[80];
			WeightsStore6[25] <= WeightsStore6[81];
			WeightsStore6[26] <= WeightsStore6[82];
			WeightsStore6[27] <= WeightsStore6[83];
			WeightsStore7[0] <= WeightsStore7[56];
			WeightsStore7[1] <= WeightsStore7[57];
			WeightsStore7[2] <= WeightsStore7[58];
			WeightsStore7[3] <= WeightsStore7[59];
			WeightsStore7[4] <= WeightsStore7[60];
			WeightsStore7[5] <= WeightsStore7[61];
			WeightsStore7[6] <= WeightsStore7[62];
			WeightsStore7[7] <= WeightsStore7[63];
			WeightsStore7[8] <= WeightsStore7[64];
			WeightsStore7[9] <= WeightsStore7[65];
			WeightsStore7[10] <= WeightsStore7[66];
			WeightsStore7[11] <= WeightsStore7[67];
			WeightsStore7[12] <= WeightsStore7[68];
			WeightsStore7[13] <= WeightsStore7[69];
			WeightsStore7[14] <= WeightsStore7[70];
			WeightsStore7[15] <= WeightsStore7[71];
			WeightsStore7[16] <= WeightsStore7[72];
			WeightsStore7[17] <= WeightsStore7[73];
			WeightsStore7[18] <= WeightsStore7[74];
			WeightsStore7[19] <= WeightsStore7[75];
			WeightsStore7[20] <= WeightsStore7[76];
			WeightsStore7[21] <= WeightsStore7[77];
			WeightsStore7[22] <= WeightsStore7[78];
			WeightsStore7[23] <= WeightsStore7[79];
			WeightsStore7[24] <= WeightsStore7[80];
			WeightsStore7[25] <= WeightsStore7[81];
			WeightsStore7[26] <= WeightsStore7[82];
			WeightsStore7[27] <= WeightsStore7[83];
			WeightsStore8[0] <= WeightsStore8[56];
			WeightsStore8[1] <= WeightsStore8[57];
			WeightsStore8[2] <= WeightsStore8[58];
			WeightsStore8[3] <= WeightsStore8[59];
			WeightsStore8[4] <= WeightsStore8[60];
			WeightsStore8[5] <= WeightsStore8[61];
			WeightsStore8[6] <= WeightsStore8[62];
			WeightsStore8[7] <= WeightsStore8[63];
			WeightsStore8[8] <= WeightsStore8[64];
			WeightsStore8[9] <= WeightsStore8[65];
			WeightsStore8[10] <= WeightsStore8[66];
			WeightsStore8[11] <= WeightsStore8[67];
			WeightsStore8[12] <= WeightsStore8[68];
			WeightsStore8[13] <= WeightsStore8[69];
			WeightsStore8[14] <= WeightsStore8[70];
			WeightsStore8[15] <= WeightsStore8[71];
			WeightsStore8[16] <= WeightsStore8[72];
			WeightsStore8[17] <= WeightsStore8[73];
			WeightsStore8[18] <= WeightsStore8[74];
			WeightsStore8[19] <= WeightsStore8[75];
			WeightsStore8[20] <= WeightsStore8[76];
			WeightsStore8[21] <= WeightsStore8[77];
			WeightsStore8[22] <= WeightsStore8[78];
			WeightsStore8[23] <= WeightsStore8[79];
			WeightsStore8[24] <= WeightsStore8[80];
			WeightsStore8[25] <= WeightsStore8[81];
			WeightsStore8[26] <= WeightsStore8[82];
			WeightsStore8[27] <= WeightsStore8[83];
			WeightsStore9[0] <= WeightsStore9[56];
			WeightsStore9[1] <= WeightsStore9[57];
			WeightsStore9[2] <= WeightsStore9[58];
			WeightsStore9[3] <= WeightsStore9[59];
			WeightsStore9[4] <= WeightsStore9[60];
			WeightsStore9[5] <= WeightsStore9[61];
			WeightsStore9[6] <= WeightsStore9[62];
			WeightsStore9[7] <= WeightsStore9[63];
			WeightsStore9[8] <= WeightsStore9[64];
			WeightsStore9[9] <= WeightsStore9[65];
			WeightsStore9[10] <= WeightsStore9[66];
			WeightsStore9[11] <= WeightsStore9[67];
			WeightsStore9[12] <= WeightsStore9[68];
			WeightsStore9[13] <= WeightsStore9[69];
			WeightsStore9[14] <= WeightsStore9[70];
			WeightsStore9[15] <= WeightsStore9[71];
			WeightsStore9[16] <= WeightsStore9[72];
			WeightsStore9[17] <= WeightsStore9[73];
			WeightsStore9[18] <= WeightsStore9[74];
			WeightsStore9[19] <= WeightsStore9[75];
			WeightsStore9[20] <= WeightsStore9[76];
			WeightsStore9[21] <= WeightsStore9[77];
			WeightsStore9[22] <= WeightsStore9[78];
			WeightsStore9[23] <= WeightsStore9[79];
			WeightsStore9[24] <= WeightsStore9[80];
			WeightsStore9[25] <= WeightsStore9[81];
			WeightsStore9[26] <= WeightsStore9[82];
			WeightsStore9[27] <= WeightsStore9[83];
		end else if(switchCounter == 32'd20)begin
			PixelsStore[0] <= PixelsStore[84];
			PixelsStore[1] <= PixelsStore[85];
			PixelsStore[2] <= PixelsStore[86];
			PixelsStore[3] <= PixelsStore[87];
			PixelsStore[4] <= PixelsStore[88];
			PixelsStore[5] <= PixelsStore[89];
			PixelsStore[6] <= PixelsStore[90];
			PixelsStore[7] <= PixelsStore[91];
			PixelsStore[8] <= PixelsStore[92];
			PixelsStore[9] <= PixelsStore[93];
			PixelsStore[10] <= PixelsStore[94];
			PixelsStore[11] <= PixelsStore[95];
			PixelsStore[12] <= PixelsStore[96];
			PixelsStore[13] <= PixelsStore[97];
			PixelsStore[14] <= PixelsStore[98];
			PixelsStore[15] <= PixelsStore[99];
			PixelsStore[16] <= PixelsStore[100];
			PixelsStore[17] <= PixelsStore[101];
			PixelsStore[18] <= PixelsStore[102];
			PixelsStore[19] <= PixelsStore[103];
			PixelsStore[20] <= PixelsStore[104];
			PixelsStore[21] <= PixelsStore[105];
			PixelsStore[22] <= PixelsStore[106];
			PixelsStore[23] <= PixelsStore[107];
			PixelsStore[24] <= PixelsStore[108];
			PixelsStore[25] <= PixelsStore[109];
			PixelsStore[26] <= PixelsStore[110];
			PixelsStore[27] <= PixelsStore[111];
			WeightsStore0[0] <= WeightsStore0[84];
			WeightsStore0[1] <= WeightsStore0[85];
			WeightsStore0[2] <= WeightsStore0[86];
			WeightsStore0[3] <= WeightsStore0[87];
			WeightsStore0[4] <= WeightsStore0[88];
			WeightsStore0[5] <= WeightsStore0[89];
			WeightsStore0[6] <= WeightsStore0[90];
			WeightsStore0[7] <= WeightsStore0[91];
			WeightsStore0[8] <= WeightsStore0[92];
			WeightsStore0[9] <= WeightsStore0[93];
			WeightsStore0[10] <= WeightsStore0[94];
			WeightsStore0[11] <= WeightsStore0[95];
			WeightsStore0[12] <= WeightsStore0[96];
			WeightsStore0[13] <= WeightsStore0[97];
			WeightsStore0[14] <= WeightsStore0[98];
			WeightsStore0[15] <= WeightsStore0[99];
			WeightsStore0[16] <= WeightsStore0[100];
			WeightsStore0[17] <= WeightsStore0[101];
			WeightsStore0[18] <= WeightsStore0[102];
			WeightsStore0[19] <= WeightsStore0[103];
			WeightsStore0[20] <= WeightsStore0[104];
			WeightsStore0[21] <= WeightsStore0[105];
			WeightsStore0[22] <= WeightsStore0[106];
			WeightsStore0[23] <= WeightsStore0[107];
			WeightsStore0[24] <= WeightsStore0[108];
			WeightsStore0[25] <= WeightsStore0[109];
			WeightsStore0[26] <= WeightsStore0[110];
			WeightsStore0[27] <= WeightsStore0[111];
			WeightsStore1[0] <= WeightsStore1[84];
			WeightsStore1[1] <= WeightsStore1[85];
			WeightsStore1[2] <= WeightsStore1[86];
			WeightsStore1[3] <= WeightsStore1[87];
			WeightsStore1[4] <= WeightsStore1[88];
			WeightsStore1[5] <= WeightsStore1[89];
			WeightsStore1[6] <= WeightsStore1[90];
			WeightsStore1[7] <= WeightsStore1[91];
			WeightsStore1[8] <= WeightsStore1[92];
			WeightsStore1[9] <= WeightsStore1[93];
			WeightsStore1[10] <= WeightsStore1[94];
			WeightsStore1[11] <= WeightsStore1[95];
			WeightsStore1[12] <= WeightsStore1[96];
			WeightsStore1[13] <= WeightsStore1[97];
			WeightsStore1[14] <= WeightsStore1[98];
			WeightsStore1[15] <= WeightsStore1[99];
			WeightsStore1[16] <= WeightsStore1[100];
			WeightsStore1[17] <= WeightsStore1[101];
			WeightsStore1[18] <= WeightsStore1[102];
			WeightsStore1[19] <= WeightsStore1[103];
			WeightsStore1[20] <= WeightsStore1[104];
			WeightsStore1[21] <= WeightsStore1[105];
			WeightsStore1[22] <= WeightsStore1[106];
			WeightsStore1[23] <= WeightsStore1[107];
			WeightsStore1[24] <= WeightsStore1[108];
			WeightsStore1[25] <= WeightsStore1[109];
			WeightsStore1[26] <= WeightsStore1[110];
			WeightsStore1[27] <= WeightsStore1[111];
			WeightsStore2[0] <= WeightsStore2[84];
			WeightsStore2[1] <= WeightsStore2[85];
			WeightsStore2[2] <= WeightsStore2[86];
			WeightsStore2[3] <= WeightsStore2[87];
			WeightsStore2[4] <= WeightsStore2[88];
			WeightsStore2[5] <= WeightsStore2[89];
			WeightsStore2[6] <= WeightsStore2[90];
			WeightsStore2[7] <= WeightsStore2[91];
			WeightsStore2[8] <= WeightsStore2[92];
			WeightsStore2[9] <= WeightsStore2[93];
			WeightsStore2[10] <= WeightsStore2[94];
			WeightsStore2[11] <= WeightsStore2[95];
			WeightsStore2[12] <= WeightsStore2[96];
			WeightsStore2[13] <= WeightsStore2[97];
			WeightsStore2[14] <= WeightsStore2[98];
			WeightsStore2[15] <= WeightsStore2[99];
			WeightsStore2[16] <= WeightsStore2[100];
			WeightsStore2[17] <= WeightsStore2[101];
			WeightsStore2[18] <= WeightsStore2[102];
			WeightsStore2[19] <= WeightsStore2[103];
			WeightsStore2[20] <= WeightsStore2[104];
			WeightsStore2[21] <= WeightsStore2[105];
			WeightsStore2[22] <= WeightsStore2[106];
			WeightsStore2[23] <= WeightsStore2[107];
			WeightsStore2[24] <= WeightsStore2[108];
			WeightsStore2[25] <= WeightsStore2[109];
			WeightsStore2[26] <= WeightsStore2[110];
			WeightsStore2[27] <= WeightsStore2[111];
			WeightsStore3[0] <= WeightsStore3[84];
			WeightsStore3[1] <= WeightsStore3[85];
			WeightsStore3[2] <= WeightsStore3[86];
			WeightsStore3[3] <= WeightsStore3[87];
			WeightsStore3[4] <= WeightsStore3[88];
			WeightsStore3[5] <= WeightsStore3[89];
			WeightsStore3[6] <= WeightsStore3[90];
			WeightsStore3[7] <= WeightsStore3[91];
			WeightsStore3[8] <= WeightsStore3[92];
			WeightsStore3[9] <= WeightsStore3[93];
			WeightsStore3[10] <= WeightsStore3[94];
			WeightsStore3[11] <= WeightsStore3[95];
			WeightsStore3[12] <= WeightsStore3[96];
			WeightsStore3[13] <= WeightsStore3[97];
			WeightsStore3[14] <= WeightsStore3[98];
			WeightsStore3[15] <= WeightsStore3[99];
			WeightsStore3[16] <= WeightsStore3[100];
			WeightsStore3[17] <= WeightsStore3[101];
			WeightsStore3[18] <= WeightsStore3[102];
			WeightsStore3[19] <= WeightsStore3[103];
			WeightsStore3[20] <= WeightsStore3[104];
			WeightsStore3[21] <= WeightsStore3[105];
			WeightsStore3[22] <= WeightsStore3[106];
			WeightsStore3[23] <= WeightsStore3[107];
			WeightsStore3[24] <= WeightsStore3[108];
			WeightsStore3[25] <= WeightsStore3[109];
			WeightsStore3[26] <= WeightsStore3[110];
			WeightsStore3[27] <= WeightsStore3[111];
			WeightsStore4[0] <= WeightsStore4[84];
			WeightsStore4[1] <= WeightsStore4[85];
			WeightsStore4[2] <= WeightsStore4[86];
			WeightsStore4[3] <= WeightsStore4[87];
			WeightsStore4[4] <= WeightsStore4[88];
			WeightsStore4[5] <= WeightsStore4[89];
			WeightsStore4[6] <= WeightsStore4[90];
			WeightsStore4[7] <= WeightsStore4[91];
			WeightsStore4[8] <= WeightsStore4[92];
			WeightsStore4[9] <= WeightsStore4[93];
			WeightsStore4[10] <= WeightsStore4[94];
			WeightsStore4[11] <= WeightsStore4[95];
			WeightsStore4[12] <= WeightsStore4[96];
			WeightsStore4[13] <= WeightsStore4[97];
			WeightsStore4[14] <= WeightsStore4[98];
			WeightsStore4[15] <= WeightsStore4[99];
			WeightsStore4[16] <= WeightsStore4[100];
			WeightsStore4[17] <= WeightsStore4[101];
			WeightsStore4[18] <= WeightsStore4[102];
			WeightsStore4[19] <= WeightsStore4[103];
			WeightsStore4[20] <= WeightsStore4[104];
			WeightsStore4[21] <= WeightsStore4[105];
			WeightsStore4[22] <= WeightsStore4[106];
			WeightsStore4[23] <= WeightsStore4[107];
			WeightsStore4[24] <= WeightsStore4[108];
			WeightsStore4[25] <= WeightsStore4[109];
			WeightsStore4[26] <= WeightsStore4[110];
			WeightsStore4[27] <= WeightsStore4[111];
			WeightsStore5[0] <= WeightsStore5[84];
			WeightsStore5[1] <= WeightsStore5[85];
			WeightsStore5[2] <= WeightsStore5[86];
			WeightsStore5[3] <= WeightsStore5[87];
			WeightsStore5[4] <= WeightsStore5[88];
			WeightsStore5[5] <= WeightsStore5[89];
			WeightsStore5[6] <= WeightsStore5[90];
			WeightsStore5[7] <= WeightsStore5[91];
			WeightsStore5[8] <= WeightsStore5[92];
			WeightsStore5[9] <= WeightsStore5[93];
			WeightsStore5[10] <= WeightsStore5[94];
			WeightsStore5[11] <= WeightsStore5[95];
			WeightsStore5[12] <= WeightsStore5[96];
			WeightsStore5[13] <= WeightsStore5[97];
			WeightsStore5[14] <= WeightsStore5[98];
			WeightsStore5[15] <= WeightsStore5[99];
			WeightsStore5[16] <= WeightsStore5[100];
			WeightsStore5[17] <= WeightsStore5[101];
			WeightsStore5[18] <= WeightsStore5[102];
			WeightsStore5[19] <= WeightsStore5[103];
			WeightsStore5[20] <= WeightsStore5[104];
			WeightsStore5[21] <= WeightsStore5[105];
			WeightsStore5[22] <= WeightsStore5[106];
			WeightsStore5[23] <= WeightsStore5[107];
			WeightsStore5[24] <= WeightsStore5[108];
			WeightsStore5[25] <= WeightsStore5[109];
			WeightsStore5[26] <= WeightsStore5[110];
			WeightsStore5[27] <= WeightsStore5[111];
			WeightsStore6[0] <= WeightsStore6[84];
			WeightsStore6[1] <= WeightsStore6[85];
			WeightsStore6[2] <= WeightsStore6[86];
			WeightsStore6[3] <= WeightsStore6[87];
			WeightsStore6[4] <= WeightsStore6[88];
			WeightsStore6[5] <= WeightsStore6[89];
			WeightsStore6[6] <= WeightsStore6[90];
			WeightsStore6[7] <= WeightsStore6[91];
			WeightsStore6[8] <= WeightsStore6[92];
			WeightsStore6[9] <= WeightsStore6[93];
			WeightsStore6[10] <= WeightsStore6[94];
			WeightsStore6[11] <= WeightsStore6[95];
			WeightsStore6[12] <= WeightsStore6[96];
			WeightsStore6[13] <= WeightsStore6[97];
			WeightsStore6[14] <= WeightsStore6[98];
			WeightsStore6[15] <= WeightsStore6[99];
			WeightsStore6[16] <= WeightsStore6[100];
			WeightsStore6[17] <= WeightsStore6[101];
			WeightsStore6[18] <= WeightsStore6[102];
			WeightsStore6[19] <= WeightsStore6[103];
			WeightsStore6[20] <= WeightsStore6[104];
			WeightsStore6[21] <= WeightsStore6[105];
			WeightsStore6[22] <= WeightsStore6[106];
			WeightsStore6[23] <= WeightsStore6[107];
			WeightsStore6[24] <= WeightsStore6[108];
			WeightsStore6[25] <= WeightsStore6[109];
			WeightsStore6[26] <= WeightsStore6[110];
			WeightsStore6[27] <= WeightsStore6[111];
			WeightsStore7[0] <= WeightsStore7[84];
			WeightsStore7[1] <= WeightsStore7[85];
			WeightsStore7[2] <= WeightsStore7[86];
			WeightsStore7[3] <= WeightsStore7[87];
			WeightsStore7[4] <= WeightsStore7[88];
			WeightsStore7[5] <= WeightsStore7[89];
			WeightsStore7[6] <= WeightsStore7[90];
			WeightsStore7[7] <= WeightsStore7[91];
			WeightsStore7[8] <= WeightsStore7[92];
			WeightsStore7[9] <= WeightsStore7[93];
			WeightsStore7[10] <= WeightsStore7[94];
			WeightsStore7[11] <= WeightsStore7[95];
			WeightsStore7[12] <= WeightsStore7[96];
			WeightsStore7[13] <= WeightsStore7[97];
			WeightsStore7[14] <= WeightsStore7[98];
			WeightsStore7[15] <= WeightsStore7[99];
			WeightsStore7[16] <= WeightsStore7[100];
			WeightsStore7[17] <= WeightsStore7[101];
			WeightsStore7[18] <= WeightsStore7[102];
			WeightsStore7[19] <= WeightsStore7[103];
			WeightsStore7[20] <= WeightsStore7[104];
			WeightsStore7[21] <= WeightsStore7[105];
			WeightsStore7[22] <= WeightsStore7[106];
			WeightsStore7[23] <= WeightsStore7[107];
			WeightsStore7[24] <= WeightsStore7[108];
			WeightsStore7[25] <= WeightsStore7[109];
			WeightsStore7[26] <= WeightsStore7[110];
			WeightsStore7[27] <= WeightsStore7[111];
			WeightsStore8[0] <= WeightsStore8[84];
			WeightsStore8[1] <= WeightsStore8[85];
			WeightsStore8[2] <= WeightsStore8[86];
			WeightsStore8[3] <= WeightsStore8[87];
			WeightsStore8[4] <= WeightsStore8[88];
			WeightsStore8[5] <= WeightsStore8[89];
			WeightsStore8[6] <= WeightsStore8[90];
			WeightsStore8[7] <= WeightsStore8[91];
			WeightsStore8[8] <= WeightsStore8[92];
			WeightsStore8[9] <= WeightsStore8[93];
			WeightsStore8[10] <= WeightsStore8[94];
			WeightsStore8[11] <= WeightsStore8[95];
			WeightsStore8[12] <= WeightsStore8[96];
			WeightsStore8[13] <= WeightsStore8[97];
			WeightsStore8[14] <= WeightsStore8[98];
			WeightsStore8[15] <= WeightsStore8[99];
			WeightsStore8[16] <= WeightsStore8[100];
			WeightsStore8[17] <= WeightsStore8[101];
			WeightsStore8[18] <= WeightsStore8[102];
			WeightsStore8[19] <= WeightsStore8[103];
			WeightsStore8[20] <= WeightsStore8[104];
			WeightsStore8[21] <= WeightsStore8[105];
			WeightsStore8[22] <= WeightsStore8[106];
			WeightsStore8[23] <= WeightsStore8[107];
			WeightsStore8[24] <= WeightsStore8[108];
			WeightsStore8[25] <= WeightsStore8[109];
			WeightsStore8[26] <= WeightsStore8[110];
			WeightsStore8[27] <= WeightsStore8[111];
			WeightsStore9[0] <= WeightsStore9[84];
			WeightsStore9[1] <= WeightsStore9[85];
			WeightsStore9[2] <= WeightsStore9[86];
			WeightsStore9[3] <= WeightsStore9[87];
			WeightsStore9[4] <= WeightsStore9[88];
			WeightsStore9[5] <= WeightsStore9[89];
			WeightsStore9[6] <= WeightsStore9[90];
			WeightsStore9[7] <= WeightsStore9[91];
			WeightsStore9[8] <= WeightsStore9[92];
			WeightsStore9[9] <= WeightsStore9[93];
			WeightsStore9[10] <= WeightsStore9[94];
			WeightsStore9[11] <= WeightsStore9[95];
			WeightsStore9[12] <= WeightsStore9[96];
			WeightsStore9[13] <= WeightsStore9[97];
			WeightsStore9[14] <= WeightsStore9[98];
			WeightsStore9[15] <= WeightsStore9[99];
			WeightsStore9[16] <= WeightsStore9[100];
			WeightsStore9[17] <= WeightsStore9[101];
			WeightsStore9[18] <= WeightsStore9[102];
			WeightsStore9[19] <= WeightsStore9[103];
			WeightsStore9[20] <= WeightsStore9[104];
			WeightsStore9[21] <= WeightsStore9[105];
			WeightsStore9[22] <= WeightsStore9[106];
			WeightsStore9[23] <= WeightsStore9[107];
			WeightsStore9[24] <= WeightsStore9[108];
			WeightsStore9[25] <= WeightsStore9[109];
			WeightsStore9[26] <= WeightsStore9[110];
			WeightsStore9[27] <= WeightsStore9[111];
		end else if(switchCounter == 32'd27)begin
			PixelsStore[0] <= PixelsStore[112];
			PixelsStore[1] <= PixelsStore[113];
			PixelsStore[2] <= PixelsStore[114];
			PixelsStore[3] <= PixelsStore[115];
			PixelsStore[4] <= PixelsStore[116];
			PixelsStore[5] <= PixelsStore[117];
			PixelsStore[6] <= PixelsStore[118];
			PixelsStore[7] <= PixelsStore[119];
			PixelsStore[8] <= PixelsStore[120];
			PixelsStore[9] <= PixelsStore[121];
			PixelsStore[10] <= PixelsStore[122];
			PixelsStore[11] <= PixelsStore[123];
			PixelsStore[12] <= PixelsStore[124];
			PixelsStore[13] <= PixelsStore[125];
			PixelsStore[14] <= PixelsStore[126];
			PixelsStore[15] <= PixelsStore[127];
			PixelsStore[16] <= PixelsStore[128];
			PixelsStore[17] <= PixelsStore[129];
			PixelsStore[18] <= PixelsStore[130];
			PixelsStore[19] <= PixelsStore[131];
			PixelsStore[20] <= PixelsStore[132];
			PixelsStore[21] <= PixelsStore[133];
			PixelsStore[22] <= PixelsStore[134];
			PixelsStore[23] <= PixelsStore[135];
			PixelsStore[24] <= PixelsStore[136];
			PixelsStore[25] <= PixelsStore[137];
			PixelsStore[26] <= PixelsStore[138];
			PixelsStore[27] <= PixelsStore[139];
			WeightsStore0[0] <= WeightsStore0[112];
			WeightsStore0[1] <= WeightsStore0[113];
			WeightsStore0[2] <= WeightsStore0[114];
			WeightsStore0[3] <= WeightsStore0[115];
			WeightsStore0[4] <= WeightsStore0[116];
			WeightsStore0[5] <= WeightsStore0[117];
			WeightsStore0[6] <= WeightsStore0[118];
			WeightsStore0[7] <= WeightsStore0[119];
			WeightsStore0[8] <= WeightsStore0[120];
			WeightsStore0[9] <= WeightsStore0[121];
			WeightsStore0[10] <= WeightsStore0[122];
			WeightsStore0[11] <= WeightsStore0[123];
			WeightsStore0[12] <= WeightsStore0[124];
			WeightsStore0[13] <= WeightsStore0[125];
			WeightsStore0[14] <= WeightsStore0[126];
			WeightsStore0[15] <= WeightsStore0[127];
			WeightsStore0[16] <= WeightsStore0[128];
			WeightsStore0[17] <= WeightsStore0[129];
			WeightsStore0[18] <= WeightsStore0[130];
			WeightsStore0[19] <= WeightsStore0[131];
			WeightsStore0[20] <= WeightsStore0[132];
			WeightsStore0[21] <= WeightsStore0[133];
			WeightsStore0[22] <= WeightsStore0[134];
			WeightsStore0[23] <= WeightsStore0[135];
			WeightsStore0[24] <= WeightsStore0[136];
			WeightsStore0[25] <= WeightsStore0[137];
			WeightsStore0[26] <= WeightsStore0[138];
			WeightsStore0[27] <= WeightsStore0[139];
			WeightsStore1[0] <= WeightsStore1[112];
			WeightsStore1[1] <= WeightsStore1[113];
			WeightsStore1[2] <= WeightsStore1[114];
			WeightsStore1[3] <= WeightsStore1[115];
			WeightsStore1[4] <= WeightsStore1[116];
			WeightsStore1[5] <= WeightsStore1[117];
			WeightsStore1[6] <= WeightsStore1[118];
			WeightsStore1[7] <= WeightsStore1[119];
			WeightsStore1[8] <= WeightsStore1[120];
			WeightsStore1[9] <= WeightsStore1[121];
			WeightsStore1[10] <= WeightsStore1[122];
			WeightsStore1[11] <= WeightsStore1[123];
			WeightsStore1[12] <= WeightsStore1[124];
			WeightsStore1[13] <= WeightsStore1[125];
			WeightsStore1[14] <= WeightsStore1[126];
			WeightsStore1[15] <= WeightsStore1[127];
			WeightsStore1[16] <= WeightsStore1[128];
			WeightsStore1[17] <= WeightsStore1[129];
			WeightsStore1[18] <= WeightsStore1[130];
			WeightsStore1[19] <= WeightsStore1[131];
			WeightsStore1[20] <= WeightsStore1[132];
			WeightsStore1[21] <= WeightsStore1[133];
			WeightsStore1[22] <= WeightsStore1[134];
			WeightsStore1[23] <= WeightsStore1[135];
			WeightsStore1[24] <= WeightsStore1[136];
			WeightsStore1[25] <= WeightsStore1[137];
			WeightsStore1[26] <= WeightsStore1[138];
			WeightsStore1[27] <= WeightsStore1[139];
			WeightsStore2[0] <= WeightsStore2[112];
			WeightsStore2[1] <= WeightsStore2[113];
			WeightsStore2[2] <= WeightsStore2[114];
			WeightsStore2[3] <= WeightsStore2[115];
			WeightsStore2[4] <= WeightsStore2[116];
			WeightsStore2[5] <= WeightsStore2[117];
			WeightsStore2[6] <= WeightsStore2[118];
			WeightsStore2[7] <= WeightsStore2[119];
			WeightsStore2[8] <= WeightsStore2[120];
			WeightsStore2[9] <= WeightsStore2[121];
			WeightsStore2[10] <= WeightsStore2[122];
			WeightsStore2[11] <= WeightsStore2[123];
			WeightsStore2[12] <= WeightsStore2[124];
			WeightsStore2[13] <= WeightsStore2[125];
			WeightsStore2[14] <= WeightsStore2[126];
			WeightsStore2[15] <= WeightsStore2[127];
			WeightsStore2[16] <= WeightsStore2[128];
			WeightsStore2[17] <= WeightsStore2[129];
			WeightsStore2[18] <= WeightsStore2[130];
			WeightsStore2[19] <= WeightsStore2[131];
			WeightsStore2[20] <= WeightsStore2[132];
			WeightsStore2[21] <= WeightsStore2[133];
			WeightsStore2[22] <= WeightsStore2[134];
			WeightsStore2[23] <= WeightsStore2[135];
			WeightsStore2[24] <= WeightsStore2[136];
			WeightsStore2[25] <= WeightsStore2[137];
			WeightsStore2[26] <= WeightsStore2[138];
			WeightsStore2[27] <= WeightsStore2[139];
			WeightsStore3[0] <= WeightsStore3[112];
			WeightsStore3[1] <= WeightsStore3[113];
			WeightsStore3[2] <= WeightsStore3[114];
			WeightsStore3[3] <= WeightsStore3[115];
			WeightsStore3[4] <= WeightsStore3[116];
			WeightsStore3[5] <= WeightsStore3[117];
			WeightsStore3[6] <= WeightsStore3[118];
			WeightsStore3[7] <= WeightsStore3[119];
			WeightsStore3[8] <= WeightsStore3[120];
			WeightsStore3[9] <= WeightsStore3[121];
			WeightsStore3[10] <= WeightsStore3[122];
			WeightsStore3[11] <= WeightsStore3[123];
			WeightsStore3[12] <= WeightsStore3[124];
			WeightsStore3[13] <= WeightsStore3[125];
			WeightsStore3[14] <= WeightsStore3[126];
			WeightsStore3[15] <= WeightsStore3[127];
			WeightsStore3[16] <= WeightsStore3[128];
			WeightsStore3[17] <= WeightsStore3[129];
			WeightsStore3[18] <= WeightsStore3[130];
			WeightsStore3[19] <= WeightsStore3[131];
			WeightsStore3[20] <= WeightsStore3[132];
			WeightsStore3[21] <= WeightsStore3[133];
			WeightsStore3[22] <= WeightsStore3[134];
			WeightsStore3[23] <= WeightsStore3[135];
			WeightsStore3[24] <= WeightsStore3[136];
			WeightsStore3[25] <= WeightsStore3[137];
			WeightsStore3[26] <= WeightsStore3[138];
			WeightsStore3[27] <= WeightsStore3[139];
			WeightsStore4[0] <= WeightsStore4[112];
			WeightsStore4[1] <= WeightsStore4[113];
			WeightsStore4[2] <= WeightsStore4[114];
			WeightsStore4[3] <= WeightsStore4[115];
			WeightsStore4[4] <= WeightsStore4[116];
			WeightsStore4[5] <= WeightsStore4[117];
			WeightsStore4[6] <= WeightsStore4[118];
			WeightsStore4[7] <= WeightsStore4[119];
			WeightsStore4[8] <= WeightsStore4[120];
			WeightsStore4[9] <= WeightsStore4[121];
			WeightsStore4[10] <= WeightsStore4[122];
			WeightsStore4[11] <= WeightsStore4[123];
			WeightsStore4[12] <= WeightsStore4[124];
			WeightsStore4[13] <= WeightsStore4[125];
			WeightsStore4[14] <= WeightsStore4[126];
			WeightsStore4[15] <= WeightsStore4[127];
			WeightsStore4[16] <= WeightsStore4[128];
			WeightsStore4[17] <= WeightsStore4[129];
			WeightsStore4[18] <= WeightsStore4[130];
			WeightsStore4[19] <= WeightsStore4[131];
			WeightsStore4[20] <= WeightsStore4[132];
			WeightsStore4[21] <= WeightsStore4[133];
			WeightsStore4[22] <= WeightsStore4[134];
			WeightsStore4[23] <= WeightsStore4[135];
			WeightsStore4[24] <= WeightsStore4[136];
			WeightsStore4[25] <= WeightsStore4[137];
			WeightsStore4[26] <= WeightsStore4[138];
			WeightsStore4[27] <= WeightsStore4[139];
			WeightsStore5[0] <= WeightsStore5[112];
			WeightsStore5[1] <= WeightsStore5[113];
			WeightsStore5[2] <= WeightsStore5[114];
			WeightsStore5[3] <= WeightsStore5[115];
			WeightsStore5[4] <= WeightsStore5[116];
			WeightsStore5[5] <= WeightsStore5[117];
			WeightsStore5[6] <= WeightsStore5[118];
			WeightsStore5[7] <= WeightsStore5[119];
			WeightsStore5[8] <= WeightsStore5[120];
			WeightsStore5[9] <= WeightsStore5[121];
			WeightsStore5[10] <= WeightsStore5[122];
			WeightsStore5[11] <= WeightsStore5[123];
			WeightsStore5[12] <= WeightsStore5[124];
			WeightsStore5[13] <= WeightsStore5[125];
			WeightsStore5[14] <= WeightsStore5[126];
			WeightsStore5[15] <= WeightsStore5[127];
			WeightsStore5[16] <= WeightsStore5[128];
			WeightsStore5[17] <= WeightsStore5[129];
			WeightsStore5[18] <= WeightsStore5[130];
			WeightsStore5[19] <= WeightsStore5[131];
			WeightsStore5[20] <= WeightsStore5[132];
			WeightsStore5[21] <= WeightsStore5[133];
			WeightsStore5[22] <= WeightsStore5[134];
			WeightsStore5[23] <= WeightsStore5[135];
			WeightsStore5[24] <= WeightsStore5[136];
			WeightsStore5[25] <= WeightsStore5[137];
			WeightsStore5[26] <= WeightsStore5[138];
			WeightsStore5[27] <= WeightsStore5[139];
			WeightsStore6[0] <= WeightsStore6[112];
			WeightsStore6[1] <= WeightsStore6[113];
			WeightsStore6[2] <= WeightsStore6[114];
			WeightsStore6[3] <= WeightsStore6[115];
			WeightsStore6[4] <= WeightsStore6[116];
			WeightsStore6[5] <= WeightsStore6[117];
			WeightsStore6[6] <= WeightsStore6[118];
			WeightsStore6[7] <= WeightsStore6[119];
			WeightsStore6[8] <= WeightsStore6[120];
			WeightsStore6[9] <= WeightsStore6[121];
			WeightsStore6[10] <= WeightsStore6[122];
			WeightsStore6[11] <= WeightsStore6[123];
			WeightsStore6[12] <= WeightsStore6[124];
			WeightsStore6[13] <= WeightsStore6[125];
			WeightsStore6[14] <= WeightsStore6[126];
			WeightsStore6[15] <= WeightsStore6[127];
			WeightsStore6[16] <= WeightsStore6[128];
			WeightsStore6[17] <= WeightsStore6[129];
			WeightsStore6[18] <= WeightsStore6[130];
			WeightsStore6[19] <= WeightsStore6[131];
			WeightsStore6[20] <= WeightsStore6[132];
			WeightsStore6[21] <= WeightsStore6[133];
			WeightsStore6[22] <= WeightsStore6[134];
			WeightsStore6[23] <= WeightsStore6[135];
			WeightsStore6[24] <= WeightsStore6[136];
			WeightsStore6[25] <= WeightsStore6[137];
			WeightsStore6[26] <= WeightsStore6[138];
			WeightsStore6[27] <= WeightsStore6[139];
			WeightsStore7[0] <= WeightsStore7[112];
			WeightsStore7[1] <= WeightsStore7[113];
			WeightsStore7[2] <= WeightsStore7[114];
			WeightsStore7[3] <= WeightsStore7[115];
			WeightsStore7[4] <= WeightsStore7[116];
			WeightsStore7[5] <= WeightsStore7[117];
			WeightsStore7[6] <= WeightsStore7[118];
			WeightsStore7[7] <= WeightsStore7[119];
			WeightsStore7[8] <= WeightsStore7[120];
			WeightsStore7[9] <= WeightsStore7[121];
			WeightsStore7[10] <= WeightsStore7[122];
			WeightsStore7[11] <= WeightsStore7[123];
			WeightsStore7[12] <= WeightsStore7[124];
			WeightsStore7[13] <= WeightsStore7[125];
			WeightsStore7[14] <= WeightsStore7[126];
			WeightsStore7[15] <= WeightsStore7[127];
			WeightsStore7[16] <= WeightsStore7[128];
			WeightsStore7[17] <= WeightsStore7[129];
			WeightsStore7[18] <= WeightsStore7[130];
			WeightsStore7[19] <= WeightsStore7[131];
			WeightsStore7[20] <= WeightsStore7[132];
			WeightsStore7[21] <= WeightsStore7[133];
			WeightsStore7[22] <= WeightsStore7[134];
			WeightsStore7[23] <= WeightsStore7[135];
			WeightsStore7[24] <= WeightsStore7[136];
			WeightsStore7[25] <= WeightsStore7[137];
			WeightsStore7[26] <= WeightsStore7[138];
			WeightsStore7[27] <= WeightsStore7[139];
			WeightsStore8[0] <= WeightsStore8[112];
			WeightsStore8[1] <= WeightsStore8[113];
			WeightsStore8[2] <= WeightsStore8[114];
			WeightsStore8[3] <= WeightsStore8[115];
			WeightsStore8[4] <= WeightsStore8[116];
			WeightsStore8[5] <= WeightsStore8[117];
			WeightsStore8[6] <= WeightsStore8[118];
			WeightsStore8[7] <= WeightsStore8[119];
			WeightsStore8[8] <= WeightsStore8[120];
			WeightsStore8[9] <= WeightsStore8[121];
			WeightsStore8[10] <= WeightsStore8[122];
			WeightsStore8[11] <= WeightsStore8[123];
			WeightsStore8[12] <= WeightsStore8[124];
			WeightsStore8[13] <= WeightsStore8[125];
			WeightsStore8[14] <= WeightsStore8[126];
			WeightsStore8[15] <= WeightsStore8[127];
			WeightsStore8[16] <= WeightsStore8[128];
			WeightsStore8[17] <= WeightsStore8[129];
			WeightsStore8[18] <= WeightsStore8[130];
			WeightsStore8[19] <= WeightsStore8[131];
			WeightsStore8[20] <= WeightsStore8[132];
			WeightsStore8[21] <= WeightsStore8[133];
			WeightsStore8[22] <= WeightsStore8[134];
			WeightsStore8[23] <= WeightsStore8[135];
			WeightsStore8[24] <= WeightsStore8[136];
			WeightsStore8[25] <= WeightsStore8[137];
			WeightsStore8[26] <= WeightsStore8[138];
			WeightsStore8[27] <= WeightsStore8[139];
			WeightsStore9[0] <= WeightsStore9[112];
			WeightsStore9[1] <= WeightsStore9[113];
			WeightsStore9[2] <= WeightsStore9[114];
			WeightsStore9[3] <= WeightsStore9[115];
			WeightsStore9[4] <= WeightsStore9[116];
			WeightsStore9[5] <= WeightsStore9[117];
			WeightsStore9[6] <= WeightsStore9[118];
			WeightsStore9[7] <= WeightsStore9[119];
			WeightsStore9[8] <= WeightsStore9[120];
			WeightsStore9[9] <= WeightsStore9[121];
			WeightsStore9[10] <= WeightsStore9[122];
			WeightsStore9[11] <= WeightsStore9[123];
			WeightsStore9[12] <= WeightsStore9[124];
			WeightsStore9[13] <= WeightsStore9[125];
			WeightsStore9[14] <= WeightsStore9[126];
			WeightsStore9[15] <= WeightsStore9[127];
			WeightsStore9[16] <= WeightsStore9[128];
			WeightsStore9[17] <= WeightsStore9[129];
			WeightsStore9[18] <= WeightsStore9[130];
			WeightsStore9[19] <= WeightsStore9[131];
			WeightsStore9[20] <= WeightsStore9[132];
			WeightsStore9[21] <= WeightsStore9[133];
			WeightsStore9[22] <= WeightsStore9[134];
			WeightsStore9[23] <= WeightsStore9[135];
			WeightsStore9[24] <= WeightsStore9[136];
			WeightsStore9[25] <= WeightsStore9[137];
			WeightsStore9[26] <= WeightsStore9[138];
			WeightsStore9[27] <= WeightsStore9[139];
		end else if(switchCounter == 32'd34)begin
			PixelsStore[0] <= PixelsStore[140];
			PixelsStore[1] <= PixelsStore[141];
			PixelsStore[2] <= PixelsStore[142];
			PixelsStore[3] <= PixelsStore[143];
			PixelsStore[4] <= PixelsStore[144];
			PixelsStore[5] <= PixelsStore[145];
			PixelsStore[6] <= PixelsStore[146];
			PixelsStore[7] <= PixelsStore[147];
			PixelsStore[8] <= PixelsStore[148];
			PixelsStore[9] <= PixelsStore[149];
			PixelsStore[10] <= PixelsStore[150];
			PixelsStore[11] <= PixelsStore[151];
			PixelsStore[12] <= PixelsStore[152];
			PixelsStore[13] <= PixelsStore[153];
			PixelsStore[14] <= PixelsStore[154];
			PixelsStore[15] <= PixelsStore[155];
			PixelsStore[16] <= PixelsStore[156];
			PixelsStore[17] <= PixelsStore[157];
			PixelsStore[18] <= PixelsStore[158];
			PixelsStore[19] <= PixelsStore[159];
			PixelsStore[20] <= PixelsStore[160];
			PixelsStore[21] <= PixelsStore[161];
			PixelsStore[22] <= PixelsStore[162];
			PixelsStore[23] <= PixelsStore[163];
			PixelsStore[24] <= PixelsStore[164];
			PixelsStore[25] <= PixelsStore[165];
			PixelsStore[26] <= PixelsStore[166];
			PixelsStore[27] <= PixelsStore[167];
			WeightsStore0[0] <= WeightsStore0[140];
			WeightsStore0[1] <= WeightsStore0[141];
			WeightsStore0[2] <= WeightsStore0[142];
			WeightsStore0[3] <= WeightsStore0[143];
			WeightsStore0[4] <= WeightsStore0[144];
			WeightsStore0[5] <= WeightsStore0[145];
			WeightsStore0[6] <= WeightsStore0[146];
			WeightsStore0[7] <= WeightsStore0[147];
			WeightsStore0[8] <= WeightsStore0[148];
			WeightsStore0[9] <= WeightsStore0[149];
			WeightsStore0[10] <= WeightsStore0[150];
			WeightsStore0[11] <= WeightsStore0[151];
			WeightsStore0[12] <= WeightsStore0[152];
			WeightsStore0[13] <= WeightsStore0[153];
			WeightsStore0[14] <= WeightsStore0[154];
			WeightsStore0[15] <= WeightsStore0[155];
			WeightsStore0[16] <= WeightsStore0[156];
			WeightsStore0[17] <= WeightsStore0[157];
			WeightsStore0[18] <= WeightsStore0[158];
			WeightsStore0[19] <= WeightsStore0[159];
			WeightsStore0[20] <= WeightsStore0[160];
			WeightsStore0[21] <= WeightsStore0[161];
			WeightsStore0[22] <= WeightsStore0[162];
			WeightsStore0[23] <= WeightsStore0[163];
			WeightsStore0[24] <= WeightsStore0[164];
			WeightsStore0[25] <= WeightsStore0[165];
			WeightsStore0[26] <= WeightsStore0[166];
			WeightsStore0[27] <= WeightsStore0[167];
			WeightsStore1[0] <= WeightsStore1[140];
			WeightsStore1[1] <= WeightsStore1[141];
			WeightsStore1[2] <= WeightsStore1[142];
			WeightsStore1[3] <= WeightsStore1[143];
			WeightsStore1[4] <= WeightsStore1[144];
			WeightsStore1[5] <= WeightsStore1[145];
			WeightsStore1[6] <= WeightsStore1[146];
			WeightsStore1[7] <= WeightsStore1[147];
			WeightsStore1[8] <= WeightsStore1[148];
			WeightsStore1[9] <= WeightsStore1[149];
			WeightsStore1[10] <= WeightsStore1[150];
			WeightsStore1[11] <= WeightsStore1[151];
			WeightsStore1[12] <= WeightsStore1[152];
			WeightsStore1[13] <= WeightsStore1[153];
			WeightsStore1[14] <= WeightsStore1[154];
			WeightsStore1[15] <= WeightsStore1[155];
			WeightsStore1[16] <= WeightsStore1[156];
			WeightsStore1[17] <= WeightsStore1[157];
			WeightsStore1[18] <= WeightsStore1[158];
			WeightsStore1[19] <= WeightsStore1[159];
			WeightsStore1[20] <= WeightsStore1[160];
			WeightsStore1[21] <= WeightsStore1[161];
			WeightsStore1[22] <= WeightsStore1[162];
			WeightsStore1[23] <= WeightsStore1[163];
			WeightsStore1[24] <= WeightsStore1[164];
			WeightsStore1[25] <= WeightsStore1[165];
			WeightsStore1[26] <= WeightsStore1[166];
			WeightsStore1[27] <= WeightsStore1[167];
			WeightsStore2[0] <= WeightsStore2[140];
			WeightsStore2[1] <= WeightsStore2[141];
			WeightsStore2[2] <= WeightsStore2[142];
			WeightsStore2[3] <= WeightsStore2[143];
			WeightsStore2[4] <= WeightsStore2[144];
			WeightsStore2[5] <= WeightsStore2[145];
			WeightsStore2[6] <= WeightsStore2[146];
			WeightsStore2[7] <= WeightsStore2[147];
			WeightsStore2[8] <= WeightsStore2[148];
			WeightsStore2[9] <= WeightsStore2[149];
			WeightsStore2[10] <= WeightsStore2[150];
			WeightsStore2[11] <= WeightsStore2[151];
			WeightsStore2[12] <= WeightsStore2[152];
			WeightsStore2[13] <= WeightsStore2[153];
			WeightsStore2[14] <= WeightsStore2[154];
			WeightsStore2[15] <= WeightsStore2[155];
			WeightsStore2[16] <= WeightsStore2[156];
			WeightsStore2[17] <= WeightsStore2[157];
			WeightsStore2[18] <= WeightsStore2[158];
			WeightsStore2[19] <= WeightsStore2[159];
			WeightsStore2[20] <= WeightsStore2[160];
			WeightsStore2[21] <= WeightsStore2[161];
			WeightsStore2[22] <= WeightsStore2[162];
			WeightsStore2[23] <= WeightsStore2[163];
			WeightsStore2[24] <= WeightsStore2[164];
			WeightsStore2[25] <= WeightsStore2[165];
			WeightsStore2[26] <= WeightsStore2[166];
			WeightsStore2[27] <= WeightsStore2[167];
			WeightsStore3[0] <= WeightsStore3[140];
			WeightsStore3[1] <= WeightsStore3[141];
			WeightsStore3[2] <= WeightsStore3[142];
			WeightsStore3[3] <= WeightsStore3[143];
			WeightsStore3[4] <= WeightsStore3[144];
			WeightsStore3[5] <= WeightsStore3[145];
			WeightsStore3[6] <= WeightsStore3[146];
			WeightsStore3[7] <= WeightsStore3[147];
			WeightsStore3[8] <= WeightsStore3[148];
			WeightsStore3[9] <= WeightsStore3[149];
			WeightsStore3[10] <= WeightsStore3[150];
			WeightsStore3[11] <= WeightsStore3[151];
			WeightsStore3[12] <= WeightsStore3[152];
			WeightsStore3[13] <= WeightsStore3[153];
			WeightsStore3[14] <= WeightsStore3[154];
			WeightsStore3[15] <= WeightsStore3[155];
			WeightsStore3[16] <= WeightsStore3[156];
			WeightsStore3[17] <= WeightsStore3[157];
			WeightsStore3[18] <= WeightsStore3[158];
			WeightsStore3[19] <= WeightsStore3[159];
			WeightsStore3[20] <= WeightsStore3[160];
			WeightsStore3[21] <= WeightsStore3[161];
			WeightsStore3[22] <= WeightsStore3[162];
			WeightsStore3[23] <= WeightsStore3[163];
			WeightsStore3[24] <= WeightsStore3[164];
			WeightsStore3[25] <= WeightsStore3[165];
			WeightsStore3[26] <= WeightsStore3[166];
			WeightsStore3[27] <= WeightsStore3[167];
			WeightsStore4[0] <= WeightsStore4[140];
			WeightsStore4[1] <= WeightsStore4[141];
			WeightsStore4[2] <= WeightsStore4[142];
			WeightsStore4[3] <= WeightsStore4[143];
			WeightsStore4[4] <= WeightsStore4[144];
			WeightsStore4[5] <= WeightsStore4[145];
			WeightsStore4[6] <= WeightsStore4[146];
			WeightsStore4[7] <= WeightsStore4[147];
			WeightsStore4[8] <= WeightsStore4[148];
			WeightsStore4[9] <= WeightsStore4[149];
			WeightsStore4[10] <= WeightsStore4[150];
			WeightsStore4[11] <= WeightsStore4[151];
			WeightsStore4[12] <= WeightsStore4[152];
			WeightsStore4[13] <= WeightsStore4[153];
			WeightsStore4[14] <= WeightsStore4[154];
			WeightsStore4[15] <= WeightsStore4[155];
			WeightsStore4[16] <= WeightsStore4[156];
			WeightsStore4[17] <= WeightsStore4[157];
			WeightsStore4[18] <= WeightsStore4[158];
			WeightsStore4[19] <= WeightsStore4[159];
			WeightsStore4[20] <= WeightsStore4[160];
			WeightsStore4[21] <= WeightsStore4[161];
			WeightsStore4[22] <= WeightsStore4[162];
			WeightsStore4[23] <= WeightsStore4[163];
			WeightsStore4[24] <= WeightsStore4[164];
			WeightsStore4[25] <= WeightsStore4[165];
			WeightsStore4[26] <= WeightsStore4[166];
			WeightsStore4[27] <= WeightsStore4[167];
			WeightsStore5[0] <= WeightsStore5[140];
			WeightsStore5[1] <= WeightsStore5[141];
			WeightsStore5[2] <= WeightsStore5[142];
			WeightsStore5[3] <= WeightsStore5[143];
			WeightsStore5[4] <= WeightsStore5[144];
			WeightsStore5[5] <= WeightsStore5[145];
			WeightsStore5[6] <= WeightsStore5[146];
			WeightsStore5[7] <= WeightsStore5[147];
			WeightsStore5[8] <= WeightsStore5[148];
			WeightsStore5[9] <= WeightsStore5[149];
			WeightsStore5[10] <= WeightsStore5[150];
			WeightsStore5[11] <= WeightsStore5[151];
			WeightsStore5[12] <= WeightsStore5[152];
			WeightsStore5[13] <= WeightsStore5[153];
			WeightsStore5[14] <= WeightsStore5[154];
			WeightsStore5[15] <= WeightsStore5[155];
			WeightsStore5[16] <= WeightsStore5[156];
			WeightsStore5[17] <= WeightsStore5[157];
			WeightsStore5[18] <= WeightsStore5[158];
			WeightsStore5[19] <= WeightsStore5[159];
			WeightsStore5[20] <= WeightsStore5[160];
			WeightsStore5[21] <= WeightsStore5[161];
			WeightsStore5[22] <= WeightsStore5[162];
			WeightsStore5[23] <= WeightsStore5[163];
			WeightsStore5[24] <= WeightsStore5[164];
			WeightsStore5[25] <= WeightsStore5[165];
			WeightsStore5[26] <= WeightsStore5[166];
			WeightsStore5[27] <= WeightsStore5[167];
			WeightsStore6[0] <= WeightsStore6[140];
			WeightsStore6[1] <= WeightsStore6[141];
			WeightsStore6[2] <= WeightsStore6[142];
			WeightsStore6[3] <= WeightsStore6[143];
			WeightsStore6[4] <= WeightsStore6[144];
			WeightsStore6[5] <= WeightsStore6[145];
			WeightsStore6[6] <= WeightsStore6[146];
			WeightsStore6[7] <= WeightsStore6[147];
			WeightsStore6[8] <= WeightsStore6[148];
			WeightsStore6[9] <= WeightsStore6[149];
			WeightsStore6[10] <= WeightsStore6[150];
			WeightsStore6[11] <= WeightsStore6[151];
			WeightsStore6[12] <= WeightsStore6[152];
			WeightsStore6[13] <= WeightsStore6[153];
			WeightsStore6[14] <= WeightsStore6[154];
			WeightsStore6[15] <= WeightsStore6[155];
			WeightsStore6[16] <= WeightsStore6[156];
			WeightsStore6[17] <= WeightsStore6[157];
			WeightsStore6[18] <= WeightsStore6[158];
			WeightsStore6[19] <= WeightsStore6[159];
			WeightsStore6[20] <= WeightsStore6[160];
			WeightsStore6[21] <= WeightsStore6[161];
			WeightsStore6[22] <= WeightsStore6[162];
			WeightsStore6[23] <= WeightsStore6[163];
			WeightsStore6[24] <= WeightsStore6[164];
			WeightsStore6[25] <= WeightsStore6[165];
			WeightsStore6[26] <= WeightsStore6[166];
			WeightsStore6[27] <= WeightsStore6[167];
			WeightsStore7[0] <= WeightsStore7[140];
			WeightsStore7[1] <= WeightsStore7[141];
			WeightsStore7[2] <= WeightsStore7[142];
			WeightsStore7[3] <= WeightsStore7[143];
			WeightsStore7[4] <= WeightsStore7[144];
			WeightsStore7[5] <= WeightsStore7[145];
			WeightsStore7[6] <= WeightsStore7[146];
			WeightsStore7[7] <= WeightsStore7[147];
			WeightsStore7[8] <= WeightsStore7[148];
			WeightsStore7[9] <= WeightsStore7[149];
			WeightsStore7[10] <= WeightsStore7[150];
			WeightsStore7[11] <= WeightsStore7[151];
			WeightsStore7[12] <= WeightsStore7[152];
			WeightsStore7[13] <= WeightsStore7[153];
			WeightsStore7[14] <= WeightsStore7[154];
			WeightsStore7[15] <= WeightsStore7[155];
			WeightsStore7[16] <= WeightsStore7[156];
			WeightsStore7[17] <= WeightsStore7[157];
			WeightsStore7[18] <= WeightsStore7[158];
			WeightsStore7[19] <= WeightsStore7[159];
			WeightsStore7[20] <= WeightsStore7[160];
			WeightsStore7[21] <= WeightsStore7[161];
			WeightsStore7[22] <= WeightsStore7[162];
			WeightsStore7[23] <= WeightsStore7[163];
			WeightsStore7[24] <= WeightsStore7[164];
			WeightsStore7[25] <= WeightsStore7[165];
			WeightsStore7[26] <= WeightsStore7[166];
			WeightsStore7[27] <= WeightsStore7[167];
			WeightsStore8[0] <= WeightsStore8[140];
			WeightsStore8[1] <= WeightsStore8[141];
			WeightsStore8[2] <= WeightsStore8[142];
			WeightsStore8[3] <= WeightsStore8[143];
			WeightsStore8[4] <= WeightsStore8[144];
			WeightsStore8[5] <= WeightsStore8[145];
			WeightsStore8[6] <= WeightsStore8[146];
			WeightsStore8[7] <= WeightsStore8[147];
			WeightsStore8[8] <= WeightsStore8[148];
			WeightsStore8[9] <= WeightsStore8[149];
			WeightsStore8[10] <= WeightsStore8[150];
			WeightsStore8[11] <= WeightsStore8[151];
			WeightsStore8[12] <= WeightsStore8[152];
			WeightsStore8[13] <= WeightsStore8[153];
			WeightsStore8[14] <= WeightsStore8[154];
			WeightsStore8[15] <= WeightsStore8[155];
			WeightsStore8[16] <= WeightsStore8[156];
			WeightsStore8[17] <= WeightsStore8[157];
			WeightsStore8[18] <= WeightsStore8[158];
			WeightsStore8[19] <= WeightsStore8[159];
			WeightsStore8[20] <= WeightsStore8[160];
			WeightsStore8[21] <= WeightsStore8[161];
			WeightsStore8[22] <= WeightsStore8[162];
			WeightsStore8[23] <= WeightsStore8[163];
			WeightsStore8[24] <= WeightsStore8[164];
			WeightsStore8[25] <= WeightsStore8[165];
			WeightsStore8[26] <= WeightsStore8[166];
			WeightsStore8[27] <= WeightsStore8[167];
			WeightsStore9[0] <= WeightsStore9[140];
			WeightsStore9[1] <= WeightsStore9[141];
			WeightsStore9[2] <= WeightsStore9[142];
			WeightsStore9[3] <= WeightsStore9[143];
			WeightsStore9[4] <= WeightsStore9[144];
			WeightsStore9[5] <= WeightsStore9[145];
			WeightsStore9[6] <= WeightsStore9[146];
			WeightsStore9[7] <= WeightsStore9[147];
			WeightsStore9[8] <= WeightsStore9[148];
			WeightsStore9[9] <= WeightsStore9[149];
			WeightsStore9[10] <= WeightsStore9[150];
			WeightsStore9[11] <= WeightsStore9[151];
			WeightsStore9[12] <= WeightsStore9[152];
			WeightsStore9[13] <= WeightsStore9[153];
			WeightsStore9[14] <= WeightsStore9[154];
			WeightsStore9[15] <= WeightsStore9[155];
			WeightsStore9[16] <= WeightsStore9[156];
			WeightsStore9[17] <= WeightsStore9[157];
			WeightsStore9[18] <= WeightsStore9[158];
			WeightsStore9[19] <= WeightsStore9[159];
			WeightsStore9[20] <= WeightsStore9[160];
			WeightsStore9[21] <= WeightsStore9[161];
			WeightsStore9[22] <= WeightsStore9[162];
			WeightsStore9[23] <= WeightsStore9[163];
			WeightsStore9[24] <= WeightsStore9[164];
			WeightsStore9[25] <= WeightsStore9[165];
			WeightsStore9[26] <= WeightsStore9[166];
			WeightsStore9[27] <= WeightsStore9[167];
		end else if(switchCounter == 32'd41)begin
			PixelsStore[0] <= PixelsStore[168];
			PixelsStore[1] <= PixelsStore[169];
			PixelsStore[2] <= PixelsStore[170];
			PixelsStore[3] <= PixelsStore[171];
			PixelsStore[4] <= PixelsStore[172];
			PixelsStore[5] <= PixelsStore[173];
			PixelsStore[6] <= PixelsStore[174];
			PixelsStore[7] <= PixelsStore[175];
			PixelsStore[8] <= PixelsStore[176];
			PixelsStore[9] <= PixelsStore[177];
			PixelsStore[10] <= PixelsStore[178];
			PixelsStore[11] <= PixelsStore[179];
			PixelsStore[12] <= PixelsStore[180];
			PixelsStore[13] <= PixelsStore[181];
			PixelsStore[14] <= PixelsStore[182];
			PixelsStore[15] <= PixelsStore[183];
			PixelsStore[16] <= PixelsStore[184];
			PixelsStore[17] <= PixelsStore[185];
			PixelsStore[18] <= PixelsStore[186];
			PixelsStore[19] <= PixelsStore[187];
			PixelsStore[20] <= PixelsStore[188];
			PixelsStore[21] <= PixelsStore[189];
			PixelsStore[22] <= PixelsStore[190];
			PixelsStore[23] <= PixelsStore[191];
			PixelsStore[24] <= PixelsStore[192];
			PixelsStore[25] <= PixelsStore[193];
			PixelsStore[26] <= PixelsStore[194];
			PixelsStore[27] <= PixelsStore[195];
			WeightsStore0[0] <= WeightsStore0[168];
			WeightsStore0[1] <= WeightsStore0[169];
			WeightsStore0[2] <= WeightsStore0[170];
			WeightsStore0[3] <= WeightsStore0[171];
			WeightsStore0[4] <= WeightsStore0[172];
			WeightsStore0[5] <= WeightsStore0[173];
			WeightsStore0[6] <= WeightsStore0[174];
			WeightsStore0[7] <= WeightsStore0[175];
			WeightsStore0[8] <= WeightsStore0[176];
			WeightsStore0[9] <= WeightsStore0[177];
			WeightsStore0[10] <= WeightsStore0[178];
			WeightsStore0[11] <= WeightsStore0[179];
			WeightsStore0[12] <= WeightsStore0[180];
			WeightsStore0[13] <= WeightsStore0[181];
			WeightsStore0[14] <= WeightsStore0[182];
			WeightsStore0[15] <= WeightsStore0[183];
			WeightsStore0[16] <= WeightsStore0[184];
			WeightsStore0[17] <= WeightsStore0[185];
			WeightsStore0[18] <= WeightsStore0[186];
			WeightsStore0[19] <= WeightsStore0[187];
			WeightsStore0[20] <= WeightsStore0[188];
			WeightsStore0[21] <= WeightsStore0[189];
			WeightsStore0[22] <= WeightsStore0[190];
			WeightsStore0[23] <= WeightsStore0[191];
			WeightsStore0[24] <= WeightsStore0[192];
			WeightsStore0[25] <= WeightsStore0[193];
			WeightsStore0[26] <= WeightsStore0[194];
			WeightsStore0[27] <= WeightsStore0[195];
			WeightsStore1[0] <= WeightsStore1[168];
			WeightsStore1[1] <= WeightsStore1[169];
			WeightsStore1[2] <= WeightsStore1[170];
			WeightsStore1[3] <= WeightsStore1[171];
			WeightsStore1[4] <= WeightsStore1[172];
			WeightsStore1[5] <= WeightsStore1[173];
			WeightsStore1[6] <= WeightsStore1[174];
			WeightsStore1[7] <= WeightsStore1[175];
			WeightsStore1[8] <= WeightsStore1[176];
			WeightsStore1[9] <= WeightsStore1[177];
			WeightsStore1[10] <= WeightsStore1[178];
			WeightsStore1[11] <= WeightsStore1[179];
			WeightsStore1[12] <= WeightsStore1[180];
			WeightsStore1[13] <= WeightsStore1[181];
			WeightsStore1[14] <= WeightsStore1[182];
			WeightsStore1[15] <= WeightsStore1[183];
			WeightsStore1[16] <= WeightsStore1[184];
			WeightsStore1[17] <= WeightsStore1[185];
			WeightsStore1[18] <= WeightsStore1[186];
			WeightsStore1[19] <= WeightsStore1[187];
			WeightsStore1[20] <= WeightsStore1[188];
			WeightsStore1[21] <= WeightsStore1[189];
			WeightsStore1[22] <= WeightsStore1[190];
			WeightsStore1[23] <= WeightsStore1[191];
			WeightsStore1[24] <= WeightsStore1[192];
			WeightsStore1[25] <= WeightsStore1[193];
			WeightsStore1[26] <= WeightsStore1[194];
			WeightsStore1[27] <= WeightsStore1[195];
			WeightsStore2[0] <= WeightsStore2[168];
			WeightsStore2[1] <= WeightsStore2[169];
			WeightsStore2[2] <= WeightsStore2[170];
			WeightsStore2[3] <= WeightsStore2[171];
			WeightsStore2[4] <= WeightsStore2[172];
			WeightsStore2[5] <= WeightsStore2[173];
			WeightsStore2[6] <= WeightsStore2[174];
			WeightsStore2[7] <= WeightsStore2[175];
			WeightsStore2[8] <= WeightsStore2[176];
			WeightsStore2[9] <= WeightsStore2[177];
			WeightsStore2[10] <= WeightsStore2[178];
			WeightsStore2[11] <= WeightsStore2[179];
			WeightsStore2[12] <= WeightsStore2[180];
			WeightsStore2[13] <= WeightsStore2[181];
			WeightsStore2[14] <= WeightsStore2[182];
			WeightsStore2[15] <= WeightsStore2[183];
			WeightsStore2[16] <= WeightsStore2[184];
			WeightsStore2[17] <= WeightsStore2[185];
			WeightsStore2[18] <= WeightsStore2[186];
			WeightsStore2[19] <= WeightsStore2[187];
			WeightsStore2[20] <= WeightsStore2[188];
			WeightsStore2[21] <= WeightsStore2[189];
			WeightsStore2[22] <= WeightsStore2[190];
			WeightsStore2[23] <= WeightsStore2[191];
			WeightsStore2[24] <= WeightsStore2[192];
			WeightsStore2[25] <= WeightsStore2[193];
			WeightsStore2[26] <= WeightsStore2[194];
			WeightsStore2[27] <= WeightsStore2[195];
			WeightsStore3[0] <= WeightsStore3[168];
			WeightsStore3[1] <= WeightsStore3[169];
			WeightsStore3[2] <= WeightsStore3[170];
			WeightsStore3[3] <= WeightsStore3[171];
			WeightsStore3[4] <= WeightsStore3[172];
			WeightsStore3[5] <= WeightsStore3[173];
			WeightsStore3[6] <= WeightsStore3[174];
			WeightsStore3[7] <= WeightsStore3[175];
			WeightsStore3[8] <= WeightsStore3[176];
			WeightsStore3[9] <= WeightsStore3[177];
			WeightsStore3[10] <= WeightsStore3[178];
			WeightsStore3[11] <= WeightsStore3[179];
			WeightsStore3[12] <= WeightsStore3[180];
			WeightsStore3[13] <= WeightsStore3[181];
			WeightsStore3[14] <= WeightsStore3[182];
			WeightsStore3[15] <= WeightsStore3[183];
			WeightsStore3[16] <= WeightsStore3[184];
			WeightsStore3[17] <= WeightsStore3[185];
			WeightsStore3[18] <= WeightsStore3[186];
			WeightsStore3[19] <= WeightsStore3[187];
			WeightsStore3[20] <= WeightsStore3[188];
			WeightsStore3[21] <= WeightsStore3[189];
			WeightsStore3[22] <= WeightsStore3[190];
			WeightsStore3[23] <= WeightsStore3[191];
			WeightsStore3[24] <= WeightsStore3[192];
			WeightsStore3[25] <= WeightsStore3[193];
			WeightsStore3[26] <= WeightsStore3[194];
			WeightsStore3[27] <= WeightsStore3[195];
			WeightsStore4[0] <= WeightsStore4[168];
			WeightsStore4[1] <= WeightsStore4[169];
			WeightsStore4[2] <= WeightsStore4[170];
			WeightsStore4[3] <= WeightsStore4[171];
			WeightsStore4[4] <= WeightsStore4[172];
			WeightsStore4[5] <= WeightsStore4[173];
			WeightsStore4[6] <= WeightsStore4[174];
			WeightsStore4[7] <= WeightsStore4[175];
			WeightsStore4[8] <= WeightsStore4[176];
			WeightsStore4[9] <= WeightsStore4[177];
			WeightsStore4[10] <= WeightsStore4[178];
			WeightsStore4[11] <= WeightsStore4[179];
			WeightsStore4[12] <= WeightsStore4[180];
			WeightsStore4[13] <= WeightsStore4[181];
			WeightsStore4[14] <= WeightsStore4[182];
			WeightsStore4[15] <= WeightsStore4[183];
			WeightsStore4[16] <= WeightsStore4[184];
			WeightsStore4[17] <= WeightsStore4[185];
			WeightsStore4[18] <= WeightsStore4[186];
			WeightsStore4[19] <= WeightsStore4[187];
			WeightsStore4[20] <= WeightsStore4[188];
			WeightsStore4[21] <= WeightsStore4[189];
			WeightsStore4[22] <= WeightsStore4[190];
			WeightsStore4[23] <= WeightsStore4[191];
			WeightsStore4[24] <= WeightsStore4[192];
			WeightsStore4[25] <= WeightsStore4[193];
			WeightsStore4[26] <= WeightsStore4[194];
			WeightsStore4[27] <= WeightsStore4[195];
			WeightsStore5[0] <= WeightsStore5[168];
			WeightsStore5[1] <= WeightsStore5[169];
			WeightsStore5[2] <= WeightsStore5[170];
			WeightsStore5[3] <= WeightsStore5[171];
			WeightsStore5[4] <= WeightsStore5[172];
			WeightsStore5[5] <= WeightsStore5[173];
			WeightsStore5[6] <= WeightsStore5[174];
			WeightsStore5[7] <= WeightsStore5[175];
			WeightsStore5[8] <= WeightsStore5[176];
			WeightsStore5[9] <= WeightsStore5[177];
			WeightsStore5[10] <= WeightsStore5[178];
			WeightsStore5[11] <= WeightsStore5[179];
			WeightsStore5[12] <= WeightsStore5[180];
			WeightsStore5[13] <= WeightsStore5[181];
			WeightsStore5[14] <= WeightsStore5[182];
			WeightsStore5[15] <= WeightsStore5[183];
			WeightsStore5[16] <= WeightsStore5[184];
			WeightsStore5[17] <= WeightsStore5[185];
			WeightsStore5[18] <= WeightsStore5[186];
			WeightsStore5[19] <= WeightsStore5[187];
			WeightsStore5[20] <= WeightsStore5[188];
			WeightsStore5[21] <= WeightsStore5[189];
			WeightsStore5[22] <= WeightsStore5[190];
			WeightsStore5[23] <= WeightsStore5[191];
			WeightsStore5[24] <= WeightsStore5[192];
			WeightsStore5[25] <= WeightsStore5[193];
			WeightsStore5[26] <= WeightsStore5[194];
			WeightsStore5[27] <= WeightsStore5[195];
			WeightsStore6[0] <= WeightsStore6[168];
			WeightsStore6[1] <= WeightsStore6[169];
			WeightsStore6[2] <= WeightsStore6[170];
			WeightsStore6[3] <= WeightsStore6[171];
			WeightsStore6[4] <= WeightsStore6[172];
			WeightsStore6[5] <= WeightsStore6[173];
			WeightsStore6[6] <= WeightsStore6[174];
			WeightsStore6[7] <= WeightsStore6[175];
			WeightsStore6[8] <= WeightsStore6[176];
			WeightsStore6[9] <= WeightsStore6[177];
			WeightsStore6[10] <= WeightsStore6[178];
			WeightsStore6[11] <= WeightsStore6[179];
			WeightsStore6[12] <= WeightsStore6[180];
			WeightsStore6[13] <= WeightsStore6[181];
			WeightsStore6[14] <= WeightsStore6[182];
			WeightsStore6[15] <= WeightsStore6[183];
			WeightsStore6[16] <= WeightsStore6[184];
			WeightsStore6[17] <= WeightsStore6[185];
			WeightsStore6[18] <= WeightsStore6[186];
			WeightsStore6[19] <= WeightsStore6[187];
			WeightsStore6[20] <= WeightsStore6[188];
			WeightsStore6[21] <= WeightsStore6[189];
			WeightsStore6[22] <= WeightsStore6[190];
			WeightsStore6[23] <= WeightsStore6[191];
			WeightsStore6[24] <= WeightsStore6[192];
			WeightsStore6[25] <= WeightsStore6[193];
			WeightsStore6[26] <= WeightsStore6[194];
			WeightsStore6[27] <= WeightsStore6[195];
			WeightsStore7[0] <= WeightsStore7[168];
			WeightsStore7[1] <= WeightsStore7[169];
			WeightsStore7[2] <= WeightsStore7[170];
			WeightsStore7[3] <= WeightsStore7[171];
			WeightsStore7[4] <= WeightsStore7[172];
			WeightsStore7[5] <= WeightsStore7[173];
			WeightsStore7[6] <= WeightsStore7[174];
			WeightsStore7[7] <= WeightsStore7[175];
			WeightsStore7[8] <= WeightsStore7[176];
			WeightsStore7[9] <= WeightsStore7[177];
			WeightsStore7[10] <= WeightsStore7[178];
			WeightsStore7[11] <= WeightsStore7[179];
			WeightsStore7[12] <= WeightsStore7[180];
			WeightsStore7[13] <= WeightsStore7[181];
			WeightsStore7[14] <= WeightsStore7[182];
			WeightsStore7[15] <= WeightsStore7[183];
			WeightsStore7[16] <= WeightsStore7[184];
			WeightsStore7[17] <= WeightsStore7[185];
			WeightsStore7[18] <= WeightsStore7[186];
			WeightsStore7[19] <= WeightsStore7[187];
			WeightsStore7[20] <= WeightsStore7[188];
			WeightsStore7[21] <= WeightsStore7[189];
			WeightsStore7[22] <= WeightsStore7[190];
			WeightsStore7[23] <= WeightsStore7[191];
			WeightsStore7[24] <= WeightsStore7[192];
			WeightsStore7[25] <= WeightsStore7[193];
			WeightsStore7[26] <= WeightsStore7[194];
			WeightsStore7[27] <= WeightsStore7[195];
			WeightsStore8[0] <= WeightsStore8[168];
			WeightsStore8[1] <= WeightsStore8[169];
			WeightsStore8[2] <= WeightsStore8[170];
			WeightsStore8[3] <= WeightsStore8[171];
			WeightsStore8[4] <= WeightsStore8[172];
			WeightsStore8[5] <= WeightsStore8[173];
			WeightsStore8[6] <= WeightsStore8[174];
			WeightsStore8[7] <= WeightsStore8[175];
			WeightsStore8[8] <= WeightsStore8[176];
			WeightsStore8[9] <= WeightsStore8[177];
			WeightsStore8[10] <= WeightsStore8[178];
			WeightsStore8[11] <= WeightsStore8[179];
			WeightsStore8[12] <= WeightsStore8[180];
			WeightsStore8[13] <= WeightsStore8[181];
			WeightsStore8[14] <= WeightsStore8[182];
			WeightsStore8[15] <= WeightsStore8[183];
			WeightsStore8[16] <= WeightsStore8[184];
			WeightsStore8[17] <= WeightsStore8[185];
			WeightsStore8[18] <= WeightsStore8[186];
			WeightsStore8[19] <= WeightsStore8[187];
			WeightsStore8[20] <= WeightsStore8[188];
			WeightsStore8[21] <= WeightsStore8[189];
			WeightsStore8[22] <= WeightsStore8[190];
			WeightsStore8[23] <= WeightsStore8[191];
			WeightsStore8[24] <= WeightsStore8[192];
			WeightsStore8[25] <= WeightsStore8[193];
			WeightsStore8[26] <= WeightsStore8[194];
			WeightsStore8[27] <= WeightsStore8[195];
			WeightsStore9[0] <= WeightsStore9[168];
			WeightsStore9[1] <= WeightsStore9[169];
			WeightsStore9[2] <= WeightsStore9[170];
			WeightsStore9[3] <= WeightsStore9[171];
			WeightsStore9[4] <= WeightsStore9[172];
			WeightsStore9[5] <= WeightsStore9[173];
			WeightsStore9[6] <= WeightsStore9[174];
			WeightsStore9[7] <= WeightsStore9[175];
			WeightsStore9[8] <= WeightsStore9[176];
			WeightsStore9[9] <= WeightsStore9[177];
			WeightsStore9[10] <= WeightsStore9[178];
			WeightsStore9[11] <= WeightsStore9[179];
			WeightsStore9[12] <= WeightsStore9[180];
			WeightsStore9[13] <= WeightsStore9[181];
			WeightsStore9[14] <= WeightsStore9[182];
			WeightsStore9[15] <= WeightsStore9[183];
			WeightsStore9[16] <= WeightsStore9[184];
			WeightsStore9[17] <= WeightsStore9[185];
			WeightsStore9[18] <= WeightsStore9[186];
			WeightsStore9[19] <= WeightsStore9[187];
			WeightsStore9[20] <= WeightsStore9[188];
			WeightsStore9[21] <= WeightsStore9[189];
			WeightsStore9[22] <= WeightsStore9[190];
			WeightsStore9[23] <= WeightsStore9[191];
			WeightsStore9[24] <= WeightsStore9[192];
			WeightsStore9[25] <= WeightsStore9[193];
			WeightsStore9[26] <= WeightsStore9[194];
			WeightsStore9[27] <= WeightsStore9[195];
		end else if(switchCounter == 32'd48)begin
			PixelsStore[0] <= PixelsStore[196];
			PixelsStore[1] <= PixelsStore[197];
			PixelsStore[2] <= PixelsStore[198];
			PixelsStore[3] <= PixelsStore[199];
			PixelsStore[4] <= PixelsStore[200];
			PixelsStore[5] <= PixelsStore[201];
			PixelsStore[6] <= PixelsStore[202];
			PixelsStore[7] <= PixelsStore[203];
			PixelsStore[8] <= PixelsStore[204];
			PixelsStore[9] <= PixelsStore[205];
			PixelsStore[10] <= PixelsStore[206];
			PixelsStore[11] <= PixelsStore[207];
			PixelsStore[12] <= PixelsStore[208];
			PixelsStore[13] <= PixelsStore[209];
			PixelsStore[14] <= PixelsStore[210];
			PixelsStore[15] <= PixelsStore[211];
			PixelsStore[16] <= PixelsStore[212];
			PixelsStore[17] <= PixelsStore[213];
			PixelsStore[18] <= PixelsStore[214];
			PixelsStore[19] <= PixelsStore[215];
			PixelsStore[20] <= PixelsStore[216];
			PixelsStore[21] <= PixelsStore[217];
			PixelsStore[22] <= PixelsStore[218];
			PixelsStore[23] <= PixelsStore[219];
			PixelsStore[24] <= PixelsStore[220];
			PixelsStore[25] <= PixelsStore[221];
			PixelsStore[26] <= PixelsStore[222];
			PixelsStore[27] <= PixelsStore[223];
			WeightsStore0[0] <= WeightsStore0[196];
			WeightsStore0[1] <= WeightsStore0[197];
			WeightsStore0[2] <= WeightsStore0[198];
			WeightsStore0[3] <= WeightsStore0[199];
			WeightsStore0[4] <= WeightsStore0[200];
			WeightsStore0[5] <= WeightsStore0[201];
			WeightsStore0[6] <= WeightsStore0[202];
			WeightsStore0[7] <= WeightsStore0[203];
			WeightsStore0[8] <= WeightsStore0[204];
			WeightsStore0[9] <= WeightsStore0[205];
			WeightsStore0[10] <= WeightsStore0[206];
			WeightsStore0[11] <= WeightsStore0[207];
			WeightsStore0[12] <= WeightsStore0[208];
			WeightsStore0[13] <= WeightsStore0[209];
			WeightsStore0[14] <= WeightsStore0[210];
			WeightsStore0[15] <= WeightsStore0[211];
			WeightsStore0[16] <= WeightsStore0[212];
			WeightsStore0[17] <= WeightsStore0[213];
			WeightsStore0[18] <= WeightsStore0[214];
			WeightsStore0[19] <= WeightsStore0[215];
			WeightsStore0[20] <= WeightsStore0[216];
			WeightsStore0[21] <= WeightsStore0[217];
			WeightsStore0[22] <= WeightsStore0[218];
			WeightsStore0[23] <= WeightsStore0[219];
			WeightsStore0[24] <= WeightsStore0[220];
			WeightsStore0[25] <= WeightsStore0[221];
			WeightsStore0[26] <= WeightsStore0[222];
			WeightsStore0[27] <= WeightsStore0[223];
			WeightsStore1[0] <= WeightsStore1[196];
			WeightsStore1[1] <= WeightsStore1[197];
			WeightsStore1[2] <= WeightsStore1[198];
			WeightsStore1[3] <= WeightsStore1[199];
			WeightsStore1[4] <= WeightsStore1[200];
			WeightsStore1[5] <= WeightsStore1[201];
			WeightsStore1[6] <= WeightsStore1[202];
			WeightsStore1[7] <= WeightsStore1[203];
			WeightsStore1[8] <= WeightsStore1[204];
			WeightsStore1[9] <= WeightsStore1[205];
			WeightsStore1[10] <= WeightsStore1[206];
			WeightsStore1[11] <= WeightsStore1[207];
			WeightsStore1[12] <= WeightsStore1[208];
			WeightsStore1[13] <= WeightsStore1[209];
			WeightsStore1[14] <= WeightsStore1[210];
			WeightsStore1[15] <= WeightsStore1[211];
			WeightsStore1[16] <= WeightsStore1[212];
			WeightsStore1[17] <= WeightsStore1[213];
			WeightsStore1[18] <= WeightsStore1[214];
			WeightsStore1[19] <= WeightsStore1[215];
			WeightsStore1[20] <= WeightsStore1[216];
			WeightsStore1[21] <= WeightsStore1[217];
			WeightsStore1[22] <= WeightsStore1[218];
			WeightsStore1[23] <= WeightsStore1[219];
			WeightsStore1[24] <= WeightsStore1[220];
			WeightsStore1[25] <= WeightsStore1[221];
			WeightsStore1[26] <= WeightsStore1[222];
			WeightsStore1[27] <= WeightsStore1[223];
			WeightsStore2[0] <= WeightsStore2[196];
			WeightsStore2[1] <= WeightsStore2[197];
			WeightsStore2[2] <= WeightsStore2[198];
			WeightsStore2[3] <= WeightsStore2[199];
			WeightsStore2[4] <= WeightsStore2[200];
			WeightsStore2[5] <= WeightsStore2[201];
			WeightsStore2[6] <= WeightsStore2[202];
			WeightsStore2[7] <= WeightsStore2[203];
			WeightsStore2[8] <= WeightsStore2[204];
			WeightsStore2[9] <= WeightsStore2[205];
			WeightsStore2[10] <= WeightsStore2[206];
			WeightsStore2[11] <= WeightsStore2[207];
			WeightsStore2[12] <= WeightsStore2[208];
			WeightsStore2[13] <= WeightsStore2[209];
			WeightsStore2[14] <= WeightsStore2[210];
			WeightsStore2[15] <= WeightsStore2[211];
			WeightsStore2[16] <= WeightsStore2[212];
			WeightsStore2[17] <= WeightsStore2[213];
			WeightsStore2[18] <= WeightsStore2[214];
			WeightsStore2[19] <= WeightsStore2[215];
			WeightsStore2[20] <= WeightsStore2[216];
			WeightsStore2[21] <= WeightsStore2[217];
			WeightsStore2[22] <= WeightsStore2[218];
			WeightsStore2[23] <= WeightsStore2[219];
			WeightsStore2[24] <= WeightsStore2[220];
			WeightsStore2[25] <= WeightsStore2[221];
			WeightsStore2[26] <= WeightsStore2[222];
			WeightsStore2[27] <= WeightsStore2[223];
			WeightsStore3[0] <= WeightsStore3[196];
			WeightsStore3[1] <= WeightsStore3[197];
			WeightsStore3[2] <= WeightsStore3[198];
			WeightsStore3[3] <= WeightsStore3[199];
			WeightsStore3[4] <= WeightsStore3[200];
			WeightsStore3[5] <= WeightsStore3[201];
			WeightsStore3[6] <= WeightsStore3[202];
			WeightsStore3[7] <= WeightsStore3[203];
			WeightsStore3[8] <= WeightsStore3[204];
			WeightsStore3[9] <= WeightsStore3[205];
			WeightsStore3[10] <= WeightsStore3[206];
			WeightsStore3[11] <= WeightsStore3[207];
			WeightsStore3[12] <= WeightsStore3[208];
			WeightsStore3[13] <= WeightsStore3[209];
			WeightsStore3[14] <= WeightsStore3[210];
			WeightsStore3[15] <= WeightsStore3[211];
			WeightsStore3[16] <= WeightsStore3[212];
			WeightsStore3[17] <= WeightsStore3[213];
			WeightsStore3[18] <= WeightsStore3[214];
			WeightsStore3[19] <= WeightsStore3[215];
			WeightsStore3[20] <= WeightsStore3[216];
			WeightsStore3[21] <= WeightsStore3[217];
			WeightsStore3[22] <= WeightsStore3[218];
			WeightsStore3[23] <= WeightsStore3[219];
			WeightsStore3[24] <= WeightsStore3[220];
			WeightsStore3[25] <= WeightsStore3[221];
			WeightsStore3[26] <= WeightsStore3[222];
			WeightsStore3[27] <= WeightsStore3[223];
			WeightsStore4[0] <= WeightsStore4[196];
			WeightsStore4[1] <= WeightsStore4[197];
			WeightsStore4[2] <= WeightsStore4[198];
			WeightsStore4[3] <= WeightsStore4[199];
			WeightsStore4[4] <= WeightsStore4[200];
			WeightsStore4[5] <= WeightsStore4[201];
			WeightsStore4[6] <= WeightsStore4[202];
			WeightsStore4[7] <= WeightsStore4[203];
			WeightsStore4[8] <= WeightsStore4[204];
			WeightsStore4[9] <= WeightsStore4[205];
			WeightsStore4[10] <= WeightsStore4[206];
			WeightsStore4[11] <= WeightsStore4[207];
			WeightsStore4[12] <= WeightsStore4[208];
			WeightsStore4[13] <= WeightsStore4[209];
			WeightsStore4[14] <= WeightsStore4[210];
			WeightsStore4[15] <= WeightsStore4[211];
			WeightsStore4[16] <= WeightsStore4[212];
			WeightsStore4[17] <= WeightsStore4[213];
			WeightsStore4[18] <= WeightsStore4[214];
			WeightsStore4[19] <= WeightsStore4[215];
			WeightsStore4[20] <= WeightsStore4[216];
			WeightsStore4[21] <= WeightsStore4[217];
			WeightsStore4[22] <= WeightsStore4[218];
			WeightsStore4[23] <= WeightsStore4[219];
			WeightsStore4[24] <= WeightsStore4[220];
			WeightsStore4[25] <= WeightsStore4[221];
			WeightsStore4[26] <= WeightsStore4[222];
			WeightsStore4[27] <= WeightsStore4[223];
			WeightsStore5[0] <= WeightsStore5[196];
			WeightsStore5[1] <= WeightsStore5[197];
			WeightsStore5[2] <= WeightsStore5[198];
			WeightsStore5[3] <= WeightsStore5[199];
			WeightsStore5[4] <= WeightsStore5[200];
			WeightsStore5[5] <= WeightsStore5[201];
			WeightsStore5[6] <= WeightsStore5[202];
			WeightsStore5[7] <= WeightsStore5[203];
			WeightsStore5[8] <= WeightsStore5[204];
			WeightsStore5[9] <= WeightsStore5[205];
			WeightsStore5[10] <= WeightsStore5[206];
			WeightsStore5[11] <= WeightsStore5[207];
			WeightsStore5[12] <= WeightsStore5[208];
			WeightsStore5[13] <= WeightsStore5[209];
			WeightsStore5[14] <= WeightsStore5[210];
			WeightsStore5[15] <= WeightsStore5[211];
			WeightsStore5[16] <= WeightsStore5[212];
			WeightsStore5[17] <= WeightsStore5[213];
			WeightsStore5[18] <= WeightsStore5[214];
			WeightsStore5[19] <= WeightsStore5[215];
			WeightsStore5[20] <= WeightsStore5[216];
			WeightsStore5[21] <= WeightsStore5[217];
			WeightsStore5[22] <= WeightsStore5[218];
			WeightsStore5[23] <= WeightsStore5[219];
			WeightsStore5[24] <= WeightsStore5[220];
			WeightsStore5[25] <= WeightsStore5[221];
			WeightsStore5[26] <= WeightsStore5[222];
			WeightsStore5[27] <= WeightsStore5[223];
			WeightsStore6[0] <= WeightsStore6[196];
			WeightsStore6[1] <= WeightsStore6[197];
			WeightsStore6[2] <= WeightsStore6[198];
			WeightsStore6[3] <= WeightsStore6[199];
			WeightsStore6[4] <= WeightsStore6[200];
			WeightsStore6[5] <= WeightsStore6[201];
			WeightsStore6[6] <= WeightsStore6[202];
			WeightsStore6[7] <= WeightsStore6[203];
			WeightsStore6[8] <= WeightsStore6[204];
			WeightsStore6[9] <= WeightsStore6[205];
			WeightsStore6[10] <= WeightsStore6[206];
			WeightsStore6[11] <= WeightsStore6[207];
			WeightsStore6[12] <= WeightsStore6[208];
			WeightsStore6[13] <= WeightsStore6[209];
			WeightsStore6[14] <= WeightsStore6[210];
			WeightsStore6[15] <= WeightsStore6[211];
			WeightsStore6[16] <= WeightsStore6[212];
			WeightsStore6[17] <= WeightsStore6[213];
			WeightsStore6[18] <= WeightsStore6[214];
			WeightsStore6[19] <= WeightsStore6[215];
			WeightsStore6[20] <= WeightsStore6[216];
			WeightsStore6[21] <= WeightsStore6[217];
			WeightsStore6[22] <= WeightsStore6[218];
			WeightsStore6[23] <= WeightsStore6[219];
			WeightsStore6[24] <= WeightsStore6[220];
			WeightsStore6[25] <= WeightsStore6[221];
			WeightsStore6[26] <= WeightsStore6[222];
			WeightsStore6[27] <= WeightsStore6[223];
			WeightsStore7[0] <= WeightsStore7[196];
			WeightsStore7[1] <= WeightsStore7[197];
			WeightsStore7[2] <= WeightsStore7[198];
			WeightsStore7[3] <= WeightsStore7[199];
			WeightsStore7[4] <= WeightsStore7[200];
			WeightsStore7[5] <= WeightsStore7[201];
			WeightsStore7[6] <= WeightsStore7[202];
			WeightsStore7[7] <= WeightsStore7[203];
			WeightsStore7[8] <= WeightsStore7[204];
			WeightsStore7[9] <= WeightsStore7[205];
			WeightsStore7[10] <= WeightsStore7[206];
			WeightsStore7[11] <= WeightsStore7[207];
			WeightsStore7[12] <= WeightsStore7[208];
			WeightsStore7[13] <= WeightsStore7[209];
			WeightsStore7[14] <= WeightsStore7[210];
			WeightsStore7[15] <= WeightsStore7[211];
			WeightsStore7[16] <= WeightsStore7[212];
			WeightsStore7[17] <= WeightsStore7[213];
			WeightsStore7[18] <= WeightsStore7[214];
			WeightsStore7[19] <= WeightsStore7[215];
			WeightsStore7[20] <= WeightsStore7[216];
			WeightsStore7[21] <= WeightsStore7[217];
			WeightsStore7[22] <= WeightsStore7[218];
			WeightsStore7[23] <= WeightsStore7[219];
			WeightsStore7[24] <= WeightsStore7[220];
			WeightsStore7[25] <= WeightsStore7[221];
			WeightsStore7[26] <= WeightsStore7[222];
			WeightsStore7[27] <= WeightsStore7[223];
			WeightsStore8[0] <= WeightsStore8[196];
			WeightsStore8[1] <= WeightsStore8[197];
			WeightsStore8[2] <= WeightsStore8[198];
			WeightsStore8[3] <= WeightsStore8[199];
			WeightsStore8[4] <= WeightsStore8[200];
			WeightsStore8[5] <= WeightsStore8[201];
			WeightsStore8[6] <= WeightsStore8[202];
			WeightsStore8[7] <= WeightsStore8[203];
			WeightsStore8[8] <= WeightsStore8[204];
			WeightsStore8[9] <= WeightsStore8[205];
			WeightsStore8[10] <= WeightsStore8[206];
			WeightsStore8[11] <= WeightsStore8[207];
			WeightsStore8[12] <= WeightsStore8[208];
			WeightsStore8[13] <= WeightsStore8[209];
			WeightsStore8[14] <= WeightsStore8[210];
			WeightsStore8[15] <= WeightsStore8[211];
			WeightsStore8[16] <= WeightsStore8[212];
			WeightsStore8[17] <= WeightsStore8[213];
			WeightsStore8[18] <= WeightsStore8[214];
			WeightsStore8[19] <= WeightsStore8[215];
			WeightsStore8[20] <= WeightsStore8[216];
			WeightsStore8[21] <= WeightsStore8[217];
			WeightsStore8[22] <= WeightsStore8[218];
			WeightsStore8[23] <= WeightsStore8[219];
			WeightsStore8[24] <= WeightsStore8[220];
			WeightsStore8[25] <= WeightsStore8[221];
			WeightsStore8[26] <= WeightsStore8[222];
			WeightsStore8[27] <= WeightsStore8[223];
			WeightsStore9[0] <= WeightsStore9[196];
			WeightsStore9[1] <= WeightsStore9[197];
			WeightsStore9[2] <= WeightsStore9[198];
			WeightsStore9[3] <= WeightsStore9[199];
			WeightsStore9[4] <= WeightsStore9[200];
			WeightsStore9[5] <= WeightsStore9[201];
			WeightsStore9[6] <= WeightsStore9[202];
			WeightsStore9[7] <= WeightsStore9[203];
			WeightsStore9[8] <= WeightsStore9[204];
			WeightsStore9[9] <= WeightsStore9[205];
			WeightsStore9[10] <= WeightsStore9[206];
			WeightsStore9[11] <= WeightsStore9[207];
			WeightsStore9[12] <= WeightsStore9[208];
			WeightsStore9[13] <= WeightsStore9[209];
			WeightsStore9[14] <= WeightsStore9[210];
			WeightsStore9[15] <= WeightsStore9[211];
			WeightsStore9[16] <= WeightsStore9[212];
			WeightsStore9[17] <= WeightsStore9[213];
			WeightsStore9[18] <= WeightsStore9[214];
			WeightsStore9[19] <= WeightsStore9[215];
			WeightsStore9[20] <= WeightsStore9[216];
			WeightsStore9[21] <= WeightsStore9[217];
			WeightsStore9[22] <= WeightsStore9[218];
			WeightsStore9[23] <= WeightsStore9[219];
			WeightsStore9[24] <= WeightsStore9[220];
			WeightsStore9[25] <= WeightsStore9[221];
			WeightsStore9[26] <= WeightsStore9[222];
			WeightsStore9[27] <= WeightsStore9[223];
		end else if(switchCounter == 32'd55)begin
			PixelsStore[0] <= PixelsStore[224];
			PixelsStore[1] <= PixelsStore[225];
			PixelsStore[2] <= PixelsStore[226];
			PixelsStore[3] <= PixelsStore[227];
			PixelsStore[4] <= PixelsStore[228];
			PixelsStore[5] <= PixelsStore[229];
			PixelsStore[6] <= PixelsStore[230];
			PixelsStore[7] <= PixelsStore[231];
			PixelsStore[8] <= PixelsStore[232];
			PixelsStore[9] <= PixelsStore[233];
			PixelsStore[10] <= PixelsStore[234];
			PixelsStore[11] <= PixelsStore[235];
			PixelsStore[12] <= PixelsStore[236];
			PixelsStore[13] <= PixelsStore[237];
			PixelsStore[14] <= PixelsStore[238];
			PixelsStore[15] <= PixelsStore[239];
			PixelsStore[16] <= PixelsStore[240];
			PixelsStore[17] <= PixelsStore[241];
			PixelsStore[18] <= PixelsStore[242];
			PixelsStore[19] <= PixelsStore[243];
			PixelsStore[20] <= PixelsStore[244];
			PixelsStore[21] <= PixelsStore[245];
			PixelsStore[22] <= PixelsStore[246];
			PixelsStore[23] <= PixelsStore[247];
			PixelsStore[24] <= PixelsStore[248];
			PixelsStore[25] <= PixelsStore[249];
			PixelsStore[26] <= PixelsStore[250];
			PixelsStore[27] <= PixelsStore[251];
			WeightsStore0[0] <= WeightsStore0[224];
			WeightsStore0[1] <= WeightsStore0[225];
			WeightsStore0[2] <= WeightsStore0[226];
			WeightsStore0[3] <= WeightsStore0[227];
			WeightsStore0[4] <= WeightsStore0[228];
			WeightsStore0[5] <= WeightsStore0[229];
			WeightsStore0[6] <= WeightsStore0[230];
			WeightsStore0[7] <= WeightsStore0[231];
			WeightsStore0[8] <= WeightsStore0[232];
			WeightsStore0[9] <= WeightsStore0[233];
			WeightsStore0[10] <= WeightsStore0[234];
			WeightsStore0[11] <= WeightsStore0[235];
			WeightsStore0[12] <= WeightsStore0[236];
			WeightsStore0[13] <= WeightsStore0[237];
			WeightsStore0[14] <= WeightsStore0[238];
			WeightsStore0[15] <= WeightsStore0[239];
			WeightsStore0[16] <= WeightsStore0[240];
			WeightsStore0[17] <= WeightsStore0[241];
			WeightsStore0[18] <= WeightsStore0[242];
			WeightsStore0[19] <= WeightsStore0[243];
			WeightsStore0[20] <= WeightsStore0[244];
			WeightsStore0[21] <= WeightsStore0[245];
			WeightsStore0[22] <= WeightsStore0[246];
			WeightsStore0[23] <= WeightsStore0[247];
			WeightsStore0[24] <= WeightsStore0[248];
			WeightsStore0[25] <= WeightsStore0[249];
			WeightsStore0[26] <= WeightsStore0[250];
			WeightsStore0[27] <= WeightsStore0[251];
			WeightsStore1[0] <= WeightsStore1[224];
			WeightsStore1[1] <= WeightsStore1[225];
			WeightsStore1[2] <= WeightsStore1[226];
			WeightsStore1[3] <= WeightsStore1[227];
			WeightsStore1[4] <= WeightsStore1[228];
			WeightsStore1[5] <= WeightsStore1[229];
			WeightsStore1[6] <= WeightsStore1[230];
			WeightsStore1[7] <= WeightsStore1[231];
			WeightsStore1[8] <= WeightsStore1[232];
			WeightsStore1[9] <= WeightsStore1[233];
			WeightsStore1[10] <= WeightsStore1[234];
			WeightsStore1[11] <= WeightsStore1[235];
			WeightsStore1[12] <= WeightsStore1[236];
			WeightsStore1[13] <= WeightsStore1[237];
			WeightsStore1[14] <= WeightsStore1[238];
			WeightsStore1[15] <= WeightsStore1[239];
			WeightsStore1[16] <= WeightsStore1[240];
			WeightsStore1[17] <= WeightsStore1[241];
			WeightsStore1[18] <= WeightsStore1[242];
			WeightsStore1[19] <= WeightsStore1[243];
			WeightsStore1[20] <= WeightsStore1[244];
			WeightsStore1[21] <= WeightsStore1[245];
			WeightsStore1[22] <= WeightsStore1[246];
			WeightsStore1[23] <= WeightsStore1[247];
			WeightsStore1[24] <= WeightsStore1[248];
			WeightsStore1[25] <= WeightsStore1[249];
			WeightsStore1[26] <= WeightsStore1[250];
			WeightsStore1[27] <= WeightsStore1[251];
			WeightsStore2[0] <= WeightsStore2[224];
			WeightsStore2[1] <= WeightsStore2[225];
			WeightsStore2[2] <= WeightsStore2[226];
			WeightsStore2[3] <= WeightsStore2[227];
			WeightsStore2[4] <= WeightsStore2[228];
			WeightsStore2[5] <= WeightsStore2[229];
			WeightsStore2[6] <= WeightsStore2[230];
			WeightsStore2[7] <= WeightsStore2[231];
			WeightsStore2[8] <= WeightsStore2[232];
			WeightsStore2[9] <= WeightsStore2[233];
			WeightsStore2[10] <= WeightsStore2[234];
			WeightsStore2[11] <= WeightsStore2[235];
			WeightsStore2[12] <= WeightsStore2[236];
			WeightsStore2[13] <= WeightsStore2[237];
			WeightsStore2[14] <= WeightsStore2[238];
			WeightsStore2[15] <= WeightsStore2[239];
			WeightsStore2[16] <= WeightsStore2[240];
			WeightsStore2[17] <= WeightsStore2[241];
			WeightsStore2[18] <= WeightsStore2[242];
			WeightsStore2[19] <= WeightsStore2[243];
			WeightsStore2[20] <= WeightsStore2[244];
			WeightsStore2[21] <= WeightsStore2[245];
			WeightsStore2[22] <= WeightsStore2[246];
			WeightsStore2[23] <= WeightsStore2[247];
			WeightsStore2[24] <= WeightsStore2[248];
			WeightsStore2[25] <= WeightsStore2[249];
			WeightsStore2[26] <= WeightsStore2[250];
			WeightsStore2[27] <= WeightsStore2[251];
			WeightsStore3[0] <= WeightsStore3[224];
			WeightsStore3[1] <= WeightsStore3[225];
			WeightsStore3[2] <= WeightsStore3[226];
			WeightsStore3[3] <= WeightsStore3[227];
			WeightsStore3[4] <= WeightsStore3[228];
			WeightsStore3[5] <= WeightsStore3[229];
			WeightsStore3[6] <= WeightsStore3[230];
			WeightsStore3[7] <= WeightsStore3[231];
			WeightsStore3[8] <= WeightsStore3[232];
			WeightsStore3[9] <= WeightsStore3[233];
			WeightsStore3[10] <= WeightsStore3[234];
			WeightsStore3[11] <= WeightsStore3[235];
			WeightsStore3[12] <= WeightsStore3[236];
			WeightsStore3[13] <= WeightsStore3[237];
			WeightsStore3[14] <= WeightsStore3[238];
			WeightsStore3[15] <= WeightsStore3[239];
			WeightsStore3[16] <= WeightsStore3[240];
			WeightsStore3[17] <= WeightsStore3[241];
			WeightsStore3[18] <= WeightsStore3[242];
			WeightsStore3[19] <= WeightsStore3[243];
			WeightsStore3[20] <= WeightsStore3[244];
			WeightsStore3[21] <= WeightsStore3[245];
			WeightsStore3[22] <= WeightsStore3[246];
			WeightsStore3[23] <= WeightsStore3[247];
			WeightsStore3[24] <= WeightsStore3[248];
			WeightsStore3[25] <= WeightsStore3[249];
			WeightsStore3[26] <= WeightsStore3[250];
			WeightsStore3[27] <= WeightsStore3[251];
			WeightsStore4[0] <= WeightsStore4[224];
			WeightsStore4[1] <= WeightsStore4[225];
			WeightsStore4[2] <= WeightsStore4[226];
			WeightsStore4[3] <= WeightsStore4[227];
			WeightsStore4[4] <= WeightsStore4[228];
			WeightsStore4[5] <= WeightsStore4[229];
			WeightsStore4[6] <= WeightsStore4[230];
			WeightsStore4[7] <= WeightsStore4[231];
			WeightsStore4[8] <= WeightsStore4[232];
			WeightsStore4[9] <= WeightsStore4[233];
			WeightsStore4[10] <= WeightsStore4[234];
			WeightsStore4[11] <= WeightsStore4[235];
			WeightsStore4[12] <= WeightsStore4[236];
			WeightsStore4[13] <= WeightsStore4[237];
			WeightsStore4[14] <= WeightsStore4[238];
			WeightsStore4[15] <= WeightsStore4[239];
			WeightsStore4[16] <= WeightsStore4[240];
			WeightsStore4[17] <= WeightsStore4[241];
			WeightsStore4[18] <= WeightsStore4[242];
			WeightsStore4[19] <= WeightsStore4[243];
			WeightsStore4[20] <= WeightsStore4[244];
			WeightsStore4[21] <= WeightsStore4[245];
			WeightsStore4[22] <= WeightsStore4[246];
			WeightsStore4[23] <= WeightsStore4[247];
			WeightsStore4[24] <= WeightsStore4[248];
			WeightsStore4[25] <= WeightsStore4[249];
			WeightsStore4[26] <= WeightsStore4[250];
			WeightsStore4[27] <= WeightsStore4[251];
			WeightsStore5[0] <= WeightsStore5[224];
			WeightsStore5[1] <= WeightsStore5[225];
			WeightsStore5[2] <= WeightsStore5[226];
			WeightsStore5[3] <= WeightsStore5[227];
			WeightsStore5[4] <= WeightsStore5[228];
			WeightsStore5[5] <= WeightsStore5[229];
			WeightsStore5[6] <= WeightsStore5[230];
			WeightsStore5[7] <= WeightsStore5[231];
			WeightsStore5[8] <= WeightsStore5[232];
			WeightsStore5[9] <= WeightsStore5[233];
			WeightsStore5[10] <= WeightsStore5[234];
			WeightsStore5[11] <= WeightsStore5[235];
			WeightsStore5[12] <= WeightsStore5[236];
			WeightsStore5[13] <= WeightsStore5[237];
			WeightsStore5[14] <= WeightsStore5[238];
			WeightsStore5[15] <= WeightsStore5[239];
			WeightsStore5[16] <= WeightsStore5[240];
			WeightsStore5[17] <= WeightsStore5[241];
			WeightsStore5[18] <= WeightsStore5[242];
			WeightsStore5[19] <= WeightsStore5[243];
			WeightsStore5[20] <= WeightsStore5[244];
			WeightsStore5[21] <= WeightsStore5[245];
			WeightsStore5[22] <= WeightsStore5[246];
			WeightsStore5[23] <= WeightsStore5[247];
			WeightsStore5[24] <= WeightsStore5[248];
			WeightsStore5[25] <= WeightsStore5[249];
			WeightsStore5[26] <= WeightsStore5[250];
			WeightsStore5[27] <= WeightsStore5[251];
			WeightsStore6[0] <= WeightsStore6[224];
			WeightsStore6[1] <= WeightsStore6[225];
			WeightsStore6[2] <= WeightsStore6[226];
			WeightsStore6[3] <= WeightsStore6[227];
			WeightsStore6[4] <= WeightsStore6[228];
			WeightsStore6[5] <= WeightsStore6[229];
			WeightsStore6[6] <= WeightsStore6[230];
			WeightsStore6[7] <= WeightsStore6[231];
			WeightsStore6[8] <= WeightsStore6[232];
			WeightsStore6[9] <= WeightsStore6[233];
			WeightsStore6[10] <= WeightsStore6[234];
			WeightsStore6[11] <= WeightsStore6[235];
			WeightsStore6[12] <= WeightsStore6[236];
			WeightsStore6[13] <= WeightsStore6[237];
			WeightsStore6[14] <= WeightsStore6[238];
			WeightsStore6[15] <= WeightsStore6[239];
			WeightsStore6[16] <= WeightsStore6[240];
			WeightsStore6[17] <= WeightsStore6[241];
			WeightsStore6[18] <= WeightsStore6[242];
			WeightsStore6[19] <= WeightsStore6[243];
			WeightsStore6[20] <= WeightsStore6[244];
			WeightsStore6[21] <= WeightsStore6[245];
			WeightsStore6[22] <= WeightsStore6[246];
			WeightsStore6[23] <= WeightsStore6[247];
			WeightsStore6[24] <= WeightsStore6[248];
			WeightsStore6[25] <= WeightsStore6[249];
			WeightsStore6[26] <= WeightsStore6[250];
			WeightsStore6[27] <= WeightsStore6[251];
			WeightsStore7[0] <= WeightsStore7[224];
			WeightsStore7[1] <= WeightsStore7[225];
			WeightsStore7[2] <= WeightsStore7[226];
			WeightsStore7[3] <= WeightsStore7[227];
			WeightsStore7[4] <= WeightsStore7[228];
			WeightsStore7[5] <= WeightsStore7[229];
			WeightsStore7[6] <= WeightsStore7[230];
			WeightsStore7[7] <= WeightsStore7[231];
			WeightsStore7[8] <= WeightsStore7[232];
			WeightsStore7[9] <= WeightsStore7[233];
			WeightsStore7[10] <= WeightsStore7[234];
			WeightsStore7[11] <= WeightsStore7[235];
			WeightsStore7[12] <= WeightsStore7[236];
			WeightsStore7[13] <= WeightsStore7[237];
			WeightsStore7[14] <= WeightsStore7[238];
			WeightsStore7[15] <= WeightsStore7[239];
			WeightsStore7[16] <= WeightsStore7[240];
			WeightsStore7[17] <= WeightsStore7[241];
			WeightsStore7[18] <= WeightsStore7[242];
			WeightsStore7[19] <= WeightsStore7[243];
			WeightsStore7[20] <= WeightsStore7[244];
			WeightsStore7[21] <= WeightsStore7[245];
			WeightsStore7[22] <= WeightsStore7[246];
			WeightsStore7[23] <= WeightsStore7[247];
			WeightsStore7[24] <= WeightsStore7[248];
			WeightsStore7[25] <= WeightsStore7[249];
			WeightsStore7[26] <= WeightsStore7[250];
			WeightsStore7[27] <= WeightsStore7[251];
			WeightsStore8[0] <= WeightsStore8[224];
			WeightsStore8[1] <= WeightsStore8[225];
			WeightsStore8[2] <= WeightsStore8[226];
			WeightsStore8[3] <= WeightsStore8[227];
			WeightsStore8[4] <= WeightsStore8[228];
			WeightsStore8[5] <= WeightsStore8[229];
			WeightsStore8[6] <= WeightsStore8[230];
			WeightsStore8[7] <= WeightsStore8[231];
			WeightsStore8[8] <= WeightsStore8[232];
			WeightsStore8[9] <= WeightsStore8[233];
			WeightsStore8[10] <= WeightsStore8[234];
			WeightsStore8[11] <= WeightsStore8[235];
			WeightsStore8[12] <= WeightsStore8[236];
			WeightsStore8[13] <= WeightsStore8[237];
			WeightsStore8[14] <= WeightsStore8[238];
			WeightsStore8[15] <= WeightsStore8[239];
			WeightsStore8[16] <= WeightsStore8[240];
			WeightsStore8[17] <= WeightsStore8[241];
			WeightsStore8[18] <= WeightsStore8[242];
			WeightsStore8[19] <= WeightsStore8[243];
			WeightsStore8[20] <= WeightsStore8[244];
			WeightsStore8[21] <= WeightsStore8[245];
			WeightsStore8[22] <= WeightsStore8[246];
			WeightsStore8[23] <= WeightsStore8[247];
			WeightsStore8[24] <= WeightsStore8[248];
			WeightsStore8[25] <= WeightsStore8[249];
			WeightsStore8[26] <= WeightsStore8[250];
			WeightsStore8[27] <= WeightsStore8[251];
			WeightsStore9[0] <= WeightsStore9[224];
			WeightsStore9[1] <= WeightsStore9[225];
			WeightsStore9[2] <= WeightsStore9[226];
			WeightsStore9[3] <= WeightsStore9[227];
			WeightsStore9[4] <= WeightsStore9[228];
			WeightsStore9[5] <= WeightsStore9[229];
			WeightsStore9[6] <= WeightsStore9[230];
			WeightsStore9[7] <= WeightsStore9[231];
			WeightsStore9[8] <= WeightsStore9[232];
			WeightsStore9[9] <= WeightsStore9[233];
			WeightsStore9[10] <= WeightsStore9[234];
			WeightsStore9[11] <= WeightsStore9[235];
			WeightsStore9[12] <= WeightsStore9[236];
			WeightsStore9[13] <= WeightsStore9[237];
			WeightsStore9[14] <= WeightsStore9[238];
			WeightsStore9[15] <= WeightsStore9[239];
			WeightsStore9[16] <= WeightsStore9[240];
			WeightsStore9[17] <= WeightsStore9[241];
			WeightsStore9[18] <= WeightsStore9[242];
			WeightsStore9[19] <= WeightsStore9[243];
			WeightsStore9[20] <= WeightsStore9[244];
			WeightsStore9[21] <= WeightsStore9[245];
			WeightsStore9[22] <= WeightsStore9[246];
			WeightsStore9[23] <= WeightsStore9[247];
			WeightsStore9[24] <= WeightsStore9[248];
			WeightsStore9[25] <= WeightsStore9[249];
			WeightsStore9[26] <= WeightsStore9[250];
			WeightsStore9[27] <= WeightsStore9[251];
		end else if(switchCounter == 32'd62)begin
			PixelsStore[0] <= PixelsStore[252];
			PixelsStore[1] <= PixelsStore[253];
			PixelsStore[2] <= PixelsStore[254];
			PixelsStore[3] <= PixelsStore[255];
			PixelsStore[4] <= PixelsStore[256];
			PixelsStore[5] <= PixelsStore[257];
			PixelsStore[6] <= PixelsStore[258];
			PixelsStore[7] <= PixelsStore[259];
			PixelsStore[8] <= PixelsStore[260];
			PixelsStore[9] <= PixelsStore[261];
			PixelsStore[10] <= PixelsStore[262];
			PixelsStore[11] <= PixelsStore[263];
			PixelsStore[12] <= PixelsStore[264];
			PixelsStore[13] <= PixelsStore[265];
			PixelsStore[14] <= PixelsStore[266];
			PixelsStore[15] <= PixelsStore[267];
			PixelsStore[16] <= PixelsStore[268];
			PixelsStore[17] <= PixelsStore[269];
			PixelsStore[18] <= PixelsStore[270];
			PixelsStore[19] <= PixelsStore[271];
			PixelsStore[20] <= PixelsStore[272];
			PixelsStore[21] <= PixelsStore[273];
			PixelsStore[22] <= PixelsStore[274];
			PixelsStore[23] <= PixelsStore[275];
			PixelsStore[24] <= PixelsStore[276];
			PixelsStore[25] <= PixelsStore[277];
			PixelsStore[26] <= PixelsStore[278];
			PixelsStore[27] <= PixelsStore[279];
			WeightsStore0[0] <= WeightsStore0[252];
			WeightsStore0[1] <= WeightsStore0[253];
			WeightsStore0[2] <= WeightsStore0[254];
			WeightsStore0[3] <= WeightsStore0[255];
			WeightsStore0[4] <= WeightsStore0[256];
			WeightsStore0[5] <= WeightsStore0[257];
			WeightsStore0[6] <= WeightsStore0[258];
			WeightsStore0[7] <= WeightsStore0[259];
			WeightsStore0[8] <= WeightsStore0[260];
			WeightsStore0[9] <= WeightsStore0[261];
			WeightsStore0[10] <= WeightsStore0[262];
			WeightsStore0[11] <= WeightsStore0[263];
			WeightsStore0[12] <= WeightsStore0[264];
			WeightsStore0[13] <= WeightsStore0[265];
			WeightsStore0[14] <= WeightsStore0[266];
			WeightsStore0[15] <= WeightsStore0[267];
			WeightsStore0[16] <= WeightsStore0[268];
			WeightsStore0[17] <= WeightsStore0[269];
			WeightsStore0[18] <= WeightsStore0[270];
			WeightsStore0[19] <= WeightsStore0[271];
			WeightsStore0[20] <= WeightsStore0[272];
			WeightsStore0[21] <= WeightsStore0[273];
			WeightsStore0[22] <= WeightsStore0[274];
			WeightsStore0[23] <= WeightsStore0[275];
			WeightsStore0[24] <= WeightsStore0[276];
			WeightsStore0[25] <= WeightsStore0[277];
			WeightsStore0[26] <= WeightsStore0[278];
			WeightsStore0[27] <= WeightsStore0[279];
			WeightsStore1[0] <= WeightsStore1[252];
			WeightsStore1[1] <= WeightsStore1[253];
			WeightsStore1[2] <= WeightsStore1[254];
			WeightsStore1[3] <= WeightsStore1[255];
			WeightsStore1[4] <= WeightsStore1[256];
			WeightsStore1[5] <= WeightsStore1[257];
			WeightsStore1[6] <= WeightsStore1[258];
			WeightsStore1[7] <= WeightsStore1[259];
			WeightsStore1[8] <= WeightsStore1[260];
			WeightsStore1[9] <= WeightsStore1[261];
			WeightsStore1[10] <= WeightsStore1[262];
			WeightsStore1[11] <= WeightsStore1[263];
			WeightsStore1[12] <= WeightsStore1[264];
			WeightsStore1[13] <= WeightsStore1[265];
			WeightsStore1[14] <= WeightsStore1[266];
			WeightsStore1[15] <= WeightsStore1[267];
			WeightsStore1[16] <= WeightsStore1[268];
			WeightsStore1[17] <= WeightsStore1[269];
			WeightsStore1[18] <= WeightsStore1[270];
			WeightsStore1[19] <= WeightsStore1[271];
			WeightsStore1[20] <= WeightsStore1[272];
			WeightsStore1[21] <= WeightsStore1[273];
			WeightsStore1[22] <= WeightsStore1[274];
			WeightsStore1[23] <= WeightsStore1[275];
			WeightsStore1[24] <= WeightsStore1[276];
			WeightsStore1[25] <= WeightsStore1[277];
			WeightsStore1[26] <= WeightsStore1[278];
			WeightsStore1[27] <= WeightsStore1[279];
			WeightsStore2[0] <= WeightsStore2[252];
			WeightsStore2[1] <= WeightsStore2[253];
			WeightsStore2[2] <= WeightsStore2[254];
			WeightsStore2[3] <= WeightsStore2[255];
			WeightsStore2[4] <= WeightsStore2[256];
			WeightsStore2[5] <= WeightsStore2[257];
			WeightsStore2[6] <= WeightsStore2[258];
			WeightsStore2[7] <= WeightsStore2[259];
			WeightsStore2[8] <= WeightsStore2[260];
			WeightsStore2[9] <= WeightsStore2[261];
			WeightsStore2[10] <= WeightsStore2[262];
			WeightsStore2[11] <= WeightsStore2[263];
			WeightsStore2[12] <= WeightsStore2[264];
			WeightsStore2[13] <= WeightsStore2[265];
			WeightsStore2[14] <= WeightsStore2[266];
			WeightsStore2[15] <= WeightsStore2[267];
			WeightsStore2[16] <= WeightsStore2[268];
			WeightsStore2[17] <= WeightsStore2[269];
			WeightsStore2[18] <= WeightsStore2[270];
			WeightsStore2[19] <= WeightsStore2[271];
			WeightsStore2[20] <= WeightsStore2[272];
			WeightsStore2[21] <= WeightsStore2[273];
			WeightsStore2[22] <= WeightsStore2[274];
			WeightsStore2[23] <= WeightsStore2[275];
			WeightsStore2[24] <= WeightsStore2[276];
			WeightsStore2[25] <= WeightsStore2[277];
			WeightsStore2[26] <= WeightsStore2[278];
			WeightsStore2[27] <= WeightsStore2[279];
			WeightsStore3[0] <= WeightsStore3[252];
			WeightsStore3[1] <= WeightsStore3[253];
			WeightsStore3[2] <= WeightsStore3[254];
			WeightsStore3[3] <= WeightsStore3[255];
			WeightsStore3[4] <= WeightsStore3[256];
			WeightsStore3[5] <= WeightsStore3[257];
			WeightsStore3[6] <= WeightsStore3[258];
			WeightsStore3[7] <= WeightsStore3[259];
			WeightsStore3[8] <= WeightsStore3[260];
			WeightsStore3[9] <= WeightsStore3[261];
			WeightsStore3[10] <= WeightsStore3[262];
			WeightsStore3[11] <= WeightsStore3[263];
			WeightsStore3[12] <= WeightsStore3[264];
			WeightsStore3[13] <= WeightsStore3[265];
			WeightsStore3[14] <= WeightsStore3[266];
			WeightsStore3[15] <= WeightsStore3[267];
			WeightsStore3[16] <= WeightsStore3[268];
			WeightsStore3[17] <= WeightsStore3[269];
			WeightsStore3[18] <= WeightsStore3[270];
			WeightsStore3[19] <= WeightsStore3[271];
			WeightsStore3[20] <= WeightsStore3[272];
			WeightsStore3[21] <= WeightsStore3[273];
			WeightsStore3[22] <= WeightsStore3[274];
			WeightsStore3[23] <= WeightsStore3[275];
			WeightsStore3[24] <= WeightsStore3[276];
			WeightsStore3[25] <= WeightsStore3[277];
			WeightsStore3[26] <= WeightsStore3[278];
			WeightsStore3[27] <= WeightsStore3[279];
			WeightsStore4[0] <= WeightsStore4[252];
			WeightsStore4[1] <= WeightsStore4[253];
			WeightsStore4[2] <= WeightsStore4[254];
			WeightsStore4[3] <= WeightsStore4[255];
			WeightsStore4[4] <= WeightsStore4[256];
			WeightsStore4[5] <= WeightsStore4[257];
			WeightsStore4[6] <= WeightsStore4[258];
			WeightsStore4[7] <= WeightsStore4[259];
			WeightsStore4[8] <= WeightsStore4[260];
			WeightsStore4[9] <= WeightsStore4[261];
			WeightsStore4[10] <= WeightsStore4[262];
			WeightsStore4[11] <= WeightsStore4[263];
			WeightsStore4[12] <= WeightsStore4[264];
			WeightsStore4[13] <= WeightsStore4[265];
			WeightsStore4[14] <= WeightsStore4[266];
			WeightsStore4[15] <= WeightsStore4[267];
			WeightsStore4[16] <= WeightsStore4[268];
			WeightsStore4[17] <= WeightsStore4[269];
			WeightsStore4[18] <= WeightsStore4[270];
			WeightsStore4[19] <= WeightsStore4[271];
			WeightsStore4[20] <= WeightsStore4[272];
			WeightsStore4[21] <= WeightsStore4[273];
			WeightsStore4[22] <= WeightsStore4[274];
			WeightsStore4[23] <= WeightsStore4[275];
			WeightsStore4[24] <= WeightsStore4[276];
			WeightsStore4[25] <= WeightsStore4[277];
			WeightsStore4[26] <= WeightsStore4[278];
			WeightsStore4[27] <= WeightsStore4[279];
			WeightsStore5[0] <= WeightsStore5[252];
			WeightsStore5[1] <= WeightsStore5[253];
			WeightsStore5[2] <= WeightsStore5[254];
			WeightsStore5[3] <= WeightsStore5[255];
			WeightsStore5[4] <= WeightsStore5[256];
			WeightsStore5[5] <= WeightsStore5[257];
			WeightsStore5[6] <= WeightsStore5[258];
			WeightsStore5[7] <= WeightsStore5[259];
			WeightsStore5[8] <= WeightsStore5[260];
			WeightsStore5[9] <= WeightsStore5[261];
			WeightsStore5[10] <= WeightsStore5[262];
			WeightsStore5[11] <= WeightsStore5[263];
			WeightsStore5[12] <= WeightsStore5[264];
			WeightsStore5[13] <= WeightsStore5[265];
			WeightsStore5[14] <= WeightsStore5[266];
			WeightsStore5[15] <= WeightsStore5[267];
			WeightsStore5[16] <= WeightsStore5[268];
			WeightsStore5[17] <= WeightsStore5[269];
			WeightsStore5[18] <= WeightsStore5[270];
			WeightsStore5[19] <= WeightsStore5[271];
			WeightsStore5[20] <= WeightsStore5[272];
			WeightsStore5[21] <= WeightsStore5[273];
			WeightsStore5[22] <= WeightsStore5[274];
			WeightsStore5[23] <= WeightsStore5[275];
			WeightsStore5[24] <= WeightsStore5[276];
			WeightsStore5[25] <= WeightsStore5[277];
			WeightsStore5[26] <= WeightsStore5[278];
			WeightsStore5[27] <= WeightsStore5[279];
			WeightsStore6[0] <= WeightsStore6[252];
			WeightsStore6[1] <= WeightsStore6[253];
			WeightsStore6[2] <= WeightsStore6[254];
			WeightsStore6[3] <= WeightsStore6[255];
			WeightsStore6[4] <= WeightsStore6[256];
			WeightsStore6[5] <= WeightsStore6[257];
			WeightsStore6[6] <= WeightsStore6[258];
			WeightsStore6[7] <= WeightsStore6[259];
			WeightsStore6[8] <= WeightsStore6[260];
			WeightsStore6[9] <= WeightsStore6[261];
			WeightsStore6[10] <= WeightsStore6[262];
			WeightsStore6[11] <= WeightsStore6[263];
			WeightsStore6[12] <= WeightsStore6[264];
			WeightsStore6[13] <= WeightsStore6[265];
			WeightsStore6[14] <= WeightsStore6[266];
			WeightsStore6[15] <= WeightsStore6[267];
			WeightsStore6[16] <= WeightsStore6[268];
			WeightsStore6[17] <= WeightsStore6[269];
			WeightsStore6[18] <= WeightsStore6[270];
			WeightsStore6[19] <= WeightsStore6[271];
			WeightsStore6[20] <= WeightsStore6[272];
			WeightsStore6[21] <= WeightsStore6[273];
			WeightsStore6[22] <= WeightsStore6[274];
			WeightsStore6[23] <= WeightsStore6[275];
			WeightsStore6[24] <= WeightsStore6[276];
			WeightsStore6[25] <= WeightsStore6[277];
			WeightsStore6[26] <= WeightsStore6[278];
			WeightsStore6[27] <= WeightsStore6[279];
			WeightsStore7[0] <= WeightsStore7[252];
			WeightsStore7[1] <= WeightsStore7[253];
			WeightsStore7[2] <= WeightsStore7[254];
			WeightsStore7[3] <= WeightsStore7[255];
			WeightsStore7[4] <= WeightsStore7[256];
			WeightsStore7[5] <= WeightsStore7[257];
			WeightsStore7[6] <= WeightsStore7[258];
			WeightsStore7[7] <= WeightsStore7[259];
			WeightsStore7[8] <= WeightsStore7[260];
			WeightsStore7[9] <= WeightsStore7[261];
			WeightsStore7[10] <= WeightsStore7[262];
			WeightsStore7[11] <= WeightsStore7[263];
			WeightsStore7[12] <= WeightsStore7[264];
			WeightsStore7[13] <= WeightsStore7[265];
			WeightsStore7[14] <= WeightsStore7[266];
			WeightsStore7[15] <= WeightsStore7[267];
			WeightsStore7[16] <= WeightsStore7[268];
			WeightsStore7[17] <= WeightsStore7[269];
			WeightsStore7[18] <= WeightsStore7[270];
			WeightsStore7[19] <= WeightsStore7[271];
			WeightsStore7[20] <= WeightsStore7[272];
			WeightsStore7[21] <= WeightsStore7[273];
			WeightsStore7[22] <= WeightsStore7[274];
			WeightsStore7[23] <= WeightsStore7[275];
			WeightsStore7[24] <= WeightsStore7[276];
			WeightsStore7[25] <= WeightsStore7[277];
			WeightsStore7[26] <= WeightsStore7[278];
			WeightsStore7[27] <= WeightsStore7[279];
			WeightsStore8[0] <= WeightsStore8[252];
			WeightsStore8[1] <= WeightsStore8[253];
			WeightsStore8[2] <= WeightsStore8[254];
			WeightsStore8[3] <= WeightsStore8[255];
			WeightsStore8[4] <= WeightsStore8[256];
			WeightsStore8[5] <= WeightsStore8[257];
			WeightsStore8[6] <= WeightsStore8[258];
			WeightsStore8[7] <= WeightsStore8[259];
			WeightsStore8[8] <= WeightsStore8[260];
			WeightsStore8[9] <= WeightsStore8[261];
			WeightsStore8[10] <= WeightsStore8[262];
			WeightsStore8[11] <= WeightsStore8[263];
			WeightsStore8[12] <= WeightsStore8[264];
			WeightsStore8[13] <= WeightsStore8[265];
			WeightsStore8[14] <= WeightsStore8[266];
			WeightsStore8[15] <= WeightsStore8[267];
			WeightsStore8[16] <= WeightsStore8[268];
			WeightsStore8[17] <= WeightsStore8[269];
			WeightsStore8[18] <= WeightsStore8[270];
			WeightsStore8[19] <= WeightsStore8[271];
			WeightsStore8[20] <= WeightsStore8[272];
			WeightsStore8[21] <= WeightsStore8[273];
			WeightsStore8[22] <= WeightsStore8[274];
			WeightsStore8[23] <= WeightsStore8[275];
			WeightsStore8[24] <= WeightsStore8[276];
			WeightsStore8[25] <= WeightsStore8[277];
			WeightsStore8[26] <= WeightsStore8[278];
			WeightsStore8[27] <= WeightsStore8[279];
			WeightsStore9[0] <= WeightsStore9[252];
			WeightsStore9[1] <= WeightsStore9[253];
			WeightsStore9[2] <= WeightsStore9[254];
			WeightsStore9[3] <= WeightsStore9[255];
			WeightsStore9[4] <= WeightsStore9[256];
			WeightsStore9[5] <= WeightsStore9[257];
			WeightsStore9[6] <= WeightsStore9[258];
			WeightsStore9[7] <= WeightsStore9[259];
			WeightsStore9[8] <= WeightsStore9[260];
			WeightsStore9[9] <= WeightsStore9[261];
			WeightsStore9[10] <= WeightsStore9[262];
			WeightsStore9[11] <= WeightsStore9[263];
			WeightsStore9[12] <= WeightsStore9[264];
			WeightsStore9[13] <= WeightsStore9[265];
			WeightsStore9[14] <= WeightsStore9[266];
			WeightsStore9[15] <= WeightsStore9[267];
			WeightsStore9[16] <= WeightsStore9[268];
			WeightsStore9[17] <= WeightsStore9[269];
			WeightsStore9[18] <= WeightsStore9[270];
			WeightsStore9[19] <= WeightsStore9[271];
			WeightsStore9[20] <= WeightsStore9[272];
			WeightsStore9[21] <= WeightsStore9[273];
			WeightsStore9[22] <= WeightsStore9[274];
			WeightsStore9[23] <= WeightsStore9[275];
			WeightsStore9[24] <= WeightsStore9[276];
			WeightsStore9[25] <= WeightsStore9[277];
			WeightsStore9[26] <= WeightsStore9[278];
			WeightsStore9[27] <= WeightsStore9[279];
		end else if(switchCounter == 32'd69)begin
			PixelsStore[0] <= PixelsStore[280];
			PixelsStore[1] <= PixelsStore[281];
			PixelsStore[2] <= PixelsStore[282];
			PixelsStore[3] <= PixelsStore[283];
			PixelsStore[4] <= PixelsStore[284];
			PixelsStore[5] <= PixelsStore[285];
			PixelsStore[6] <= PixelsStore[286];
			PixelsStore[7] <= PixelsStore[287];
			PixelsStore[8] <= PixelsStore[288];
			PixelsStore[9] <= PixelsStore[289];
			PixelsStore[10] <= PixelsStore[290];
			PixelsStore[11] <= PixelsStore[291];
			PixelsStore[12] <= PixelsStore[292];
			PixelsStore[13] <= PixelsStore[293];
			PixelsStore[14] <= PixelsStore[294];
			PixelsStore[15] <= PixelsStore[295];
			PixelsStore[16] <= PixelsStore[296];
			PixelsStore[17] <= PixelsStore[297];
			PixelsStore[18] <= PixelsStore[298];
			PixelsStore[19] <= PixelsStore[299];
			PixelsStore[20] <= PixelsStore[300];
			PixelsStore[21] <= PixelsStore[301];
			PixelsStore[22] <= PixelsStore[302];
			PixelsStore[23] <= PixelsStore[303];
			PixelsStore[24] <= PixelsStore[304];
			PixelsStore[25] <= PixelsStore[305];
			PixelsStore[26] <= PixelsStore[306];
			PixelsStore[27] <= PixelsStore[307];
			WeightsStore0[0] <= WeightsStore0[280];
			WeightsStore0[1] <= WeightsStore0[281];
			WeightsStore0[2] <= WeightsStore0[282];
			WeightsStore0[3] <= WeightsStore0[283];
			WeightsStore0[4] <= WeightsStore0[284];
			WeightsStore0[5] <= WeightsStore0[285];
			WeightsStore0[6] <= WeightsStore0[286];
			WeightsStore0[7] <= WeightsStore0[287];
			WeightsStore0[8] <= WeightsStore0[288];
			WeightsStore0[9] <= WeightsStore0[289];
			WeightsStore0[10] <= WeightsStore0[290];
			WeightsStore0[11] <= WeightsStore0[291];
			WeightsStore0[12] <= WeightsStore0[292];
			WeightsStore0[13] <= WeightsStore0[293];
			WeightsStore0[14] <= WeightsStore0[294];
			WeightsStore0[15] <= WeightsStore0[295];
			WeightsStore0[16] <= WeightsStore0[296];
			WeightsStore0[17] <= WeightsStore0[297];
			WeightsStore0[18] <= WeightsStore0[298];
			WeightsStore0[19] <= WeightsStore0[299];
			WeightsStore0[20] <= WeightsStore0[300];
			WeightsStore0[21] <= WeightsStore0[301];
			WeightsStore0[22] <= WeightsStore0[302];
			WeightsStore0[23] <= WeightsStore0[303];
			WeightsStore0[24] <= WeightsStore0[304];
			WeightsStore0[25] <= WeightsStore0[305];
			WeightsStore0[26] <= WeightsStore0[306];
			WeightsStore0[27] <= WeightsStore0[307];
			WeightsStore1[0] <= WeightsStore1[280];
			WeightsStore1[1] <= WeightsStore1[281];
			WeightsStore1[2] <= WeightsStore1[282];
			WeightsStore1[3] <= WeightsStore1[283];
			WeightsStore1[4] <= WeightsStore1[284];
			WeightsStore1[5] <= WeightsStore1[285];
			WeightsStore1[6] <= WeightsStore1[286];
			WeightsStore1[7] <= WeightsStore1[287];
			WeightsStore1[8] <= WeightsStore1[288];
			WeightsStore1[9] <= WeightsStore1[289];
			WeightsStore1[10] <= WeightsStore1[290];
			WeightsStore1[11] <= WeightsStore1[291];
			WeightsStore1[12] <= WeightsStore1[292];
			WeightsStore1[13] <= WeightsStore1[293];
			WeightsStore1[14] <= WeightsStore1[294];
			WeightsStore1[15] <= WeightsStore1[295];
			WeightsStore1[16] <= WeightsStore1[296];
			WeightsStore1[17] <= WeightsStore1[297];
			WeightsStore1[18] <= WeightsStore1[298];
			WeightsStore1[19] <= WeightsStore1[299];
			WeightsStore1[20] <= WeightsStore1[300];
			WeightsStore1[21] <= WeightsStore1[301];
			WeightsStore1[22] <= WeightsStore1[302];
			WeightsStore1[23] <= WeightsStore1[303];
			WeightsStore1[24] <= WeightsStore1[304];
			WeightsStore1[25] <= WeightsStore1[305];
			WeightsStore1[26] <= WeightsStore1[306];
			WeightsStore1[27] <= WeightsStore1[307];
			WeightsStore2[0] <= WeightsStore2[280];
			WeightsStore2[1] <= WeightsStore2[281];
			WeightsStore2[2] <= WeightsStore2[282];
			WeightsStore2[3] <= WeightsStore2[283];
			WeightsStore2[4] <= WeightsStore2[284];
			WeightsStore2[5] <= WeightsStore2[285];
			WeightsStore2[6] <= WeightsStore2[286];
			WeightsStore2[7] <= WeightsStore2[287];
			WeightsStore2[8] <= WeightsStore2[288];
			WeightsStore2[9] <= WeightsStore2[289];
			WeightsStore2[10] <= WeightsStore2[290];
			WeightsStore2[11] <= WeightsStore2[291];
			WeightsStore2[12] <= WeightsStore2[292];
			WeightsStore2[13] <= WeightsStore2[293];
			WeightsStore2[14] <= WeightsStore2[294];
			WeightsStore2[15] <= WeightsStore2[295];
			WeightsStore2[16] <= WeightsStore2[296];
			WeightsStore2[17] <= WeightsStore2[297];
			WeightsStore2[18] <= WeightsStore2[298];
			WeightsStore2[19] <= WeightsStore2[299];
			WeightsStore2[20] <= WeightsStore2[300];
			WeightsStore2[21] <= WeightsStore2[301];
			WeightsStore2[22] <= WeightsStore2[302];
			WeightsStore2[23] <= WeightsStore2[303];
			WeightsStore2[24] <= WeightsStore2[304];
			WeightsStore2[25] <= WeightsStore2[305];
			WeightsStore2[26] <= WeightsStore2[306];
			WeightsStore2[27] <= WeightsStore2[307];
			WeightsStore3[0] <= WeightsStore3[280];
			WeightsStore3[1] <= WeightsStore3[281];
			WeightsStore3[2] <= WeightsStore3[282];
			WeightsStore3[3] <= WeightsStore3[283];
			WeightsStore3[4] <= WeightsStore3[284];
			WeightsStore3[5] <= WeightsStore3[285];
			WeightsStore3[6] <= WeightsStore3[286];
			WeightsStore3[7] <= WeightsStore3[287];
			WeightsStore3[8] <= WeightsStore3[288];
			WeightsStore3[9] <= WeightsStore3[289];
			WeightsStore3[10] <= WeightsStore3[290];
			WeightsStore3[11] <= WeightsStore3[291];
			WeightsStore3[12] <= WeightsStore3[292];
			WeightsStore3[13] <= WeightsStore3[293];
			WeightsStore3[14] <= WeightsStore3[294];
			WeightsStore3[15] <= WeightsStore3[295];
			WeightsStore3[16] <= WeightsStore3[296];
			WeightsStore3[17] <= WeightsStore3[297];
			WeightsStore3[18] <= WeightsStore3[298];
			WeightsStore3[19] <= WeightsStore3[299];
			WeightsStore3[20] <= WeightsStore3[300];
			WeightsStore3[21] <= WeightsStore3[301];
			WeightsStore3[22] <= WeightsStore3[302];
			WeightsStore3[23] <= WeightsStore3[303];
			WeightsStore3[24] <= WeightsStore3[304];
			WeightsStore3[25] <= WeightsStore3[305];
			WeightsStore3[26] <= WeightsStore3[306];
			WeightsStore3[27] <= WeightsStore3[307];
			WeightsStore4[0] <= WeightsStore4[280];
			WeightsStore4[1] <= WeightsStore4[281];
			WeightsStore4[2] <= WeightsStore4[282];
			WeightsStore4[3] <= WeightsStore4[283];
			WeightsStore4[4] <= WeightsStore4[284];
			WeightsStore4[5] <= WeightsStore4[285];
			WeightsStore4[6] <= WeightsStore4[286];
			WeightsStore4[7] <= WeightsStore4[287];
			WeightsStore4[8] <= WeightsStore4[288];
			WeightsStore4[9] <= WeightsStore4[289];
			WeightsStore4[10] <= WeightsStore4[290];
			WeightsStore4[11] <= WeightsStore4[291];
			WeightsStore4[12] <= WeightsStore4[292];
			WeightsStore4[13] <= WeightsStore4[293];
			WeightsStore4[14] <= WeightsStore4[294];
			WeightsStore4[15] <= WeightsStore4[295];
			WeightsStore4[16] <= WeightsStore4[296];
			WeightsStore4[17] <= WeightsStore4[297];
			WeightsStore4[18] <= WeightsStore4[298];
			WeightsStore4[19] <= WeightsStore4[299];
			WeightsStore4[20] <= WeightsStore4[300];
			WeightsStore4[21] <= WeightsStore4[301];
			WeightsStore4[22] <= WeightsStore4[302];
			WeightsStore4[23] <= WeightsStore4[303];
			WeightsStore4[24] <= WeightsStore4[304];
			WeightsStore4[25] <= WeightsStore4[305];
			WeightsStore4[26] <= WeightsStore4[306];
			WeightsStore4[27] <= WeightsStore4[307];
			WeightsStore5[0] <= WeightsStore5[280];
			WeightsStore5[1] <= WeightsStore5[281];
			WeightsStore5[2] <= WeightsStore5[282];
			WeightsStore5[3] <= WeightsStore5[283];
			WeightsStore5[4] <= WeightsStore5[284];
			WeightsStore5[5] <= WeightsStore5[285];
			WeightsStore5[6] <= WeightsStore5[286];
			WeightsStore5[7] <= WeightsStore5[287];
			WeightsStore5[8] <= WeightsStore5[288];
			WeightsStore5[9] <= WeightsStore5[289];
			WeightsStore5[10] <= WeightsStore5[290];
			WeightsStore5[11] <= WeightsStore5[291];
			WeightsStore5[12] <= WeightsStore5[292];
			WeightsStore5[13] <= WeightsStore5[293];
			WeightsStore5[14] <= WeightsStore5[294];
			WeightsStore5[15] <= WeightsStore5[295];
			WeightsStore5[16] <= WeightsStore5[296];
			WeightsStore5[17] <= WeightsStore5[297];
			WeightsStore5[18] <= WeightsStore5[298];
			WeightsStore5[19] <= WeightsStore5[299];
			WeightsStore5[20] <= WeightsStore5[300];
			WeightsStore5[21] <= WeightsStore5[301];
			WeightsStore5[22] <= WeightsStore5[302];
			WeightsStore5[23] <= WeightsStore5[303];
			WeightsStore5[24] <= WeightsStore5[304];
			WeightsStore5[25] <= WeightsStore5[305];
			WeightsStore5[26] <= WeightsStore5[306];
			WeightsStore5[27] <= WeightsStore5[307];
			WeightsStore6[0] <= WeightsStore6[280];
			WeightsStore6[1] <= WeightsStore6[281];
			WeightsStore6[2] <= WeightsStore6[282];
			WeightsStore6[3] <= WeightsStore6[283];
			WeightsStore6[4] <= WeightsStore6[284];
			WeightsStore6[5] <= WeightsStore6[285];
			WeightsStore6[6] <= WeightsStore6[286];
			WeightsStore6[7] <= WeightsStore6[287];
			WeightsStore6[8] <= WeightsStore6[288];
			WeightsStore6[9] <= WeightsStore6[289];
			WeightsStore6[10] <= WeightsStore6[290];
			WeightsStore6[11] <= WeightsStore6[291];
			WeightsStore6[12] <= WeightsStore6[292];
			WeightsStore6[13] <= WeightsStore6[293];
			WeightsStore6[14] <= WeightsStore6[294];
			WeightsStore6[15] <= WeightsStore6[295];
			WeightsStore6[16] <= WeightsStore6[296];
			WeightsStore6[17] <= WeightsStore6[297];
			WeightsStore6[18] <= WeightsStore6[298];
			WeightsStore6[19] <= WeightsStore6[299];
			WeightsStore6[20] <= WeightsStore6[300];
			WeightsStore6[21] <= WeightsStore6[301];
			WeightsStore6[22] <= WeightsStore6[302];
			WeightsStore6[23] <= WeightsStore6[303];
			WeightsStore6[24] <= WeightsStore6[304];
			WeightsStore6[25] <= WeightsStore6[305];
			WeightsStore6[26] <= WeightsStore6[306];
			WeightsStore6[27] <= WeightsStore6[307];
			WeightsStore7[0] <= WeightsStore7[280];
			WeightsStore7[1] <= WeightsStore7[281];
			WeightsStore7[2] <= WeightsStore7[282];
			WeightsStore7[3] <= WeightsStore7[283];
			WeightsStore7[4] <= WeightsStore7[284];
			WeightsStore7[5] <= WeightsStore7[285];
			WeightsStore7[6] <= WeightsStore7[286];
			WeightsStore7[7] <= WeightsStore7[287];
			WeightsStore7[8] <= WeightsStore7[288];
			WeightsStore7[9] <= WeightsStore7[289];
			WeightsStore7[10] <= WeightsStore7[290];
			WeightsStore7[11] <= WeightsStore7[291];
			WeightsStore7[12] <= WeightsStore7[292];
			WeightsStore7[13] <= WeightsStore7[293];
			WeightsStore7[14] <= WeightsStore7[294];
			WeightsStore7[15] <= WeightsStore7[295];
			WeightsStore7[16] <= WeightsStore7[296];
			WeightsStore7[17] <= WeightsStore7[297];
			WeightsStore7[18] <= WeightsStore7[298];
			WeightsStore7[19] <= WeightsStore7[299];
			WeightsStore7[20] <= WeightsStore7[300];
			WeightsStore7[21] <= WeightsStore7[301];
			WeightsStore7[22] <= WeightsStore7[302];
			WeightsStore7[23] <= WeightsStore7[303];
			WeightsStore7[24] <= WeightsStore7[304];
			WeightsStore7[25] <= WeightsStore7[305];
			WeightsStore7[26] <= WeightsStore7[306];
			WeightsStore7[27] <= WeightsStore7[307];
			WeightsStore8[0] <= WeightsStore8[280];
			WeightsStore8[1] <= WeightsStore8[281];
			WeightsStore8[2] <= WeightsStore8[282];
			WeightsStore8[3] <= WeightsStore8[283];
			WeightsStore8[4] <= WeightsStore8[284];
			WeightsStore8[5] <= WeightsStore8[285];
			WeightsStore8[6] <= WeightsStore8[286];
			WeightsStore8[7] <= WeightsStore8[287];
			WeightsStore8[8] <= WeightsStore8[288];
			WeightsStore8[9] <= WeightsStore8[289];
			WeightsStore8[10] <= WeightsStore8[290];
			WeightsStore8[11] <= WeightsStore8[291];
			WeightsStore8[12] <= WeightsStore8[292];
			WeightsStore8[13] <= WeightsStore8[293];
			WeightsStore8[14] <= WeightsStore8[294];
			WeightsStore8[15] <= WeightsStore8[295];
			WeightsStore8[16] <= WeightsStore8[296];
			WeightsStore8[17] <= WeightsStore8[297];
			WeightsStore8[18] <= WeightsStore8[298];
			WeightsStore8[19] <= WeightsStore8[299];
			WeightsStore8[20] <= WeightsStore8[300];
			WeightsStore8[21] <= WeightsStore8[301];
			WeightsStore8[22] <= WeightsStore8[302];
			WeightsStore8[23] <= WeightsStore8[303];
			WeightsStore8[24] <= WeightsStore8[304];
			WeightsStore8[25] <= WeightsStore8[305];
			WeightsStore8[26] <= WeightsStore8[306];
			WeightsStore8[27] <= WeightsStore8[307];
			WeightsStore9[0] <= WeightsStore9[280];
			WeightsStore9[1] <= WeightsStore9[281];
			WeightsStore9[2] <= WeightsStore9[282];
			WeightsStore9[3] <= WeightsStore9[283];
			WeightsStore9[4] <= WeightsStore9[284];
			WeightsStore9[5] <= WeightsStore9[285];
			WeightsStore9[6] <= WeightsStore9[286];
			WeightsStore9[7] <= WeightsStore9[287];
			WeightsStore9[8] <= WeightsStore9[288];
			WeightsStore9[9] <= WeightsStore9[289];
			WeightsStore9[10] <= WeightsStore9[290];
			WeightsStore9[11] <= WeightsStore9[291];
			WeightsStore9[12] <= WeightsStore9[292];
			WeightsStore9[13] <= WeightsStore9[293];
			WeightsStore9[14] <= WeightsStore9[294];
			WeightsStore9[15] <= WeightsStore9[295];
			WeightsStore9[16] <= WeightsStore9[296];
			WeightsStore9[17] <= WeightsStore9[297];
			WeightsStore9[18] <= WeightsStore9[298];
			WeightsStore9[19] <= WeightsStore9[299];
			WeightsStore9[20] <= WeightsStore9[300];
			WeightsStore9[21] <= WeightsStore9[301];
			WeightsStore9[22] <= WeightsStore9[302];
			WeightsStore9[23] <= WeightsStore9[303];
			WeightsStore9[24] <= WeightsStore9[304];
			WeightsStore9[25] <= WeightsStore9[305];
			WeightsStore9[26] <= WeightsStore9[306];
			WeightsStore9[27] <= WeightsStore9[307];
		end else if(switchCounter == 32'd76)begin
			PixelsStore[0] <= PixelsStore[308];
			PixelsStore[1] <= PixelsStore[309];
			PixelsStore[2] <= PixelsStore[310];
			PixelsStore[3] <= PixelsStore[311];
			PixelsStore[4] <= PixelsStore[312];
			PixelsStore[5] <= PixelsStore[313];
			PixelsStore[6] <= PixelsStore[314];
			PixelsStore[7] <= PixelsStore[315];
			PixelsStore[8] <= PixelsStore[316];
			PixelsStore[9] <= PixelsStore[317];
			PixelsStore[10] <= PixelsStore[318];
			PixelsStore[11] <= PixelsStore[319];
			PixelsStore[12] <= PixelsStore[320];
			PixelsStore[13] <= PixelsStore[321];
			PixelsStore[14] <= PixelsStore[322];
			PixelsStore[15] <= PixelsStore[323];
			PixelsStore[16] <= PixelsStore[324];
			PixelsStore[17] <= PixelsStore[325];
			PixelsStore[18] <= PixelsStore[326];
			PixelsStore[19] <= PixelsStore[327];
			PixelsStore[20] <= PixelsStore[328];
			PixelsStore[21] <= PixelsStore[329];
			PixelsStore[22] <= PixelsStore[330];
			PixelsStore[23] <= PixelsStore[331];
			PixelsStore[24] <= PixelsStore[332];
			PixelsStore[25] <= PixelsStore[333];
			PixelsStore[26] <= PixelsStore[334];
			PixelsStore[27] <= PixelsStore[335];
			WeightsStore0[0] <= WeightsStore0[308];
			WeightsStore0[1] <= WeightsStore0[309];
			WeightsStore0[2] <= WeightsStore0[310];
			WeightsStore0[3] <= WeightsStore0[311];
			WeightsStore0[4] <= WeightsStore0[312];
			WeightsStore0[5] <= WeightsStore0[313];
			WeightsStore0[6] <= WeightsStore0[314];
			WeightsStore0[7] <= WeightsStore0[315];
			WeightsStore0[8] <= WeightsStore0[316];
			WeightsStore0[9] <= WeightsStore0[317];
			WeightsStore0[10] <= WeightsStore0[318];
			WeightsStore0[11] <= WeightsStore0[319];
			WeightsStore0[12] <= WeightsStore0[320];
			WeightsStore0[13] <= WeightsStore0[321];
			WeightsStore0[14] <= WeightsStore0[322];
			WeightsStore0[15] <= WeightsStore0[323];
			WeightsStore0[16] <= WeightsStore0[324];
			WeightsStore0[17] <= WeightsStore0[325];
			WeightsStore0[18] <= WeightsStore0[326];
			WeightsStore0[19] <= WeightsStore0[327];
			WeightsStore0[20] <= WeightsStore0[328];
			WeightsStore0[21] <= WeightsStore0[329];
			WeightsStore0[22] <= WeightsStore0[330];
			WeightsStore0[23] <= WeightsStore0[331];
			WeightsStore0[24] <= WeightsStore0[332];
			WeightsStore0[25] <= WeightsStore0[333];
			WeightsStore0[26] <= WeightsStore0[334];
			WeightsStore0[27] <= WeightsStore0[335];
			WeightsStore1[0] <= WeightsStore1[308];
			WeightsStore1[1] <= WeightsStore1[309];
			WeightsStore1[2] <= WeightsStore1[310];
			WeightsStore1[3] <= WeightsStore1[311];
			WeightsStore1[4] <= WeightsStore1[312];
			WeightsStore1[5] <= WeightsStore1[313];
			WeightsStore1[6] <= WeightsStore1[314];
			WeightsStore1[7] <= WeightsStore1[315];
			WeightsStore1[8] <= WeightsStore1[316];
			WeightsStore1[9] <= WeightsStore1[317];
			WeightsStore1[10] <= WeightsStore1[318];
			WeightsStore1[11] <= WeightsStore1[319];
			WeightsStore1[12] <= WeightsStore1[320];
			WeightsStore1[13] <= WeightsStore1[321];
			WeightsStore1[14] <= WeightsStore1[322];
			WeightsStore1[15] <= WeightsStore1[323];
			WeightsStore1[16] <= WeightsStore1[324];
			WeightsStore1[17] <= WeightsStore1[325];
			WeightsStore1[18] <= WeightsStore1[326];
			WeightsStore1[19] <= WeightsStore1[327];
			WeightsStore1[20] <= WeightsStore1[328];
			WeightsStore1[21] <= WeightsStore1[329];
			WeightsStore1[22] <= WeightsStore1[330];
			WeightsStore1[23] <= WeightsStore1[331];
			WeightsStore1[24] <= WeightsStore1[332];
			WeightsStore1[25] <= WeightsStore1[333];
			WeightsStore1[26] <= WeightsStore1[334];
			WeightsStore1[27] <= WeightsStore1[335];
			WeightsStore2[0] <= WeightsStore2[308];
			WeightsStore2[1] <= WeightsStore2[309];
			WeightsStore2[2] <= WeightsStore2[310];
			WeightsStore2[3] <= WeightsStore2[311];
			WeightsStore2[4] <= WeightsStore2[312];
			WeightsStore2[5] <= WeightsStore2[313];
			WeightsStore2[6] <= WeightsStore2[314];
			WeightsStore2[7] <= WeightsStore2[315];
			WeightsStore2[8] <= WeightsStore2[316];
			WeightsStore2[9] <= WeightsStore2[317];
			WeightsStore2[10] <= WeightsStore2[318];
			WeightsStore2[11] <= WeightsStore2[319];
			WeightsStore2[12] <= WeightsStore2[320];
			WeightsStore2[13] <= WeightsStore2[321];
			WeightsStore2[14] <= WeightsStore2[322];
			WeightsStore2[15] <= WeightsStore2[323];
			WeightsStore2[16] <= WeightsStore2[324];
			WeightsStore2[17] <= WeightsStore2[325];
			WeightsStore2[18] <= WeightsStore2[326];
			WeightsStore2[19] <= WeightsStore2[327];
			WeightsStore2[20] <= WeightsStore2[328];
			WeightsStore2[21] <= WeightsStore2[329];
			WeightsStore2[22] <= WeightsStore2[330];
			WeightsStore2[23] <= WeightsStore2[331];
			WeightsStore2[24] <= WeightsStore2[332];
			WeightsStore2[25] <= WeightsStore2[333];
			WeightsStore2[26] <= WeightsStore2[334];
			WeightsStore2[27] <= WeightsStore2[335];
			WeightsStore3[0] <= WeightsStore3[308];
			WeightsStore3[1] <= WeightsStore3[309];
			WeightsStore3[2] <= WeightsStore3[310];
			WeightsStore3[3] <= WeightsStore3[311];
			WeightsStore3[4] <= WeightsStore3[312];
			WeightsStore3[5] <= WeightsStore3[313];
			WeightsStore3[6] <= WeightsStore3[314];
			WeightsStore3[7] <= WeightsStore3[315];
			WeightsStore3[8] <= WeightsStore3[316];
			WeightsStore3[9] <= WeightsStore3[317];
			WeightsStore3[10] <= WeightsStore3[318];
			WeightsStore3[11] <= WeightsStore3[319];
			WeightsStore3[12] <= WeightsStore3[320];
			WeightsStore3[13] <= WeightsStore3[321];
			WeightsStore3[14] <= WeightsStore3[322];
			WeightsStore3[15] <= WeightsStore3[323];
			WeightsStore3[16] <= WeightsStore3[324];
			WeightsStore3[17] <= WeightsStore3[325];
			WeightsStore3[18] <= WeightsStore3[326];
			WeightsStore3[19] <= WeightsStore3[327];
			WeightsStore3[20] <= WeightsStore3[328];
			WeightsStore3[21] <= WeightsStore3[329];
			WeightsStore3[22] <= WeightsStore3[330];
			WeightsStore3[23] <= WeightsStore3[331];
			WeightsStore3[24] <= WeightsStore3[332];
			WeightsStore3[25] <= WeightsStore3[333];
			WeightsStore3[26] <= WeightsStore3[334];
			WeightsStore3[27] <= WeightsStore3[335];
			WeightsStore4[0] <= WeightsStore4[308];
			WeightsStore4[1] <= WeightsStore4[309];
			WeightsStore4[2] <= WeightsStore4[310];
			WeightsStore4[3] <= WeightsStore4[311];
			WeightsStore4[4] <= WeightsStore4[312];
			WeightsStore4[5] <= WeightsStore4[313];
			WeightsStore4[6] <= WeightsStore4[314];
			WeightsStore4[7] <= WeightsStore4[315];
			WeightsStore4[8] <= WeightsStore4[316];
			WeightsStore4[9] <= WeightsStore4[317];
			WeightsStore4[10] <= WeightsStore4[318];
			WeightsStore4[11] <= WeightsStore4[319];
			WeightsStore4[12] <= WeightsStore4[320];
			WeightsStore4[13] <= WeightsStore4[321];
			WeightsStore4[14] <= WeightsStore4[322];
			WeightsStore4[15] <= WeightsStore4[323];
			WeightsStore4[16] <= WeightsStore4[324];
			WeightsStore4[17] <= WeightsStore4[325];
			WeightsStore4[18] <= WeightsStore4[326];
			WeightsStore4[19] <= WeightsStore4[327];
			WeightsStore4[20] <= WeightsStore4[328];
			WeightsStore4[21] <= WeightsStore4[329];
			WeightsStore4[22] <= WeightsStore4[330];
			WeightsStore4[23] <= WeightsStore4[331];
			WeightsStore4[24] <= WeightsStore4[332];
			WeightsStore4[25] <= WeightsStore4[333];
			WeightsStore4[26] <= WeightsStore4[334];
			WeightsStore4[27] <= WeightsStore4[335];
			WeightsStore5[0] <= WeightsStore5[308];
			WeightsStore5[1] <= WeightsStore5[309];
			WeightsStore5[2] <= WeightsStore5[310];
			WeightsStore5[3] <= WeightsStore5[311];
			WeightsStore5[4] <= WeightsStore5[312];
			WeightsStore5[5] <= WeightsStore5[313];
			WeightsStore5[6] <= WeightsStore5[314];
			WeightsStore5[7] <= WeightsStore5[315];
			WeightsStore5[8] <= WeightsStore5[316];
			WeightsStore5[9] <= WeightsStore5[317];
			WeightsStore5[10] <= WeightsStore5[318];
			WeightsStore5[11] <= WeightsStore5[319];
			WeightsStore5[12] <= WeightsStore5[320];
			WeightsStore5[13] <= WeightsStore5[321];
			WeightsStore5[14] <= WeightsStore5[322];
			WeightsStore5[15] <= WeightsStore5[323];
			WeightsStore5[16] <= WeightsStore5[324];
			WeightsStore5[17] <= WeightsStore5[325];
			WeightsStore5[18] <= WeightsStore5[326];
			WeightsStore5[19] <= WeightsStore5[327];
			WeightsStore5[20] <= WeightsStore5[328];
			WeightsStore5[21] <= WeightsStore5[329];
			WeightsStore5[22] <= WeightsStore5[330];
			WeightsStore5[23] <= WeightsStore5[331];
			WeightsStore5[24] <= WeightsStore5[332];
			WeightsStore5[25] <= WeightsStore5[333];
			WeightsStore5[26] <= WeightsStore5[334];
			WeightsStore5[27] <= WeightsStore5[335];
			WeightsStore6[0] <= WeightsStore6[308];
			WeightsStore6[1] <= WeightsStore6[309];
			WeightsStore6[2] <= WeightsStore6[310];
			WeightsStore6[3] <= WeightsStore6[311];
			WeightsStore6[4] <= WeightsStore6[312];
			WeightsStore6[5] <= WeightsStore6[313];
			WeightsStore6[6] <= WeightsStore6[314];
			WeightsStore6[7] <= WeightsStore6[315];
			WeightsStore6[8] <= WeightsStore6[316];
			WeightsStore6[9] <= WeightsStore6[317];
			WeightsStore6[10] <= WeightsStore6[318];
			WeightsStore6[11] <= WeightsStore6[319];
			WeightsStore6[12] <= WeightsStore6[320];
			WeightsStore6[13] <= WeightsStore6[321];
			WeightsStore6[14] <= WeightsStore6[322];
			WeightsStore6[15] <= WeightsStore6[323];
			WeightsStore6[16] <= WeightsStore6[324];
			WeightsStore6[17] <= WeightsStore6[325];
			WeightsStore6[18] <= WeightsStore6[326];
			WeightsStore6[19] <= WeightsStore6[327];
			WeightsStore6[20] <= WeightsStore6[328];
			WeightsStore6[21] <= WeightsStore6[329];
			WeightsStore6[22] <= WeightsStore6[330];
			WeightsStore6[23] <= WeightsStore6[331];
			WeightsStore6[24] <= WeightsStore6[332];
			WeightsStore6[25] <= WeightsStore6[333];
			WeightsStore6[26] <= WeightsStore6[334];
			WeightsStore6[27] <= WeightsStore6[335];
			WeightsStore7[0] <= WeightsStore7[308];
			WeightsStore7[1] <= WeightsStore7[309];
			WeightsStore7[2] <= WeightsStore7[310];
			WeightsStore7[3] <= WeightsStore7[311];
			WeightsStore7[4] <= WeightsStore7[312];
			WeightsStore7[5] <= WeightsStore7[313];
			WeightsStore7[6] <= WeightsStore7[314];
			WeightsStore7[7] <= WeightsStore7[315];
			WeightsStore7[8] <= WeightsStore7[316];
			WeightsStore7[9] <= WeightsStore7[317];
			WeightsStore7[10] <= WeightsStore7[318];
			WeightsStore7[11] <= WeightsStore7[319];
			WeightsStore7[12] <= WeightsStore7[320];
			WeightsStore7[13] <= WeightsStore7[321];
			WeightsStore7[14] <= WeightsStore7[322];
			WeightsStore7[15] <= WeightsStore7[323];
			WeightsStore7[16] <= WeightsStore7[324];
			WeightsStore7[17] <= WeightsStore7[325];
			WeightsStore7[18] <= WeightsStore7[326];
			WeightsStore7[19] <= WeightsStore7[327];
			WeightsStore7[20] <= WeightsStore7[328];
			WeightsStore7[21] <= WeightsStore7[329];
			WeightsStore7[22] <= WeightsStore7[330];
			WeightsStore7[23] <= WeightsStore7[331];
			WeightsStore7[24] <= WeightsStore7[332];
			WeightsStore7[25] <= WeightsStore7[333];
			WeightsStore7[26] <= WeightsStore7[334];
			WeightsStore7[27] <= WeightsStore7[335];
			WeightsStore8[0] <= WeightsStore8[308];
			WeightsStore8[1] <= WeightsStore8[309];
			WeightsStore8[2] <= WeightsStore8[310];
			WeightsStore8[3] <= WeightsStore8[311];
			WeightsStore8[4] <= WeightsStore8[312];
			WeightsStore8[5] <= WeightsStore8[313];
			WeightsStore8[6] <= WeightsStore8[314];
			WeightsStore8[7] <= WeightsStore8[315];
			WeightsStore8[8] <= WeightsStore8[316];
			WeightsStore8[9] <= WeightsStore8[317];
			WeightsStore8[10] <= WeightsStore8[318];
			WeightsStore8[11] <= WeightsStore8[319];
			WeightsStore8[12] <= WeightsStore8[320];
			WeightsStore8[13] <= WeightsStore8[321];
			WeightsStore8[14] <= WeightsStore8[322];
			WeightsStore8[15] <= WeightsStore8[323];
			WeightsStore8[16] <= WeightsStore8[324];
			WeightsStore8[17] <= WeightsStore8[325];
			WeightsStore8[18] <= WeightsStore8[326];
			WeightsStore8[19] <= WeightsStore8[327];
			WeightsStore8[20] <= WeightsStore8[328];
			WeightsStore8[21] <= WeightsStore8[329];
			WeightsStore8[22] <= WeightsStore8[330];
			WeightsStore8[23] <= WeightsStore8[331];
			WeightsStore8[24] <= WeightsStore8[332];
			WeightsStore8[25] <= WeightsStore8[333];
			WeightsStore8[26] <= WeightsStore8[334];
			WeightsStore8[27] <= WeightsStore8[335];
			WeightsStore9[0] <= WeightsStore9[308];
			WeightsStore9[1] <= WeightsStore9[309];
			WeightsStore9[2] <= WeightsStore9[310];
			WeightsStore9[3] <= WeightsStore9[311];
			WeightsStore9[4] <= WeightsStore9[312];
			WeightsStore9[5] <= WeightsStore9[313];
			WeightsStore9[6] <= WeightsStore9[314];
			WeightsStore9[7] <= WeightsStore9[315];
			WeightsStore9[8] <= WeightsStore9[316];
			WeightsStore9[9] <= WeightsStore9[317];
			WeightsStore9[10] <= WeightsStore9[318];
			WeightsStore9[11] <= WeightsStore9[319];
			WeightsStore9[12] <= WeightsStore9[320];
			WeightsStore9[13] <= WeightsStore9[321];
			WeightsStore9[14] <= WeightsStore9[322];
			WeightsStore9[15] <= WeightsStore9[323];
			WeightsStore9[16] <= WeightsStore9[324];
			WeightsStore9[17] <= WeightsStore9[325];
			WeightsStore9[18] <= WeightsStore9[326];
			WeightsStore9[19] <= WeightsStore9[327];
			WeightsStore9[20] <= WeightsStore9[328];
			WeightsStore9[21] <= WeightsStore9[329];
			WeightsStore9[22] <= WeightsStore9[330];
			WeightsStore9[23] <= WeightsStore9[331];
			WeightsStore9[24] <= WeightsStore9[332];
			WeightsStore9[25] <= WeightsStore9[333];
			WeightsStore9[26] <= WeightsStore9[334];
			WeightsStore9[27] <= WeightsStore9[335];
		end else if(switchCounter == 32'd83)begin
			PixelsStore[0] <= PixelsStore[336];
			PixelsStore[1] <= PixelsStore[337];
			PixelsStore[2] <= PixelsStore[338];
			PixelsStore[3] <= PixelsStore[339];
			PixelsStore[4] <= PixelsStore[340];
			PixelsStore[5] <= PixelsStore[341];
			PixelsStore[6] <= PixelsStore[342];
			PixelsStore[7] <= PixelsStore[343];
			PixelsStore[8] <= PixelsStore[344];
			PixelsStore[9] <= PixelsStore[345];
			PixelsStore[10] <= PixelsStore[346];
			PixelsStore[11] <= PixelsStore[347];
			PixelsStore[12] <= PixelsStore[348];
			PixelsStore[13] <= PixelsStore[349];
			PixelsStore[14] <= PixelsStore[350];
			PixelsStore[15] <= PixelsStore[351];
			PixelsStore[16] <= PixelsStore[352];
			PixelsStore[17] <= PixelsStore[353];
			PixelsStore[18] <= PixelsStore[354];
			PixelsStore[19] <= PixelsStore[355];
			PixelsStore[20] <= PixelsStore[356];
			PixelsStore[21] <= PixelsStore[357];
			PixelsStore[22] <= PixelsStore[358];
			PixelsStore[23] <= PixelsStore[359];
			PixelsStore[24] <= PixelsStore[360];
			PixelsStore[25] <= PixelsStore[361];
			PixelsStore[26] <= PixelsStore[362];
			PixelsStore[27] <= PixelsStore[363];
			WeightsStore0[0] <= WeightsStore0[336];
			WeightsStore0[1] <= WeightsStore0[337];
			WeightsStore0[2] <= WeightsStore0[338];
			WeightsStore0[3] <= WeightsStore0[339];
			WeightsStore0[4] <= WeightsStore0[340];
			WeightsStore0[5] <= WeightsStore0[341];
			WeightsStore0[6] <= WeightsStore0[342];
			WeightsStore0[7] <= WeightsStore0[343];
			WeightsStore0[8] <= WeightsStore0[344];
			WeightsStore0[9] <= WeightsStore0[345];
			WeightsStore0[10] <= WeightsStore0[346];
			WeightsStore0[11] <= WeightsStore0[347];
			WeightsStore0[12] <= WeightsStore0[348];
			WeightsStore0[13] <= WeightsStore0[349];
			WeightsStore0[14] <= WeightsStore0[350];
			WeightsStore0[15] <= WeightsStore0[351];
			WeightsStore0[16] <= WeightsStore0[352];
			WeightsStore0[17] <= WeightsStore0[353];
			WeightsStore0[18] <= WeightsStore0[354];
			WeightsStore0[19] <= WeightsStore0[355];
			WeightsStore0[20] <= WeightsStore0[356];
			WeightsStore0[21] <= WeightsStore0[357];
			WeightsStore0[22] <= WeightsStore0[358];
			WeightsStore0[23] <= WeightsStore0[359];
			WeightsStore0[24] <= WeightsStore0[360];
			WeightsStore0[25] <= WeightsStore0[361];
			WeightsStore0[26] <= WeightsStore0[362];
			WeightsStore0[27] <= WeightsStore0[363];
			WeightsStore1[0] <= WeightsStore1[336];
			WeightsStore1[1] <= WeightsStore1[337];
			WeightsStore1[2] <= WeightsStore1[338];
			WeightsStore1[3] <= WeightsStore1[339];
			WeightsStore1[4] <= WeightsStore1[340];
			WeightsStore1[5] <= WeightsStore1[341];
			WeightsStore1[6] <= WeightsStore1[342];
			WeightsStore1[7] <= WeightsStore1[343];
			WeightsStore1[8] <= WeightsStore1[344];
			WeightsStore1[9] <= WeightsStore1[345];
			WeightsStore1[10] <= WeightsStore1[346];
			WeightsStore1[11] <= WeightsStore1[347];
			WeightsStore1[12] <= WeightsStore1[348];
			WeightsStore1[13] <= WeightsStore1[349];
			WeightsStore1[14] <= WeightsStore1[350];
			WeightsStore1[15] <= WeightsStore1[351];
			WeightsStore1[16] <= WeightsStore1[352];
			WeightsStore1[17] <= WeightsStore1[353];
			WeightsStore1[18] <= WeightsStore1[354];
			WeightsStore1[19] <= WeightsStore1[355];
			WeightsStore1[20] <= WeightsStore1[356];
			WeightsStore1[21] <= WeightsStore1[357];
			WeightsStore1[22] <= WeightsStore1[358];
			WeightsStore1[23] <= WeightsStore1[359];
			WeightsStore1[24] <= WeightsStore1[360];
			WeightsStore1[25] <= WeightsStore1[361];
			WeightsStore1[26] <= WeightsStore1[362];
			WeightsStore1[27] <= WeightsStore1[363];
			WeightsStore2[0] <= WeightsStore2[336];
			WeightsStore2[1] <= WeightsStore2[337];
			WeightsStore2[2] <= WeightsStore2[338];
			WeightsStore2[3] <= WeightsStore2[339];
			WeightsStore2[4] <= WeightsStore2[340];
			WeightsStore2[5] <= WeightsStore2[341];
			WeightsStore2[6] <= WeightsStore2[342];
			WeightsStore2[7] <= WeightsStore2[343];
			WeightsStore2[8] <= WeightsStore2[344];
			WeightsStore2[9] <= WeightsStore2[345];
			WeightsStore2[10] <= WeightsStore2[346];
			WeightsStore2[11] <= WeightsStore2[347];
			WeightsStore2[12] <= WeightsStore2[348];
			WeightsStore2[13] <= WeightsStore2[349];
			WeightsStore2[14] <= WeightsStore2[350];
			WeightsStore2[15] <= WeightsStore2[351];
			WeightsStore2[16] <= WeightsStore2[352];
			WeightsStore2[17] <= WeightsStore2[353];
			WeightsStore2[18] <= WeightsStore2[354];
			WeightsStore2[19] <= WeightsStore2[355];
			WeightsStore2[20] <= WeightsStore2[356];
			WeightsStore2[21] <= WeightsStore2[357];
			WeightsStore2[22] <= WeightsStore2[358];
			WeightsStore2[23] <= WeightsStore2[359];
			WeightsStore2[24] <= WeightsStore2[360];
			WeightsStore2[25] <= WeightsStore2[361];
			WeightsStore2[26] <= WeightsStore2[362];
			WeightsStore2[27] <= WeightsStore2[363];
			WeightsStore3[0] <= WeightsStore3[336];
			WeightsStore3[1] <= WeightsStore3[337];
			WeightsStore3[2] <= WeightsStore3[338];
			WeightsStore3[3] <= WeightsStore3[339];
			WeightsStore3[4] <= WeightsStore3[340];
			WeightsStore3[5] <= WeightsStore3[341];
			WeightsStore3[6] <= WeightsStore3[342];
			WeightsStore3[7] <= WeightsStore3[343];
			WeightsStore3[8] <= WeightsStore3[344];
			WeightsStore3[9] <= WeightsStore3[345];
			WeightsStore3[10] <= WeightsStore3[346];
			WeightsStore3[11] <= WeightsStore3[347];
			WeightsStore3[12] <= WeightsStore3[348];
			WeightsStore3[13] <= WeightsStore3[349];
			WeightsStore3[14] <= WeightsStore3[350];
			WeightsStore3[15] <= WeightsStore3[351];
			WeightsStore3[16] <= WeightsStore3[352];
			WeightsStore3[17] <= WeightsStore3[353];
			WeightsStore3[18] <= WeightsStore3[354];
			WeightsStore3[19] <= WeightsStore3[355];
			WeightsStore3[20] <= WeightsStore3[356];
			WeightsStore3[21] <= WeightsStore3[357];
			WeightsStore3[22] <= WeightsStore3[358];
			WeightsStore3[23] <= WeightsStore3[359];
			WeightsStore3[24] <= WeightsStore3[360];
			WeightsStore3[25] <= WeightsStore3[361];
			WeightsStore3[26] <= WeightsStore3[362];
			WeightsStore3[27] <= WeightsStore3[363];
			WeightsStore4[0] <= WeightsStore4[336];
			WeightsStore4[1] <= WeightsStore4[337];
			WeightsStore4[2] <= WeightsStore4[338];
			WeightsStore4[3] <= WeightsStore4[339];
			WeightsStore4[4] <= WeightsStore4[340];
			WeightsStore4[5] <= WeightsStore4[341];
			WeightsStore4[6] <= WeightsStore4[342];
			WeightsStore4[7] <= WeightsStore4[343];
			WeightsStore4[8] <= WeightsStore4[344];
			WeightsStore4[9] <= WeightsStore4[345];
			WeightsStore4[10] <= WeightsStore4[346];
			WeightsStore4[11] <= WeightsStore4[347];
			WeightsStore4[12] <= WeightsStore4[348];
			WeightsStore4[13] <= WeightsStore4[349];
			WeightsStore4[14] <= WeightsStore4[350];
			WeightsStore4[15] <= WeightsStore4[351];
			WeightsStore4[16] <= WeightsStore4[352];
			WeightsStore4[17] <= WeightsStore4[353];
			WeightsStore4[18] <= WeightsStore4[354];
			WeightsStore4[19] <= WeightsStore4[355];
			WeightsStore4[20] <= WeightsStore4[356];
			WeightsStore4[21] <= WeightsStore4[357];
			WeightsStore4[22] <= WeightsStore4[358];
			WeightsStore4[23] <= WeightsStore4[359];
			WeightsStore4[24] <= WeightsStore4[360];
			WeightsStore4[25] <= WeightsStore4[361];
			WeightsStore4[26] <= WeightsStore4[362];
			WeightsStore4[27] <= WeightsStore4[363];
			WeightsStore5[0] <= WeightsStore5[336];
			WeightsStore5[1] <= WeightsStore5[337];
			WeightsStore5[2] <= WeightsStore5[338];
			WeightsStore5[3] <= WeightsStore5[339];
			WeightsStore5[4] <= WeightsStore5[340];
			WeightsStore5[5] <= WeightsStore5[341];
			WeightsStore5[6] <= WeightsStore5[342];
			WeightsStore5[7] <= WeightsStore5[343];
			WeightsStore5[8] <= WeightsStore5[344];
			WeightsStore5[9] <= WeightsStore5[345];
			WeightsStore5[10] <= WeightsStore5[346];
			WeightsStore5[11] <= WeightsStore5[347];
			WeightsStore5[12] <= WeightsStore5[348];
			WeightsStore5[13] <= WeightsStore5[349];
			WeightsStore5[14] <= WeightsStore5[350];
			WeightsStore5[15] <= WeightsStore5[351];
			WeightsStore5[16] <= WeightsStore5[352];
			WeightsStore5[17] <= WeightsStore5[353];
			WeightsStore5[18] <= WeightsStore5[354];
			WeightsStore5[19] <= WeightsStore5[355];
			WeightsStore5[20] <= WeightsStore5[356];
			WeightsStore5[21] <= WeightsStore5[357];
			WeightsStore5[22] <= WeightsStore5[358];
			WeightsStore5[23] <= WeightsStore5[359];
			WeightsStore5[24] <= WeightsStore5[360];
			WeightsStore5[25] <= WeightsStore5[361];
			WeightsStore5[26] <= WeightsStore5[362];
			WeightsStore5[27] <= WeightsStore5[363];
			WeightsStore6[0] <= WeightsStore6[336];
			WeightsStore6[1] <= WeightsStore6[337];
			WeightsStore6[2] <= WeightsStore6[338];
			WeightsStore6[3] <= WeightsStore6[339];
			WeightsStore6[4] <= WeightsStore6[340];
			WeightsStore6[5] <= WeightsStore6[341];
			WeightsStore6[6] <= WeightsStore6[342];
			WeightsStore6[7] <= WeightsStore6[343];
			WeightsStore6[8] <= WeightsStore6[344];
			WeightsStore6[9] <= WeightsStore6[345];
			WeightsStore6[10] <= WeightsStore6[346];
			WeightsStore6[11] <= WeightsStore6[347];
			WeightsStore6[12] <= WeightsStore6[348];
			WeightsStore6[13] <= WeightsStore6[349];
			WeightsStore6[14] <= WeightsStore6[350];
			WeightsStore6[15] <= WeightsStore6[351];
			WeightsStore6[16] <= WeightsStore6[352];
			WeightsStore6[17] <= WeightsStore6[353];
			WeightsStore6[18] <= WeightsStore6[354];
			WeightsStore6[19] <= WeightsStore6[355];
			WeightsStore6[20] <= WeightsStore6[356];
			WeightsStore6[21] <= WeightsStore6[357];
			WeightsStore6[22] <= WeightsStore6[358];
			WeightsStore6[23] <= WeightsStore6[359];
			WeightsStore6[24] <= WeightsStore6[360];
			WeightsStore6[25] <= WeightsStore6[361];
			WeightsStore6[26] <= WeightsStore6[362];
			WeightsStore6[27] <= WeightsStore6[363];
			WeightsStore7[0] <= WeightsStore7[336];
			WeightsStore7[1] <= WeightsStore7[337];
			WeightsStore7[2] <= WeightsStore7[338];
			WeightsStore7[3] <= WeightsStore7[339];
			WeightsStore7[4] <= WeightsStore7[340];
			WeightsStore7[5] <= WeightsStore7[341];
			WeightsStore7[6] <= WeightsStore7[342];
			WeightsStore7[7] <= WeightsStore7[343];
			WeightsStore7[8] <= WeightsStore7[344];
			WeightsStore7[9] <= WeightsStore7[345];
			WeightsStore7[10] <= WeightsStore7[346];
			WeightsStore7[11] <= WeightsStore7[347];
			WeightsStore7[12] <= WeightsStore7[348];
			WeightsStore7[13] <= WeightsStore7[349];
			WeightsStore7[14] <= WeightsStore7[350];
			WeightsStore7[15] <= WeightsStore7[351];
			WeightsStore7[16] <= WeightsStore7[352];
			WeightsStore7[17] <= WeightsStore7[353];
			WeightsStore7[18] <= WeightsStore7[354];
			WeightsStore7[19] <= WeightsStore7[355];
			WeightsStore7[20] <= WeightsStore7[356];
			WeightsStore7[21] <= WeightsStore7[357];
			WeightsStore7[22] <= WeightsStore7[358];
			WeightsStore7[23] <= WeightsStore7[359];
			WeightsStore7[24] <= WeightsStore7[360];
			WeightsStore7[25] <= WeightsStore7[361];
			WeightsStore7[26] <= WeightsStore7[362];
			WeightsStore7[27] <= WeightsStore7[363];
			WeightsStore8[0] <= WeightsStore8[336];
			WeightsStore8[1] <= WeightsStore8[337];
			WeightsStore8[2] <= WeightsStore8[338];
			WeightsStore8[3] <= WeightsStore8[339];
			WeightsStore8[4] <= WeightsStore8[340];
			WeightsStore8[5] <= WeightsStore8[341];
			WeightsStore8[6] <= WeightsStore8[342];
			WeightsStore8[7] <= WeightsStore8[343];
			WeightsStore8[8] <= WeightsStore8[344];
			WeightsStore8[9] <= WeightsStore8[345];
			WeightsStore8[10] <= WeightsStore8[346];
			WeightsStore8[11] <= WeightsStore8[347];
			WeightsStore8[12] <= WeightsStore8[348];
			WeightsStore8[13] <= WeightsStore8[349];
			WeightsStore8[14] <= WeightsStore8[350];
			WeightsStore8[15] <= WeightsStore8[351];
			WeightsStore8[16] <= WeightsStore8[352];
			WeightsStore8[17] <= WeightsStore8[353];
			WeightsStore8[18] <= WeightsStore8[354];
			WeightsStore8[19] <= WeightsStore8[355];
			WeightsStore8[20] <= WeightsStore8[356];
			WeightsStore8[21] <= WeightsStore8[357];
			WeightsStore8[22] <= WeightsStore8[358];
			WeightsStore8[23] <= WeightsStore8[359];
			WeightsStore8[24] <= WeightsStore8[360];
			WeightsStore8[25] <= WeightsStore8[361];
			WeightsStore8[26] <= WeightsStore8[362];
			WeightsStore8[27] <= WeightsStore8[363];
			WeightsStore9[0] <= WeightsStore9[336];
			WeightsStore9[1] <= WeightsStore9[337];
			WeightsStore9[2] <= WeightsStore9[338];
			WeightsStore9[3] <= WeightsStore9[339];
			WeightsStore9[4] <= WeightsStore9[340];
			WeightsStore9[5] <= WeightsStore9[341];
			WeightsStore9[6] <= WeightsStore9[342];
			WeightsStore9[7] <= WeightsStore9[343];
			WeightsStore9[8] <= WeightsStore9[344];
			WeightsStore9[9] <= WeightsStore9[345];
			WeightsStore9[10] <= WeightsStore9[346];
			WeightsStore9[11] <= WeightsStore9[347];
			WeightsStore9[12] <= WeightsStore9[348];
			WeightsStore9[13] <= WeightsStore9[349];
			WeightsStore9[14] <= WeightsStore9[350];
			WeightsStore9[15] <= WeightsStore9[351];
			WeightsStore9[16] <= WeightsStore9[352];
			WeightsStore9[17] <= WeightsStore9[353];
			WeightsStore9[18] <= WeightsStore9[354];
			WeightsStore9[19] <= WeightsStore9[355];
			WeightsStore9[20] <= WeightsStore9[356];
			WeightsStore9[21] <= WeightsStore9[357];
			WeightsStore9[22] <= WeightsStore9[358];
			WeightsStore9[23] <= WeightsStore9[359];
			WeightsStore9[24] <= WeightsStore9[360];
			WeightsStore9[25] <= WeightsStore9[361];
			WeightsStore9[26] <= WeightsStore9[362];
			WeightsStore9[27] <= WeightsStore9[363];
		end else if(switchCounter == 32'd90)begin
			PixelsStore[0] <= PixelsStore[364];
			PixelsStore[1] <= PixelsStore[365];
			PixelsStore[2] <= PixelsStore[366];
			PixelsStore[3] <= PixelsStore[367];
			PixelsStore[4] <= PixelsStore[368];
			PixelsStore[5] <= PixelsStore[369];
			PixelsStore[6] <= PixelsStore[370];
			PixelsStore[7] <= PixelsStore[371];
			PixelsStore[8] <= PixelsStore[372];
			PixelsStore[9] <= PixelsStore[373];
			PixelsStore[10] <= PixelsStore[374];
			PixelsStore[11] <= PixelsStore[375];
			PixelsStore[12] <= PixelsStore[376];
			PixelsStore[13] <= PixelsStore[377];
			PixelsStore[14] <= PixelsStore[378];
			PixelsStore[15] <= PixelsStore[379];
			PixelsStore[16] <= PixelsStore[380];
			PixelsStore[17] <= PixelsStore[381];
			PixelsStore[18] <= PixelsStore[382];
			PixelsStore[19] <= PixelsStore[383];
			PixelsStore[20] <= PixelsStore[384];
			PixelsStore[21] <= PixelsStore[385];
			PixelsStore[22] <= PixelsStore[386];
			PixelsStore[23] <= PixelsStore[387];
			PixelsStore[24] <= PixelsStore[388];
			PixelsStore[25] <= PixelsStore[389];
			PixelsStore[26] <= PixelsStore[390];
			PixelsStore[27] <= PixelsStore[391];
			WeightsStore0[0] <= WeightsStore0[364];
			WeightsStore0[1] <= WeightsStore0[365];
			WeightsStore0[2] <= WeightsStore0[366];
			WeightsStore0[3] <= WeightsStore0[367];
			WeightsStore0[4] <= WeightsStore0[368];
			WeightsStore0[5] <= WeightsStore0[369];
			WeightsStore0[6] <= WeightsStore0[370];
			WeightsStore0[7] <= WeightsStore0[371];
			WeightsStore0[8] <= WeightsStore0[372];
			WeightsStore0[9] <= WeightsStore0[373];
			WeightsStore0[10] <= WeightsStore0[374];
			WeightsStore0[11] <= WeightsStore0[375];
			WeightsStore0[12] <= WeightsStore0[376];
			WeightsStore0[13] <= WeightsStore0[377];
			WeightsStore0[14] <= WeightsStore0[378];
			WeightsStore0[15] <= WeightsStore0[379];
			WeightsStore0[16] <= WeightsStore0[380];
			WeightsStore0[17] <= WeightsStore0[381];
			WeightsStore0[18] <= WeightsStore0[382];
			WeightsStore0[19] <= WeightsStore0[383];
			WeightsStore0[20] <= WeightsStore0[384];
			WeightsStore0[21] <= WeightsStore0[385];
			WeightsStore0[22] <= WeightsStore0[386];
			WeightsStore0[23] <= WeightsStore0[387];
			WeightsStore0[24] <= WeightsStore0[388];
			WeightsStore0[25] <= WeightsStore0[389];
			WeightsStore0[26] <= WeightsStore0[390];
			WeightsStore0[27] <= WeightsStore0[391];
			WeightsStore1[0] <= WeightsStore1[364];
			WeightsStore1[1] <= WeightsStore1[365];
			WeightsStore1[2] <= WeightsStore1[366];
			WeightsStore1[3] <= WeightsStore1[367];
			WeightsStore1[4] <= WeightsStore1[368];
			WeightsStore1[5] <= WeightsStore1[369];
			WeightsStore1[6] <= WeightsStore1[370];
			WeightsStore1[7] <= WeightsStore1[371];
			WeightsStore1[8] <= WeightsStore1[372];
			WeightsStore1[9] <= WeightsStore1[373];
			WeightsStore1[10] <= WeightsStore1[374];
			WeightsStore1[11] <= WeightsStore1[375];
			WeightsStore1[12] <= WeightsStore1[376];
			WeightsStore1[13] <= WeightsStore1[377];
			WeightsStore1[14] <= WeightsStore1[378];
			WeightsStore1[15] <= WeightsStore1[379];
			WeightsStore1[16] <= WeightsStore1[380];
			WeightsStore1[17] <= WeightsStore1[381];
			WeightsStore1[18] <= WeightsStore1[382];
			WeightsStore1[19] <= WeightsStore1[383];
			WeightsStore1[20] <= WeightsStore1[384];
			WeightsStore1[21] <= WeightsStore1[385];
			WeightsStore1[22] <= WeightsStore1[386];
			WeightsStore1[23] <= WeightsStore1[387];
			WeightsStore1[24] <= WeightsStore1[388];
			WeightsStore1[25] <= WeightsStore1[389];
			WeightsStore1[26] <= WeightsStore1[390];
			WeightsStore1[27] <= WeightsStore1[391];
			WeightsStore2[0] <= WeightsStore2[364];
			WeightsStore2[1] <= WeightsStore2[365];
			WeightsStore2[2] <= WeightsStore2[366];
			WeightsStore2[3] <= WeightsStore2[367];
			WeightsStore2[4] <= WeightsStore2[368];
			WeightsStore2[5] <= WeightsStore2[369];
			WeightsStore2[6] <= WeightsStore2[370];
			WeightsStore2[7] <= WeightsStore2[371];
			WeightsStore2[8] <= WeightsStore2[372];
			WeightsStore2[9] <= WeightsStore2[373];
			WeightsStore2[10] <= WeightsStore2[374];
			WeightsStore2[11] <= WeightsStore2[375];
			WeightsStore2[12] <= WeightsStore2[376];
			WeightsStore2[13] <= WeightsStore2[377];
			WeightsStore2[14] <= WeightsStore2[378];
			WeightsStore2[15] <= WeightsStore2[379];
			WeightsStore2[16] <= WeightsStore2[380];
			WeightsStore2[17] <= WeightsStore2[381];
			WeightsStore2[18] <= WeightsStore2[382];
			WeightsStore2[19] <= WeightsStore2[383];
			WeightsStore2[20] <= WeightsStore2[384];
			WeightsStore2[21] <= WeightsStore2[385];
			WeightsStore2[22] <= WeightsStore2[386];
			WeightsStore2[23] <= WeightsStore2[387];
			WeightsStore2[24] <= WeightsStore2[388];
			WeightsStore2[25] <= WeightsStore2[389];
			WeightsStore2[26] <= WeightsStore2[390];
			WeightsStore2[27] <= WeightsStore2[391];
			WeightsStore3[0] <= WeightsStore3[364];
			WeightsStore3[1] <= WeightsStore3[365];
			WeightsStore3[2] <= WeightsStore3[366];
			WeightsStore3[3] <= WeightsStore3[367];
			WeightsStore3[4] <= WeightsStore3[368];
			WeightsStore3[5] <= WeightsStore3[369];
			WeightsStore3[6] <= WeightsStore3[370];
			WeightsStore3[7] <= WeightsStore3[371];
			WeightsStore3[8] <= WeightsStore3[372];
			WeightsStore3[9] <= WeightsStore3[373];
			WeightsStore3[10] <= WeightsStore3[374];
			WeightsStore3[11] <= WeightsStore3[375];
			WeightsStore3[12] <= WeightsStore3[376];
			WeightsStore3[13] <= WeightsStore3[377];
			WeightsStore3[14] <= WeightsStore3[378];
			WeightsStore3[15] <= WeightsStore3[379];
			WeightsStore3[16] <= WeightsStore3[380];
			WeightsStore3[17] <= WeightsStore3[381];
			WeightsStore3[18] <= WeightsStore3[382];
			WeightsStore3[19] <= WeightsStore3[383];
			WeightsStore3[20] <= WeightsStore3[384];
			WeightsStore3[21] <= WeightsStore3[385];
			WeightsStore3[22] <= WeightsStore3[386];
			WeightsStore3[23] <= WeightsStore3[387];
			WeightsStore3[24] <= WeightsStore3[388];
			WeightsStore3[25] <= WeightsStore3[389];
			WeightsStore3[26] <= WeightsStore3[390];
			WeightsStore3[27] <= WeightsStore3[391];
			WeightsStore4[0] <= WeightsStore4[364];
			WeightsStore4[1] <= WeightsStore4[365];
			WeightsStore4[2] <= WeightsStore4[366];
			WeightsStore4[3] <= WeightsStore4[367];
			WeightsStore4[4] <= WeightsStore4[368];
			WeightsStore4[5] <= WeightsStore4[369];
			WeightsStore4[6] <= WeightsStore4[370];
			WeightsStore4[7] <= WeightsStore4[371];
			WeightsStore4[8] <= WeightsStore4[372];
			WeightsStore4[9] <= WeightsStore4[373];
			WeightsStore4[10] <= WeightsStore4[374];
			WeightsStore4[11] <= WeightsStore4[375];
			WeightsStore4[12] <= WeightsStore4[376];
			WeightsStore4[13] <= WeightsStore4[377];
			WeightsStore4[14] <= WeightsStore4[378];
			WeightsStore4[15] <= WeightsStore4[379];
			WeightsStore4[16] <= WeightsStore4[380];
			WeightsStore4[17] <= WeightsStore4[381];
			WeightsStore4[18] <= WeightsStore4[382];
			WeightsStore4[19] <= WeightsStore4[383];
			WeightsStore4[20] <= WeightsStore4[384];
			WeightsStore4[21] <= WeightsStore4[385];
			WeightsStore4[22] <= WeightsStore4[386];
			WeightsStore4[23] <= WeightsStore4[387];
			WeightsStore4[24] <= WeightsStore4[388];
			WeightsStore4[25] <= WeightsStore4[389];
			WeightsStore4[26] <= WeightsStore4[390];
			WeightsStore4[27] <= WeightsStore4[391];
			WeightsStore5[0] <= WeightsStore5[364];
			WeightsStore5[1] <= WeightsStore5[365];
			WeightsStore5[2] <= WeightsStore5[366];
			WeightsStore5[3] <= WeightsStore5[367];
			WeightsStore5[4] <= WeightsStore5[368];
			WeightsStore5[5] <= WeightsStore5[369];
			WeightsStore5[6] <= WeightsStore5[370];
			WeightsStore5[7] <= WeightsStore5[371];
			WeightsStore5[8] <= WeightsStore5[372];
			WeightsStore5[9] <= WeightsStore5[373];
			WeightsStore5[10] <= WeightsStore5[374];
			WeightsStore5[11] <= WeightsStore5[375];
			WeightsStore5[12] <= WeightsStore5[376];
			WeightsStore5[13] <= WeightsStore5[377];
			WeightsStore5[14] <= WeightsStore5[378];
			WeightsStore5[15] <= WeightsStore5[379];
			WeightsStore5[16] <= WeightsStore5[380];
			WeightsStore5[17] <= WeightsStore5[381];
			WeightsStore5[18] <= WeightsStore5[382];
			WeightsStore5[19] <= WeightsStore5[383];
			WeightsStore5[20] <= WeightsStore5[384];
			WeightsStore5[21] <= WeightsStore5[385];
			WeightsStore5[22] <= WeightsStore5[386];
			WeightsStore5[23] <= WeightsStore5[387];
			WeightsStore5[24] <= WeightsStore5[388];
			WeightsStore5[25] <= WeightsStore5[389];
			WeightsStore5[26] <= WeightsStore5[390];
			WeightsStore5[27] <= WeightsStore5[391];
			WeightsStore6[0] <= WeightsStore6[364];
			WeightsStore6[1] <= WeightsStore6[365];
			WeightsStore6[2] <= WeightsStore6[366];
			WeightsStore6[3] <= WeightsStore6[367];
			WeightsStore6[4] <= WeightsStore6[368];
			WeightsStore6[5] <= WeightsStore6[369];
			WeightsStore6[6] <= WeightsStore6[370];
			WeightsStore6[7] <= WeightsStore6[371];
			WeightsStore6[8] <= WeightsStore6[372];
			WeightsStore6[9] <= WeightsStore6[373];
			WeightsStore6[10] <= WeightsStore6[374];
			WeightsStore6[11] <= WeightsStore6[375];
			WeightsStore6[12] <= WeightsStore6[376];
			WeightsStore6[13] <= WeightsStore6[377];
			WeightsStore6[14] <= WeightsStore6[378];
			WeightsStore6[15] <= WeightsStore6[379];
			WeightsStore6[16] <= WeightsStore6[380];
			WeightsStore6[17] <= WeightsStore6[381];
			WeightsStore6[18] <= WeightsStore6[382];
			WeightsStore6[19] <= WeightsStore6[383];
			WeightsStore6[20] <= WeightsStore6[384];
			WeightsStore6[21] <= WeightsStore6[385];
			WeightsStore6[22] <= WeightsStore6[386];
			WeightsStore6[23] <= WeightsStore6[387];
			WeightsStore6[24] <= WeightsStore6[388];
			WeightsStore6[25] <= WeightsStore6[389];
			WeightsStore6[26] <= WeightsStore6[390];
			WeightsStore6[27] <= WeightsStore6[391];
			WeightsStore7[0] <= WeightsStore7[364];
			WeightsStore7[1] <= WeightsStore7[365];
			WeightsStore7[2] <= WeightsStore7[366];
			WeightsStore7[3] <= WeightsStore7[367];
			WeightsStore7[4] <= WeightsStore7[368];
			WeightsStore7[5] <= WeightsStore7[369];
			WeightsStore7[6] <= WeightsStore7[370];
			WeightsStore7[7] <= WeightsStore7[371];
			WeightsStore7[8] <= WeightsStore7[372];
			WeightsStore7[9] <= WeightsStore7[373];
			WeightsStore7[10] <= WeightsStore7[374];
			WeightsStore7[11] <= WeightsStore7[375];
			WeightsStore7[12] <= WeightsStore7[376];
			WeightsStore7[13] <= WeightsStore7[377];
			WeightsStore7[14] <= WeightsStore7[378];
			WeightsStore7[15] <= WeightsStore7[379];
			WeightsStore7[16] <= WeightsStore7[380];
			WeightsStore7[17] <= WeightsStore7[381];
			WeightsStore7[18] <= WeightsStore7[382];
			WeightsStore7[19] <= WeightsStore7[383];
			WeightsStore7[20] <= WeightsStore7[384];
			WeightsStore7[21] <= WeightsStore7[385];
			WeightsStore7[22] <= WeightsStore7[386];
			WeightsStore7[23] <= WeightsStore7[387];
			WeightsStore7[24] <= WeightsStore7[388];
			WeightsStore7[25] <= WeightsStore7[389];
			WeightsStore7[26] <= WeightsStore7[390];
			WeightsStore7[27] <= WeightsStore7[391];
			WeightsStore8[0] <= WeightsStore8[364];
			WeightsStore8[1] <= WeightsStore8[365];
			WeightsStore8[2] <= WeightsStore8[366];
			WeightsStore8[3] <= WeightsStore8[367];
			WeightsStore8[4] <= WeightsStore8[368];
			WeightsStore8[5] <= WeightsStore8[369];
			WeightsStore8[6] <= WeightsStore8[370];
			WeightsStore8[7] <= WeightsStore8[371];
			WeightsStore8[8] <= WeightsStore8[372];
			WeightsStore8[9] <= WeightsStore8[373];
			WeightsStore8[10] <= WeightsStore8[374];
			WeightsStore8[11] <= WeightsStore8[375];
			WeightsStore8[12] <= WeightsStore8[376];
			WeightsStore8[13] <= WeightsStore8[377];
			WeightsStore8[14] <= WeightsStore8[378];
			WeightsStore8[15] <= WeightsStore8[379];
			WeightsStore8[16] <= WeightsStore8[380];
			WeightsStore8[17] <= WeightsStore8[381];
			WeightsStore8[18] <= WeightsStore8[382];
			WeightsStore8[19] <= WeightsStore8[383];
			WeightsStore8[20] <= WeightsStore8[384];
			WeightsStore8[21] <= WeightsStore8[385];
			WeightsStore8[22] <= WeightsStore8[386];
			WeightsStore8[23] <= WeightsStore8[387];
			WeightsStore8[24] <= WeightsStore8[388];
			WeightsStore8[25] <= WeightsStore8[389];
			WeightsStore8[26] <= WeightsStore8[390];
			WeightsStore8[27] <= WeightsStore8[391];
			WeightsStore9[0] <= WeightsStore9[364];
			WeightsStore9[1] <= WeightsStore9[365];
			WeightsStore9[2] <= WeightsStore9[366];
			WeightsStore9[3] <= WeightsStore9[367];
			WeightsStore9[4] <= WeightsStore9[368];
			WeightsStore9[5] <= WeightsStore9[369];
			WeightsStore9[6] <= WeightsStore9[370];
			WeightsStore9[7] <= WeightsStore9[371];
			WeightsStore9[8] <= WeightsStore9[372];
			WeightsStore9[9] <= WeightsStore9[373];
			WeightsStore9[10] <= WeightsStore9[374];
			WeightsStore9[11] <= WeightsStore9[375];
			WeightsStore9[12] <= WeightsStore9[376];
			WeightsStore9[13] <= WeightsStore9[377];
			WeightsStore9[14] <= WeightsStore9[378];
			WeightsStore9[15] <= WeightsStore9[379];
			WeightsStore9[16] <= WeightsStore9[380];
			WeightsStore9[17] <= WeightsStore9[381];
			WeightsStore9[18] <= WeightsStore9[382];
			WeightsStore9[19] <= WeightsStore9[383];
			WeightsStore9[20] <= WeightsStore9[384];
			WeightsStore9[21] <= WeightsStore9[385];
			WeightsStore9[22] <= WeightsStore9[386];
			WeightsStore9[23] <= WeightsStore9[387];
			WeightsStore9[24] <= WeightsStore9[388];
			WeightsStore9[25] <= WeightsStore9[389];
			WeightsStore9[26] <= WeightsStore9[390];
			WeightsStore9[27] <= WeightsStore9[391];
		end else if(switchCounter == 32'd97)begin
			PixelsStore[0] <= PixelsStore[392];
			PixelsStore[1] <= PixelsStore[393];
			PixelsStore[2] <= PixelsStore[394];
			PixelsStore[3] <= PixelsStore[395];
			PixelsStore[4] <= PixelsStore[396];
			PixelsStore[5] <= PixelsStore[397];
			PixelsStore[6] <= PixelsStore[398];
			PixelsStore[7] <= PixelsStore[399];
			PixelsStore[8] <= PixelsStore[400];
			PixelsStore[9] <= PixelsStore[401];
			PixelsStore[10] <= PixelsStore[402];
			PixelsStore[11] <= PixelsStore[403];
			PixelsStore[12] <= PixelsStore[404];
			PixelsStore[13] <= PixelsStore[405];
			PixelsStore[14] <= PixelsStore[406];
			PixelsStore[15] <= PixelsStore[407];
			PixelsStore[16] <= PixelsStore[408];
			PixelsStore[17] <= PixelsStore[409];
			PixelsStore[18] <= PixelsStore[410];
			PixelsStore[19] <= PixelsStore[411];
			PixelsStore[20] <= PixelsStore[412];
			PixelsStore[21] <= PixelsStore[413];
			PixelsStore[22] <= PixelsStore[414];
			PixelsStore[23] <= PixelsStore[415];
			PixelsStore[24] <= PixelsStore[416];
			PixelsStore[25] <= PixelsStore[417];
			PixelsStore[26] <= PixelsStore[418];
			PixelsStore[27] <= PixelsStore[419];
			WeightsStore0[0] <= WeightsStore0[392];
			WeightsStore0[1] <= WeightsStore0[393];
			WeightsStore0[2] <= WeightsStore0[394];
			WeightsStore0[3] <= WeightsStore0[395];
			WeightsStore0[4] <= WeightsStore0[396];
			WeightsStore0[5] <= WeightsStore0[397];
			WeightsStore0[6] <= WeightsStore0[398];
			WeightsStore0[7] <= WeightsStore0[399];
			WeightsStore0[8] <= WeightsStore0[400];
			WeightsStore0[9] <= WeightsStore0[401];
			WeightsStore0[10] <= WeightsStore0[402];
			WeightsStore0[11] <= WeightsStore0[403];
			WeightsStore0[12] <= WeightsStore0[404];
			WeightsStore0[13] <= WeightsStore0[405];
			WeightsStore0[14] <= WeightsStore0[406];
			WeightsStore0[15] <= WeightsStore0[407];
			WeightsStore0[16] <= WeightsStore0[408];
			WeightsStore0[17] <= WeightsStore0[409];
			WeightsStore0[18] <= WeightsStore0[410];
			WeightsStore0[19] <= WeightsStore0[411];
			WeightsStore0[20] <= WeightsStore0[412];
			WeightsStore0[21] <= WeightsStore0[413];
			WeightsStore0[22] <= WeightsStore0[414];
			WeightsStore0[23] <= WeightsStore0[415];
			WeightsStore0[24] <= WeightsStore0[416];
			WeightsStore0[25] <= WeightsStore0[417];
			WeightsStore0[26] <= WeightsStore0[418];
			WeightsStore0[27] <= WeightsStore0[419];
			WeightsStore1[0] <= WeightsStore1[392];
			WeightsStore1[1] <= WeightsStore1[393];
			WeightsStore1[2] <= WeightsStore1[394];
			WeightsStore1[3] <= WeightsStore1[395];
			WeightsStore1[4] <= WeightsStore1[396];
			WeightsStore1[5] <= WeightsStore1[397];
			WeightsStore1[6] <= WeightsStore1[398];
			WeightsStore1[7] <= WeightsStore1[399];
			WeightsStore1[8] <= WeightsStore1[400];
			WeightsStore1[9] <= WeightsStore1[401];
			WeightsStore1[10] <= WeightsStore1[402];
			WeightsStore1[11] <= WeightsStore1[403];
			WeightsStore1[12] <= WeightsStore1[404];
			WeightsStore1[13] <= WeightsStore1[405];
			WeightsStore1[14] <= WeightsStore1[406];
			WeightsStore1[15] <= WeightsStore1[407];
			WeightsStore1[16] <= WeightsStore1[408];
			WeightsStore1[17] <= WeightsStore1[409];
			WeightsStore1[18] <= WeightsStore1[410];
			WeightsStore1[19] <= WeightsStore1[411];
			WeightsStore1[20] <= WeightsStore1[412];
			WeightsStore1[21] <= WeightsStore1[413];
			WeightsStore1[22] <= WeightsStore1[414];
			WeightsStore1[23] <= WeightsStore1[415];
			WeightsStore1[24] <= WeightsStore1[416];
			WeightsStore1[25] <= WeightsStore1[417];
			WeightsStore1[26] <= WeightsStore1[418];
			WeightsStore1[27] <= WeightsStore1[419];
			WeightsStore2[0] <= WeightsStore2[392];
			WeightsStore2[1] <= WeightsStore2[393];
			WeightsStore2[2] <= WeightsStore2[394];
			WeightsStore2[3] <= WeightsStore2[395];
			WeightsStore2[4] <= WeightsStore2[396];
			WeightsStore2[5] <= WeightsStore2[397];
			WeightsStore2[6] <= WeightsStore2[398];
			WeightsStore2[7] <= WeightsStore2[399];
			WeightsStore2[8] <= WeightsStore2[400];
			WeightsStore2[9] <= WeightsStore2[401];
			WeightsStore2[10] <= WeightsStore2[402];
			WeightsStore2[11] <= WeightsStore2[403];
			WeightsStore2[12] <= WeightsStore2[404];
			WeightsStore2[13] <= WeightsStore2[405];
			WeightsStore2[14] <= WeightsStore2[406];
			WeightsStore2[15] <= WeightsStore2[407];
			WeightsStore2[16] <= WeightsStore2[408];
			WeightsStore2[17] <= WeightsStore2[409];
			WeightsStore2[18] <= WeightsStore2[410];
			WeightsStore2[19] <= WeightsStore2[411];
			WeightsStore2[20] <= WeightsStore2[412];
			WeightsStore2[21] <= WeightsStore2[413];
			WeightsStore2[22] <= WeightsStore2[414];
			WeightsStore2[23] <= WeightsStore2[415];
			WeightsStore2[24] <= WeightsStore2[416];
			WeightsStore2[25] <= WeightsStore2[417];
			WeightsStore2[26] <= WeightsStore2[418];
			WeightsStore2[27] <= WeightsStore2[419];
			WeightsStore3[0] <= WeightsStore3[392];
			WeightsStore3[1] <= WeightsStore3[393];
			WeightsStore3[2] <= WeightsStore3[394];
			WeightsStore3[3] <= WeightsStore3[395];
			WeightsStore3[4] <= WeightsStore3[396];
			WeightsStore3[5] <= WeightsStore3[397];
			WeightsStore3[6] <= WeightsStore3[398];
			WeightsStore3[7] <= WeightsStore3[399];
			WeightsStore3[8] <= WeightsStore3[400];
			WeightsStore3[9] <= WeightsStore3[401];
			WeightsStore3[10] <= WeightsStore3[402];
			WeightsStore3[11] <= WeightsStore3[403];
			WeightsStore3[12] <= WeightsStore3[404];
			WeightsStore3[13] <= WeightsStore3[405];
			WeightsStore3[14] <= WeightsStore3[406];
			WeightsStore3[15] <= WeightsStore3[407];
			WeightsStore3[16] <= WeightsStore3[408];
			WeightsStore3[17] <= WeightsStore3[409];
			WeightsStore3[18] <= WeightsStore3[410];
			WeightsStore3[19] <= WeightsStore3[411];
			WeightsStore3[20] <= WeightsStore3[412];
			WeightsStore3[21] <= WeightsStore3[413];
			WeightsStore3[22] <= WeightsStore3[414];
			WeightsStore3[23] <= WeightsStore3[415];
			WeightsStore3[24] <= WeightsStore3[416];
			WeightsStore3[25] <= WeightsStore3[417];
			WeightsStore3[26] <= WeightsStore3[418];
			WeightsStore3[27] <= WeightsStore3[419];
			WeightsStore4[0] <= WeightsStore4[392];
			WeightsStore4[1] <= WeightsStore4[393];
			WeightsStore4[2] <= WeightsStore4[394];
			WeightsStore4[3] <= WeightsStore4[395];
			WeightsStore4[4] <= WeightsStore4[396];
			WeightsStore4[5] <= WeightsStore4[397];
			WeightsStore4[6] <= WeightsStore4[398];
			WeightsStore4[7] <= WeightsStore4[399];
			WeightsStore4[8] <= WeightsStore4[400];
			WeightsStore4[9] <= WeightsStore4[401];
			WeightsStore4[10] <= WeightsStore4[402];
			WeightsStore4[11] <= WeightsStore4[403];
			WeightsStore4[12] <= WeightsStore4[404];
			WeightsStore4[13] <= WeightsStore4[405];
			WeightsStore4[14] <= WeightsStore4[406];
			WeightsStore4[15] <= WeightsStore4[407];
			WeightsStore4[16] <= WeightsStore4[408];
			WeightsStore4[17] <= WeightsStore4[409];
			WeightsStore4[18] <= WeightsStore4[410];
			WeightsStore4[19] <= WeightsStore4[411];
			WeightsStore4[20] <= WeightsStore4[412];
			WeightsStore4[21] <= WeightsStore4[413];
			WeightsStore4[22] <= WeightsStore4[414];
			WeightsStore4[23] <= WeightsStore4[415];
			WeightsStore4[24] <= WeightsStore4[416];
			WeightsStore4[25] <= WeightsStore4[417];
			WeightsStore4[26] <= WeightsStore4[418];
			WeightsStore4[27] <= WeightsStore4[419];
			WeightsStore5[0] <= WeightsStore5[392];
			WeightsStore5[1] <= WeightsStore5[393];
			WeightsStore5[2] <= WeightsStore5[394];
			WeightsStore5[3] <= WeightsStore5[395];
			WeightsStore5[4] <= WeightsStore5[396];
			WeightsStore5[5] <= WeightsStore5[397];
			WeightsStore5[6] <= WeightsStore5[398];
			WeightsStore5[7] <= WeightsStore5[399];
			WeightsStore5[8] <= WeightsStore5[400];
			WeightsStore5[9] <= WeightsStore5[401];
			WeightsStore5[10] <= WeightsStore5[402];
			WeightsStore5[11] <= WeightsStore5[403];
			WeightsStore5[12] <= WeightsStore5[404];
			WeightsStore5[13] <= WeightsStore5[405];
			WeightsStore5[14] <= WeightsStore5[406];
			WeightsStore5[15] <= WeightsStore5[407];
			WeightsStore5[16] <= WeightsStore5[408];
			WeightsStore5[17] <= WeightsStore5[409];
			WeightsStore5[18] <= WeightsStore5[410];
			WeightsStore5[19] <= WeightsStore5[411];
			WeightsStore5[20] <= WeightsStore5[412];
			WeightsStore5[21] <= WeightsStore5[413];
			WeightsStore5[22] <= WeightsStore5[414];
			WeightsStore5[23] <= WeightsStore5[415];
			WeightsStore5[24] <= WeightsStore5[416];
			WeightsStore5[25] <= WeightsStore5[417];
			WeightsStore5[26] <= WeightsStore5[418];
			WeightsStore5[27] <= WeightsStore5[419];
			WeightsStore6[0] <= WeightsStore6[392];
			WeightsStore6[1] <= WeightsStore6[393];
			WeightsStore6[2] <= WeightsStore6[394];
			WeightsStore6[3] <= WeightsStore6[395];
			WeightsStore6[4] <= WeightsStore6[396];
			WeightsStore6[5] <= WeightsStore6[397];
			WeightsStore6[6] <= WeightsStore6[398];
			WeightsStore6[7] <= WeightsStore6[399];
			WeightsStore6[8] <= WeightsStore6[400];
			WeightsStore6[9] <= WeightsStore6[401];
			WeightsStore6[10] <= WeightsStore6[402];
			WeightsStore6[11] <= WeightsStore6[403];
			WeightsStore6[12] <= WeightsStore6[404];
			WeightsStore6[13] <= WeightsStore6[405];
			WeightsStore6[14] <= WeightsStore6[406];
			WeightsStore6[15] <= WeightsStore6[407];
			WeightsStore6[16] <= WeightsStore6[408];
			WeightsStore6[17] <= WeightsStore6[409];
			WeightsStore6[18] <= WeightsStore6[410];
			WeightsStore6[19] <= WeightsStore6[411];
			WeightsStore6[20] <= WeightsStore6[412];
			WeightsStore6[21] <= WeightsStore6[413];
			WeightsStore6[22] <= WeightsStore6[414];
			WeightsStore6[23] <= WeightsStore6[415];
			WeightsStore6[24] <= WeightsStore6[416];
			WeightsStore6[25] <= WeightsStore6[417];
			WeightsStore6[26] <= WeightsStore6[418];
			WeightsStore6[27] <= WeightsStore6[419];
			WeightsStore7[0] <= WeightsStore7[392];
			WeightsStore7[1] <= WeightsStore7[393];
			WeightsStore7[2] <= WeightsStore7[394];
			WeightsStore7[3] <= WeightsStore7[395];
			WeightsStore7[4] <= WeightsStore7[396];
			WeightsStore7[5] <= WeightsStore7[397];
			WeightsStore7[6] <= WeightsStore7[398];
			WeightsStore7[7] <= WeightsStore7[399];
			WeightsStore7[8] <= WeightsStore7[400];
			WeightsStore7[9] <= WeightsStore7[401];
			WeightsStore7[10] <= WeightsStore7[402];
			WeightsStore7[11] <= WeightsStore7[403];
			WeightsStore7[12] <= WeightsStore7[404];
			WeightsStore7[13] <= WeightsStore7[405];
			WeightsStore7[14] <= WeightsStore7[406];
			WeightsStore7[15] <= WeightsStore7[407];
			WeightsStore7[16] <= WeightsStore7[408];
			WeightsStore7[17] <= WeightsStore7[409];
			WeightsStore7[18] <= WeightsStore7[410];
			WeightsStore7[19] <= WeightsStore7[411];
			WeightsStore7[20] <= WeightsStore7[412];
			WeightsStore7[21] <= WeightsStore7[413];
			WeightsStore7[22] <= WeightsStore7[414];
			WeightsStore7[23] <= WeightsStore7[415];
			WeightsStore7[24] <= WeightsStore7[416];
			WeightsStore7[25] <= WeightsStore7[417];
			WeightsStore7[26] <= WeightsStore7[418];
			WeightsStore7[27] <= WeightsStore7[419];
			WeightsStore8[0] <= WeightsStore8[392];
			WeightsStore8[1] <= WeightsStore8[393];
			WeightsStore8[2] <= WeightsStore8[394];
			WeightsStore8[3] <= WeightsStore8[395];
			WeightsStore8[4] <= WeightsStore8[396];
			WeightsStore8[5] <= WeightsStore8[397];
			WeightsStore8[6] <= WeightsStore8[398];
			WeightsStore8[7] <= WeightsStore8[399];
			WeightsStore8[8] <= WeightsStore8[400];
			WeightsStore8[9] <= WeightsStore8[401];
			WeightsStore8[10] <= WeightsStore8[402];
			WeightsStore8[11] <= WeightsStore8[403];
			WeightsStore8[12] <= WeightsStore8[404];
			WeightsStore8[13] <= WeightsStore8[405];
			WeightsStore8[14] <= WeightsStore8[406];
			WeightsStore8[15] <= WeightsStore8[407];
			WeightsStore8[16] <= WeightsStore8[408];
			WeightsStore8[17] <= WeightsStore8[409];
			WeightsStore8[18] <= WeightsStore8[410];
			WeightsStore8[19] <= WeightsStore8[411];
			WeightsStore8[20] <= WeightsStore8[412];
			WeightsStore8[21] <= WeightsStore8[413];
			WeightsStore8[22] <= WeightsStore8[414];
			WeightsStore8[23] <= WeightsStore8[415];
			WeightsStore8[24] <= WeightsStore8[416];
			WeightsStore8[25] <= WeightsStore8[417];
			WeightsStore8[26] <= WeightsStore8[418];
			WeightsStore8[27] <= WeightsStore8[419];
			WeightsStore9[0] <= WeightsStore9[392];
			WeightsStore9[1] <= WeightsStore9[393];
			WeightsStore9[2] <= WeightsStore9[394];
			WeightsStore9[3] <= WeightsStore9[395];
			WeightsStore9[4] <= WeightsStore9[396];
			WeightsStore9[5] <= WeightsStore9[397];
			WeightsStore9[6] <= WeightsStore9[398];
			WeightsStore9[7] <= WeightsStore9[399];
			WeightsStore9[8] <= WeightsStore9[400];
			WeightsStore9[9] <= WeightsStore9[401];
			WeightsStore9[10] <= WeightsStore9[402];
			WeightsStore9[11] <= WeightsStore9[403];
			WeightsStore9[12] <= WeightsStore9[404];
			WeightsStore9[13] <= WeightsStore9[405];
			WeightsStore9[14] <= WeightsStore9[406];
			WeightsStore9[15] <= WeightsStore9[407];
			WeightsStore9[16] <= WeightsStore9[408];
			WeightsStore9[17] <= WeightsStore9[409];
			WeightsStore9[18] <= WeightsStore9[410];
			WeightsStore9[19] <= WeightsStore9[411];
			WeightsStore9[20] <= WeightsStore9[412];
			WeightsStore9[21] <= WeightsStore9[413];
			WeightsStore9[22] <= WeightsStore9[414];
			WeightsStore9[23] <= WeightsStore9[415];
			WeightsStore9[24] <= WeightsStore9[416];
			WeightsStore9[25] <= WeightsStore9[417];
			WeightsStore9[26] <= WeightsStore9[418];
			WeightsStore9[27] <= WeightsStore9[419];
		end else if(switchCounter == 32'd104)begin
			PixelsStore[0] <= PixelsStore[420];
			PixelsStore[1] <= PixelsStore[421];
			PixelsStore[2] <= PixelsStore[422];
			PixelsStore[3] <= PixelsStore[423];
			PixelsStore[4] <= PixelsStore[424];
			PixelsStore[5] <= PixelsStore[425];
			PixelsStore[6] <= PixelsStore[426];
			PixelsStore[7] <= PixelsStore[427];
			PixelsStore[8] <= PixelsStore[428];
			PixelsStore[9] <= PixelsStore[429];
			PixelsStore[10] <= PixelsStore[430];
			PixelsStore[11] <= PixelsStore[431];
			PixelsStore[12] <= PixelsStore[432];
			PixelsStore[13] <= PixelsStore[433];
			PixelsStore[14] <= PixelsStore[434];
			PixelsStore[15] <= PixelsStore[435];
			PixelsStore[16] <= PixelsStore[436];
			PixelsStore[17] <= PixelsStore[437];
			PixelsStore[18] <= PixelsStore[438];
			PixelsStore[19] <= PixelsStore[439];
			PixelsStore[20] <= PixelsStore[440];
			PixelsStore[21] <= PixelsStore[441];
			PixelsStore[22] <= PixelsStore[442];
			PixelsStore[23] <= PixelsStore[443];
			PixelsStore[24] <= PixelsStore[444];
			PixelsStore[25] <= PixelsStore[445];
			PixelsStore[26] <= PixelsStore[446];
			PixelsStore[27] <= PixelsStore[447];
			WeightsStore0[0] <= WeightsStore0[420];
			WeightsStore0[1] <= WeightsStore0[421];
			WeightsStore0[2] <= WeightsStore0[422];
			WeightsStore0[3] <= WeightsStore0[423];
			WeightsStore0[4] <= WeightsStore0[424];
			WeightsStore0[5] <= WeightsStore0[425];
			WeightsStore0[6] <= WeightsStore0[426];
			WeightsStore0[7] <= WeightsStore0[427];
			WeightsStore0[8] <= WeightsStore0[428];
			WeightsStore0[9] <= WeightsStore0[429];
			WeightsStore0[10] <= WeightsStore0[430];
			WeightsStore0[11] <= WeightsStore0[431];
			WeightsStore0[12] <= WeightsStore0[432];
			WeightsStore0[13] <= WeightsStore0[433];
			WeightsStore0[14] <= WeightsStore0[434];
			WeightsStore0[15] <= WeightsStore0[435];
			WeightsStore0[16] <= WeightsStore0[436];
			WeightsStore0[17] <= WeightsStore0[437];
			WeightsStore0[18] <= WeightsStore0[438];
			WeightsStore0[19] <= WeightsStore0[439];
			WeightsStore0[20] <= WeightsStore0[440];
			WeightsStore0[21] <= WeightsStore0[441];
			WeightsStore0[22] <= WeightsStore0[442];
			WeightsStore0[23] <= WeightsStore0[443];
			WeightsStore0[24] <= WeightsStore0[444];
			WeightsStore0[25] <= WeightsStore0[445];
			WeightsStore0[26] <= WeightsStore0[446];
			WeightsStore0[27] <= WeightsStore0[447];
			WeightsStore1[0] <= WeightsStore1[420];
			WeightsStore1[1] <= WeightsStore1[421];
			WeightsStore1[2] <= WeightsStore1[422];
			WeightsStore1[3] <= WeightsStore1[423];
			WeightsStore1[4] <= WeightsStore1[424];
			WeightsStore1[5] <= WeightsStore1[425];
			WeightsStore1[6] <= WeightsStore1[426];
			WeightsStore1[7] <= WeightsStore1[427];
			WeightsStore1[8] <= WeightsStore1[428];
			WeightsStore1[9] <= WeightsStore1[429];
			WeightsStore1[10] <= WeightsStore1[430];
			WeightsStore1[11] <= WeightsStore1[431];
			WeightsStore1[12] <= WeightsStore1[432];
			WeightsStore1[13] <= WeightsStore1[433];
			WeightsStore1[14] <= WeightsStore1[434];
			WeightsStore1[15] <= WeightsStore1[435];
			WeightsStore1[16] <= WeightsStore1[436];
			WeightsStore1[17] <= WeightsStore1[437];
			WeightsStore1[18] <= WeightsStore1[438];
			WeightsStore1[19] <= WeightsStore1[439];
			WeightsStore1[20] <= WeightsStore1[440];
			WeightsStore1[21] <= WeightsStore1[441];
			WeightsStore1[22] <= WeightsStore1[442];
			WeightsStore1[23] <= WeightsStore1[443];
			WeightsStore1[24] <= WeightsStore1[444];
			WeightsStore1[25] <= WeightsStore1[445];
			WeightsStore1[26] <= WeightsStore1[446];
			WeightsStore1[27] <= WeightsStore1[447];
			WeightsStore2[0] <= WeightsStore2[420];
			WeightsStore2[1] <= WeightsStore2[421];
			WeightsStore2[2] <= WeightsStore2[422];
			WeightsStore2[3] <= WeightsStore2[423];
			WeightsStore2[4] <= WeightsStore2[424];
			WeightsStore2[5] <= WeightsStore2[425];
			WeightsStore2[6] <= WeightsStore2[426];
			WeightsStore2[7] <= WeightsStore2[427];
			WeightsStore2[8] <= WeightsStore2[428];
			WeightsStore2[9] <= WeightsStore2[429];
			WeightsStore2[10] <= WeightsStore2[430];
			WeightsStore2[11] <= WeightsStore2[431];
			WeightsStore2[12] <= WeightsStore2[432];
			WeightsStore2[13] <= WeightsStore2[433];
			WeightsStore2[14] <= WeightsStore2[434];
			WeightsStore2[15] <= WeightsStore2[435];
			WeightsStore2[16] <= WeightsStore2[436];
			WeightsStore2[17] <= WeightsStore2[437];
			WeightsStore2[18] <= WeightsStore2[438];
			WeightsStore2[19] <= WeightsStore2[439];
			WeightsStore2[20] <= WeightsStore2[440];
			WeightsStore2[21] <= WeightsStore2[441];
			WeightsStore2[22] <= WeightsStore2[442];
			WeightsStore2[23] <= WeightsStore2[443];
			WeightsStore2[24] <= WeightsStore2[444];
			WeightsStore2[25] <= WeightsStore2[445];
			WeightsStore2[26] <= WeightsStore2[446];
			WeightsStore2[27] <= WeightsStore2[447];
			WeightsStore3[0] <= WeightsStore3[420];
			WeightsStore3[1] <= WeightsStore3[421];
			WeightsStore3[2] <= WeightsStore3[422];
			WeightsStore3[3] <= WeightsStore3[423];
			WeightsStore3[4] <= WeightsStore3[424];
			WeightsStore3[5] <= WeightsStore3[425];
			WeightsStore3[6] <= WeightsStore3[426];
			WeightsStore3[7] <= WeightsStore3[427];
			WeightsStore3[8] <= WeightsStore3[428];
			WeightsStore3[9] <= WeightsStore3[429];
			WeightsStore3[10] <= WeightsStore3[430];
			WeightsStore3[11] <= WeightsStore3[431];
			WeightsStore3[12] <= WeightsStore3[432];
			WeightsStore3[13] <= WeightsStore3[433];
			WeightsStore3[14] <= WeightsStore3[434];
			WeightsStore3[15] <= WeightsStore3[435];
			WeightsStore3[16] <= WeightsStore3[436];
			WeightsStore3[17] <= WeightsStore3[437];
			WeightsStore3[18] <= WeightsStore3[438];
			WeightsStore3[19] <= WeightsStore3[439];
			WeightsStore3[20] <= WeightsStore3[440];
			WeightsStore3[21] <= WeightsStore3[441];
			WeightsStore3[22] <= WeightsStore3[442];
			WeightsStore3[23] <= WeightsStore3[443];
			WeightsStore3[24] <= WeightsStore3[444];
			WeightsStore3[25] <= WeightsStore3[445];
			WeightsStore3[26] <= WeightsStore3[446];
			WeightsStore3[27] <= WeightsStore3[447];
			WeightsStore4[0] <= WeightsStore4[420];
			WeightsStore4[1] <= WeightsStore4[421];
			WeightsStore4[2] <= WeightsStore4[422];
			WeightsStore4[3] <= WeightsStore4[423];
			WeightsStore4[4] <= WeightsStore4[424];
			WeightsStore4[5] <= WeightsStore4[425];
			WeightsStore4[6] <= WeightsStore4[426];
			WeightsStore4[7] <= WeightsStore4[427];
			WeightsStore4[8] <= WeightsStore4[428];
			WeightsStore4[9] <= WeightsStore4[429];
			WeightsStore4[10] <= WeightsStore4[430];
			WeightsStore4[11] <= WeightsStore4[431];
			WeightsStore4[12] <= WeightsStore4[432];
			WeightsStore4[13] <= WeightsStore4[433];
			WeightsStore4[14] <= WeightsStore4[434];
			WeightsStore4[15] <= WeightsStore4[435];
			WeightsStore4[16] <= WeightsStore4[436];
			WeightsStore4[17] <= WeightsStore4[437];
			WeightsStore4[18] <= WeightsStore4[438];
			WeightsStore4[19] <= WeightsStore4[439];
			WeightsStore4[20] <= WeightsStore4[440];
			WeightsStore4[21] <= WeightsStore4[441];
			WeightsStore4[22] <= WeightsStore4[442];
			WeightsStore4[23] <= WeightsStore4[443];
			WeightsStore4[24] <= WeightsStore4[444];
			WeightsStore4[25] <= WeightsStore4[445];
			WeightsStore4[26] <= WeightsStore4[446];
			WeightsStore4[27] <= WeightsStore4[447];
			WeightsStore5[0] <= WeightsStore5[420];
			WeightsStore5[1] <= WeightsStore5[421];
			WeightsStore5[2] <= WeightsStore5[422];
			WeightsStore5[3] <= WeightsStore5[423];
			WeightsStore5[4] <= WeightsStore5[424];
			WeightsStore5[5] <= WeightsStore5[425];
			WeightsStore5[6] <= WeightsStore5[426];
			WeightsStore5[7] <= WeightsStore5[427];
			WeightsStore5[8] <= WeightsStore5[428];
			WeightsStore5[9] <= WeightsStore5[429];
			WeightsStore5[10] <= WeightsStore5[430];
			WeightsStore5[11] <= WeightsStore5[431];
			WeightsStore5[12] <= WeightsStore5[432];
			WeightsStore5[13] <= WeightsStore5[433];
			WeightsStore5[14] <= WeightsStore5[434];
			WeightsStore5[15] <= WeightsStore5[435];
			WeightsStore5[16] <= WeightsStore5[436];
			WeightsStore5[17] <= WeightsStore5[437];
			WeightsStore5[18] <= WeightsStore5[438];
			WeightsStore5[19] <= WeightsStore5[439];
			WeightsStore5[20] <= WeightsStore5[440];
			WeightsStore5[21] <= WeightsStore5[441];
			WeightsStore5[22] <= WeightsStore5[442];
			WeightsStore5[23] <= WeightsStore5[443];
			WeightsStore5[24] <= WeightsStore5[444];
			WeightsStore5[25] <= WeightsStore5[445];
			WeightsStore5[26] <= WeightsStore5[446];
			WeightsStore5[27] <= WeightsStore5[447];
			WeightsStore6[0] <= WeightsStore6[420];
			WeightsStore6[1] <= WeightsStore6[421];
			WeightsStore6[2] <= WeightsStore6[422];
			WeightsStore6[3] <= WeightsStore6[423];
			WeightsStore6[4] <= WeightsStore6[424];
			WeightsStore6[5] <= WeightsStore6[425];
			WeightsStore6[6] <= WeightsStore6[426];
			WeightsStore6[7] <= WeightsStore6[427];
			WeightsStore6[8] <= WeightsStore6[428];
			WeightsStore6[9] <= WeightsStore6[429];
			WeightsStore6[10] <= WeightsStore6[430];
			WeightsStore6[11] <= WeightsStore6[431];
			WeightsStore6[12] <= WeightsStore6[432];
			WeightsStore6[13] <= WeightsStore6[433];
			WeightsStore6[14] <= WeightsStore6[434];
			WeightsStore6[15] <= WeightsStore6[435];
			WeightsStore6[16] <= WeightsStore6[436];
			WeightsStore6[17] <= WeightsStore6[437];
			WeightsStore6[18] <= WeightsStore6[438];
			WeightsStore6[19] <= WeightsStore6[439];
			WeightsStore6[20] <= WeightsStore6[440];
			WeightsStore6[21] <= WeightsStore6[441];
			WeightsStore6[22] <= WeightsStore6[442];
			WeightsStore6[23] <= WeightsStore6[443];
			WeightsStore6[24] <= WeightsStore6[444];
			WeightsStore6[25] <= WeightsStore6[445];
			WeightsStore6[26] <= WeightsStore6[446];
			WeightsStore6[27] <= WeightsStore6[447];
			WeightsStore7[0] <= WeightsStore7[420];
			WeightsStore7[1] <= WeightsStore7[421];
			WeightsStore7[2] <= WeightsStore7[422];
			WeightsStore7[3] <= WeightsStore7[423];
			WeightsStore7[4] <= WeightsStore7[424];
			WeightsStore7[5] <= WeightsStore7[425];
			WeightsStore7[6] <= WeightsStore7[426];
			WeightsStore7[7] <= WeightsStore7[427];
			WeightsStore7[8] <= WeightsStore7[428];
			WeightsStore7[9] <= WeightsStore7[429];
			WeightsStore7[10] <= WeightsStore7[430];
			WeightsStore7[11] <= WeightsStore7[431];
			WeightsStore7[12] <= WeightsStore7[432];
			WeightsStore7[13] <= WeightsStore7[433];
			WeightsStore7[14] <= WeightsStore7[434];
			WeightsStore7[15] <= WeightsStore7[435];
			WeightsStore7[16] <= WeightsStore7[436];
			WeightsStore7[17] <= WeightsStore7[437];
			WeightsStore7[18] <= WeightsStore7[438];
			WeightsStore7[19] <= WeightsStore7[439];
			WeightsStore7[20] <= WeightsStore7[440];
			WeightsStore7[21] <= WeightsStore7[441];
			WeightsStore7[22] <= WeightsStore7[442];
			WeightsStore7[23] <= WeightsStore7[443];
			WeightsStore7[24] <= WeightsStore7[444];
			WeightsStore7[25] <= WeightsStore7[445];
			WeightsStore7[26] <= WeightsStore7[446];
			WeightsStore7[27] <= WeightsStore7[447];
			WeightsStore8[0] <= WeightsStore8[420];
			WeightsStore8[1] <= WeightsStore8[421];
			WeightsStore8[2] <= WeightsStore8[422];
			WeightsStore8[3] <= WeightsStore8[423];
			WeightsStore8[4] <= WeightsStore8[424];
			WeightsStore8[5] <= WeightsStore8[425];
			WeightsStore8[6] <= WeightsStore8[426];
			WeightsStore8[7] <= WeightsStore8[427];
			WeightsStore8[8] <= WeightsStore8[428];
			WeightsStore8[9] <= WeightsStore8[429];
			WeightsStore8[10] <= WeightsStore8[430];
			WeightsStore8[11] <= WeightsStore8[431];
			WeightsStore8[12] <= WeightsStore8[432];
			WeightsStore8[13] <= WeightsStore8[433];
			WeightsStore8[14] <= WeightsStore8[434];
			WeightsStore8[15] <= WeightsStore8[435];
			WeightsStore8[16] <= WeightsStore8[436];
			WeightsStore8[17] <= WeightsStore8[437];
			WeightsStore8[18] <= WeightsStore8[438];
			WeightsStore8[19] <= WeightsStore8[439];
			WeightsStore8[20] <= WeightsStore8[440];
			WeightsStore8[21] <= WeightsStore8[441];
			WeightsStore8[22] <= WeightsStore8[442];
			WeightsStore8[23] <= WeightsStore8[443];
			WeightsStore8[24] <= WeightsStore8[444];
			WeightsStore8[25] <= WeightsStore8[445];
			WeightsStore8[26] <= WeightsStore8[446];
			WeightsStore8[27] <= WeightsStore8[447];
			WeightsStore9[0] <= WeightsStore9[420];
			WeightsStore9[1] <= WeightsStore9[421];
			WeightsStore9[2] <= WeightsStore9[422];
			WeightsStore9[3] <= WeightsStore9[423];
			WeightsStore9[4] <= WeightsStore9[424];
			WeightsStore9[5] <= WeightsStore9[425];
			WeightsStore9[6] <= WeightsStore9[426];
			WeightsStore9[7] <= WeightsStore9[427];
			WeightsStore9[8] <= WeightsStore9[428];
			WeightsStore9[9] <= WeightsStore9[429];
			WeightsStore9[10] <= WeightsStore9[430];
			WeightsStore9[11] <= WeightsStore9[431];
			WeightsStore9[12] <= WeightsStore9[432];
			WeightsStore9[13] <= WeightsStore9[433];
			WeightsStore9[14] <= WeightsStore9[434];
			WeightsStore9[15] <= WeightsStore9[435];
			WeightsStore9[16] <= WeightsStore9[436];
			WeightsStore9[17] <= WeightsStore9[437];
			WeightsStore9[18] <= WeightsStore9[438];
			WeightsStore9[19] <= WeightsStore9[439];
			WeightsStore9[20] <= WeightsStore9[440];
			WeightsStore9[21] <= WeightsStore9[441];
			WeightsStore9[22] <= WeightsStore9[442];
			WeightsStore9[23] <= WeightsStore9[443];
			WeightsStore9[24] <= WeightsStore9[444];
			WeightsStore9[25] <= WeightsStore9[445];
			WeightsStore9[26] <= WeightsStore9[446];
			WeightsStore9[27] <= WeightsStore9[447];
		end else if(switchCounter == 32'd111)begin
			PixelsStore[0] <= PixelsStore[448];
			PixelsStore[1] <= PixelsStore[449];
			PixelsStore[2] <= PixelsStore[450];
			PixelsStore[3] <= PixelsStore[451];
			PixelsStore[4] <= PixelsStore[452];
			PixelsStore[5] <= PixelsStore[453];
			PixelsStore[6] <= PixelsStore[454];
			PixelsStore[7] <= PixelsStore[455];
			PixelsStore[8] <= PixelsStore[456];
			PixelsStore[9] <= PixelsStore[457];
			PixelsStore[10] <= PixelsStore[458];
			PixelsStore[11] <= PixelsStore[459];
			PixelsStore[12] <= PixelsStore[460];
			PixelsStore[13] <= PixelsStore[461];
			PixelsStore[14] <= PixelsStore[462];
			PixelsStore[15] <= PixelsStore[463];
			PixelsStore[16] <= PixelsStore[464];
			PixelsStore[17] <= PixelsStore[465];
			PixelsStore[18] <= PixelsStore[466];
			PixelsStore[19] <= PixelsStore[467];
			PixelsStore[20] <= PixelsStore[468];
			PixelsStore[21] <= PixelsStore[469];
			PixelsStore[22] <= PixelsStore[470];
			PixelsStore[23] <= PixelsStore[471];
			PixelsStore[24] <= PixelsStore[472];
			PixelsStore[25] <= PixelsStore[473];
			PixelsStore[26] <= PixelsStore[474];
			PixelsStore[27] <= PixelsStore[475];
			WeightsStore0[0] <= WeightsStore0[448];
			WeightsStore0[1] <= WeightsStore0[449];
			WeightsStore0[2] <= WeightsStore0[450];
			WeightsStore0[3] <= WeightsStore0[451];
			WeightsStore0[4] <= WeightsStore0[452];
			WeightsStore0[5] <= WeightsStore0[453];
			WeightsStore0[6] <= WeightsStore0[454];
			WeightsStore0[7] <= WeightsStore0[455];
			WeightsStore0[8] <= WeightsStore0[456];
			WeightsStore0[9] <= WeightsStore0[457];
			WeightsStore0[10] <= WeightsStore0[458];
			WeightsStore0[11] <= WeightsStore0[459];
			WeightsStore0[12] <= WeightsStore0[460];
			WeightsStore0[13] <= WeightsStore0[461];
			WeightsStore0[14] <= WeightsStore0[462];
			WeightsStore0[15] <= WeightsStore0[463];
			WeightsStore0[16] <= WeightsStore0[464];
			WeightsStore0[17] <= WeightsStore0[465];
			WeightsStore0[18] <= WeightsStore0[466];
			WeightsStore0[19] <= WeightsStore0[467];
			WeightsStore0[20] <= WeightsStore0[468];
			WeightsStore0[21] <= WeightsStore0[469];
			WeightsStore0[22] <= WeightsStore0[470];
			WeightsStore0[23] <= WeightsStore0[471];
			WeightsStore0[24] <= WeightsStore0[472];
			WeightsStore0[25] <= WeightsStore0[473];
			WeightsStore0[26] <= WeightsStore0[474];
			WeightsStore0[27] <= WeightsStore0[475];
			WeightsStore1[0] <= WeightsStore1[448];
			WeightsStore1[1] <= WeightsStore1[449];
			WeightsStore1[2] <= WeightsStore1[450];
			WeightsStore1[3] <= WeightsStore1[451];
			WeightsStore1[4] <= WeightsStore1[452];
			WeightsStore1[5] <= WeightsStore1[453];
			WeightsStore1[6] <= WeightsStore1[454];
			WeightsStore1[7] <= WeightsStore1[455];
			WeightsStore1[8] <= WeightsStore1[456];
			WeightsStore1[9] <= WeightsStore1[457];
			WeightsStore1[10] <= WeightsStore1[458];
			WeightsStore1[11] <= WeightsStore1[459];
			WeightsStore1[12] <= WeightsStore1[460];
			WeightsStore1[13] <= WeightsStore1[461];
			WeightsStore1[14] <= WeightsStore1[462];
			WeightsStore1[15] <= WeightsStore1[463];
			WeightsStore1[16] <= WeightsStore1[464];
			WeightsStore1[17] <= WeightsStore1[465];
			WeightsStore1[18] <= WeightsStore1[466];
			WeightsStore1[19] <= WeightsStore1[467];
			WeightsStore1[20] <= WeightsStore1[468];
			WeightsStore1[21] <= WeightsStore1[469];
			WeightsStore1[22] <= WeightsStore1[470];
			WeightsStore1[23] <= WeightsStore1[471];
			WeightsStore1[24] <= WeightsStore1[472];
			WeightsStore1[25] <= WeightsStore1[473];
			WeightsStore1[26] <= WeightsStore1[474];
			WeightsStore1[27] <= WeightsStore1[475];
			WeightsStore2[0] <= WeightsStore2[448];
			WeightsStore2[1] <= WeightsStore2[449];
			WeightsStore2[2] <= WeightsStore2[450];
			WeightsStore2[3] <= WeightsStore2[451];
			WeightsStore2[4] <= WeightsStore2[452];
			WeightsStore2[5] <= WeightsStore2[453];
			WeightsStore2[6] <= WeightsStore2[454];
			WeightsStore2[7] <= WeightsStore2[455];
			WeightsStore2[8] <= WeightsStore2[456];
			WeightsStore2[9] <= WeightsStore2[457];
			WeightsStore2[10] <= WeightsStore2[458];
			WeightsStore2[11] <= WeightsStore2[459];
			WeightsStore2[12] <= WeightsStore2[460];
			WeightsStore2[13] <= WeightsStore2[461];
			WeightsStore2[14] <= WeightsStore2[462];
			WeightsStore2[15] <= WeightsStore2[463];
			WeightsStore2[16] <= WeightsStore2[464];
			WeightsStore2[17] <= WeightsStore2[465];
			WeightsStore2[18] <= WeightsStore2[466];
			WeightsStore2[19] <= WeightsStore2[467];
			WeightsStore2[20] <= WeightsStore2[468];
			WeightsStore2[21] <= WeightsStore2[469];
			WeightsStore2[22] <= WeightsStore2[470];
			WeightsStore2[23] <= WeightsStore2[471];
			WeightsStore2[24] <= WeightsStore2[472];
			WeightsStore2[25] <= WeightsStore2[473];
			WeightsStore2[26] <= WeightsStore2[474];
			WeightsStore2[27] <= WeightsStore2[475];
			WeightsStore3[0] <= WeightsStore3[448];
			WeightsStore3[1] <= WeightsStore3[449];
			WeightsStore3[2] <= WeightsStore3[450];
			WeightsStore3[3] <= WeightsStore3[451];
			WeightsStore3[4] <= WeightsStore3[452];
			WeightsStore3[5] <= WeightsStore3[453];
			WeightsStore3[6] <= WeightsStore3[454];
			WeightsStore3[7] <= WeightsStore3[455];
			WeightsStore3[8] <= WeightsStore3[456];
			WeightsStore3[9] <= WeightsStore3[457];
			WeightsStore3[10] <= WeightsStore3[458];
			WeightsStore3[11] <= WeightsStore3[459];
			WeightsStore3[12] <= WeightsStore3[460];
			WeightsStore3[13] <= WeightsStore3[461];
			WeightsStore3[14] <= WeightsStore3[462];
			WeightsStore3[15] <= WeightsStore3[463];
			WeightsStore3[16] <= WeightsStore3[464];
			WeightsStore3[17] <= WeightsStore3[465];
			WeightsStore3[18] <= WeightsStore3[466];
			WeightsStore3[19] <= WeightsStore3[467];
			WeightsStore3[20] <= WeightsStore3[468];
			WeightsStore3[21] <= WeightsStore3[469];
			WeightsStore3[22] <= WeightsStore3[470];
			WeightsStore3[23] <= WeightsStore3[471];
			WeightsStore3[24] <= WeightsStore3[472];
			WeightsStore3[25] <= WeightsStore3[473];
			WeightsStore3[26] <= WeightsStore3[474];
			WeightsStore3[27] <= WeightsStore3[475];
			WeightsStore4[0] <= WeightsStore4[448];
			WeightsStore4[1] <= WeightsStore4[449];
			WeightsStore4[2] <= WeightsStore4[450];
			WeightsStore4[3] <= WeightsStore4[451];
			WeightsStore4[4] <= WeightsStore4[452];
			WeightsStore4[5] <= WeightsStore4[453];
			WeightsStore4[6] <= WeightsStore4[454];
			WeightsStore4[7] <= WeightsStore4[455];
			WeightsStore4[8] <= WeightsStore4[456];
			WeightsStore4[9] <= WeightsStore4[457];
			WeightsStore4[10] <= WeightsStore4[458];
			WeightsStore4[11] <= WeightsStore4[459];
			WeightsStore4[12] <= WeightsStore4[460];
			WeightsStore4[13] <= WeightsStore4[461];
			WeightsStore4[14] <= WeightsStore4[462];
			WeightsStore4[15] <= WeightsStore4[463];
			WeightsStore4[16] <= WeightsStore4[464];
			WeightsStore4[17] <= WeightsStore4[465];
			WeightsStore4[18] <= WeightsStore4[466];
			WeightsStore4[19] <= WeightsStore4[467];
			WeightsStore4[20] <= WeightsStore4[468];
			WeightsStore4[21] <= WeightsStore4[469];
			WeightsStore4[22] <= WeightsStore4[470];
			WeightsStore4[23] <= WeightsStore4[471];
			WeightsStore4[24] <= WeightsStore4[472];
			WeightsStore4[25] <= WeightsStore4[473];
			WeightsStore4[26] <= WeightsStore4[474];
			WeightsStore4[27] <= WeightsStore4[475];
			WeightsStore5[0] <= WeightsStore5[448];
			WeightsStore5[1] <= WeightsStore5[449];
			WeightsStore5[2] <= WeightsStore5[450];
			WeightsStore5[3] <= WeightsStore5[451];
			WeightsStore5[4] <= WeightsStore5[452];
			WeightsStore5[5] <= WeightsStore5[453];
			WeightsStore5[6] <= WeightsStore5[454];
			WeightsStore5[7] <= WeightsStore5[455];
			WeightsStore5[8] <= WeightsStore5[456];
			WeightsStore5[9] <= WeightsStore5[457];
			WeightsStore5[10] <= WeightsStore5[458];
			WeightsStore5[11] <= WeightsStore5[459];
			WeightsStore5[12] <= WeightsStore5[460];
			WeightsStore5[13] <= WeightsStore5[461];
			WeightsStore5[14] <= WeightsStore5[462];
			WeightsStore5[15] <= WeightsStore5[463];
			WeightsStore5[16] <= WeightsStore5[464];
			WeightsStore5[17] <= WeightsStore5[465];
			WeightsStore5[18] <= WeightsStore5[466];
			WeightsStore5[19] <= WeightsStore5[467];
			WeightsStore5[20] <= WeightsStore5[468];
			WeightsStore5[21] <= WeightsStore5[469];
			WeightsStore5[22] <= WeightsStore5[470];
			WeightsStore5[23] <= WeightsStore5[471];
			WeightsStore5[24] <= WeightsStore5[472];
			WeightsStore5[25] <= WeightsStore5[473];
			WeightsStore5[26] <= WeightsStore5[474];
			WeightsStore5[27] <= WeightsStore5[475];
			WeightsStore6[0] <= WeightsStore6[448];
			WeightsStore6[1] <= WeightsStore6[449];
			WeightsStore6[2] <= WeightsStore6[450];
			WeightsStore6[3] <= WeightsStore6[451];
			WeightsStore6[4] <= WeightsStore6[452];
			WeightsStore6[5] <= WeightsStore6[453];
			WeightsStore6[6] <= WeightsStore6[454];
			WeightsStore6[7] <= WeightsStore6[455];
			WeightsStore6[8] <= WeightsStore6[456];
			WeightsStore6[9] <= WeightsStore6[457];
			WeightsStore6[10] <= WeightsStore6[458];
			WeightsStore6[11] <= WeightsStore6[459];
			WeightsStore6[12] <= WeightsStore6[460];
			WeightsStore6[13] <= WeightsStore6[461];
			WeightsStore6[14] <= WeightsStore6[462];
			WeightsStore6[15] <= WeightsStore6[463];
			WeightsStore6[16] <= WeightsStore6[464];
			WeightsStore6[17] <= WeightsStore6[465];
			WeightsStore6[18] <= WeightsStore6[466];
			WeightsStore6[19] <= WeightsStore6[467];
			WeightsStore6[20] <= WeightsStore6[468];
			WeightsStore6[21] <= WeightsStore6[469];
			WeightsStore6[22] <= WeightsStore6[470];
			WeightsStore6[23] <= WeightsStore6[471];
			WeightsStore6[24] <= WeightsStore6[472];
			WeightsStore6[25] <= WeightsStore6[473];
			WeightsStore6[26] <= WeightsStore6[474];
			WeightsStore6[27] <= WeightsStore6[475];
			WeightsStore7[0] <= WeightsStore7[448];
			WeightsStore7[1] <= WeightsStore7[449];
			WeightsStore7[2] <= WeightsStore7[450];
			WeightsStore7[3] <= WeightsStore7[451];
			WeightsStore7[4] <= WeightsStore7[452];
			WeightsStore7[5] <= WeightsStore7[453];
			WeightsStore7[6] <= WeightsStore7[454];
			WeightsStore7[7] <= WeightsStore7[455];
			WeightsStore7[8] <= WeightsStore7[456];
			WeightsStore7[9] <= WeightsStore7[457];
			WeightsStore7[10] <= WeightsStore7[458];
			WeightsStore7[11] <= WeightsStore7[459];
			WeightsStore7[12] <= WeightsStore7[460];
			WeightsStore7[13] <= WeightsStore7[461];
			WeightsStore7[14] <= WeightsStore7[462];
			WeightsStore7[15] <= WeightsStore7[463];
			WeightsStore7[16] <= WeightsStore7[464];
			WeightsStore7[17] <= WeightsStore7[465];
			WeightsStore7[18] <= WeightsStore7[466];
			WeightsStore7[19] <= WeightsStore7[467];
			WeightsStore7[20] <= WeightsStore7[468];
			WeightsStore7[21] <= WeightsStore7[469];
			WeightsStore7[22] <= WeightsStore7[470];
			WeightsStore7[23] <= WeightsStore7[471];
			WeightsStore7[24] <= WeightsStore7[472];
			WeightsStore7[25] <= WeightsStore7[473];
			WeightsStore7[26] <= WeightsStore7[474];
			WeightsStore7[27] <= WeightsStore7[475];
			WeightsStore8[0] <= WeightsStore8[448];
			WeightsStore8[1] <= WeightsStore8[449];
			WeightsStore8[2] <= WeightsStore8[450];
			WeightsStore8[3] <= WeightsStore8[451];
			WeightsStore8[4] <= WeightsStore8[452];
			WeightsStore8[5] <= WeightsStore8[453];
			WeightsStore8[6] <= WeightsStore8[454];
			WeightsStore8[7] <= WeightsStore8[455];
			WeightsStore8[8] <= WeightsStore8[456];
			WeightsStore8[9] <= WeightsStore8[457];
			WeightsStore8[10] <= WeightsStore8[458];
			WeightsStore8[11] <= WeightsStore8[459];
			WeightsStore8[12] <= WeightsStore8[460];
			WeightsStore8[13] <= WeightsStore8[461];
			WeightsStore8[14] <= WeightsStore8[462];
			WeightsStore8[15] <= WeightsStore8[463];
			WeightsStore8[16] <= WeightsStore8[464];
			WeightsStore8[17] <= WeightsStore8[465];
			WeightsStore8[18] <= WeightsStore8[466];
			WeightsStore8[19] <= WeightsStore8[467];
			WeightsStore8[20] <= WeightsStore8[468];
			WeightsStore8[21] <= WeightsStore8[469];
			WeightsStore8[22] <= WeightsStore8[470];
			WeightsStore8[23] <= WeightsStore8[471];
			WeightsStore8[24] <= WeightsStore8[472];
			WeightsStore8[25] <= WeightsStore8[473];
			WeightsStore8[26] <= WeightsStore8[474];
			WeightsStore8[27] <= WeightsStore8[475];
			WeightsStore9[0] <= WeightsStore9[448];
			WeightsStore9[1] <= WeightsStore9[449];
			WeightsStore9[2] <= WeightsStore9[450];
			WeightsStore9[3] <= WeightsStore9[451];
			WeightsStore9[4] <= WeightsStore9[452];
			WeightsStore9[5] <= WeightsStore9[453];
			WeightsStore9[6] <= WeightsStore9[454];
			WeightsStore9[7] <= WeightsStore9[455];
			WeightsStore9[8] <= WeightsStore9[456];
			WeightsStore9[9] <= WeightsStore9[457];
			WeightsStore9[10] <= WeightsStore9[458];
			WeightsStore9[11] <= WeightsStore9[459];
			WeightsStore9[12] <= WeightsStore9[460];
			WeightsStore9[13] <= WeightsStore9[461];
			WeightsStore9[14] <= WeightsStore9[462];
			WeightsStore9[15] <= WeightsStore9[463];
			WeightsStore9[16] <= WeightsStore9[464];
			WeightsStore9[17] <= WeightsStore9[465];
			WeightsStore9[18] <= WeightsStore9[466];
			WeightsStore9[19] <= WeightsStore9[467];
			WeightsStore9[20] <= WeightsStore9[468];
			WeightsStore9[21] <= WeightsStore9[469];
			WeightsStore9[22] <= WeightsStore9[470];
			WeightsStore9[23] <= WeightsStore9[471];
			WeightsStore9[24] <= WeightsStore9[472];
			WeightsStore9[25] <= WeightsStore9[473];
			WeightsStore9[26] <= WeightsStore9[474];
			WeightsStore9[27] <= WeightsStore9[475];
		end else if(switchCounter == 32'd118)begin
			PixelsStore[0] <= PixelsStore[476];
			PixelsStore[1] <= PixelsStore[477];
			PixelsStore[2] <= PixelsStore[478];
			PixelsStore[3] <= PixelsStore[479];
			PixelsStore[4] <= PixelsStore[480];
			PixelsStore[5] <= PixelsStore[481];
			PixelsStore[6] <= PixelsStore[482];
			PixelsStore[7] <= PixelsStore[483];
			PixelsStore[8] <= PixelsStore[484];
			PixelsStore[9] <= PixelsStore[485];
			PixelsStore[10] <= PixelsStore[486];
			PixelsStore[11] <= PixelsStore[487];
			PixelsStore[12] <= PixelsStore[488];
			PixelsStore[13] <= PixelsStore[489];
			PixelsStore[14] <= PixelsStore[490];
			PixelsStore[15] <= PixelsStore[491];
			PixelsStore[16] <= PixelsStore[492];
			PixelsStore[17] <= PixelsStore[493];
			PixelsStore[18] <= PixelsStore[494];
			PixelsStore[19] <= PixelsStore[495];
			PixelsStore[20] <= PixelsStore[496];
			PixelsStore[21] <= PixelsStore[497];
			PixelsStore[22] <= PixelsStore[498];
			PixelsStore[23] <= PixelsStore[499];
			PixelsStore[24] <= PixelsStore[500];
			PixelsStore[25] <= PixelsStore[501];
			PixelsStore[26] <= PixelsStore[502];
			PixelsStore[27] <= PixelsStore[503];
			WeightsStore0[0] <= WeightsStore0[476];
			WeightsStore0[1] <= WeightsStore0[477];
			WeightsStore0[2] <= WeightsStore0[478];
			WeightsStore0[3] <= WeightsStore0[479];
			WeightsStore0[4] <= WeightsStore0[480];
			WeightsStore0[5] <= WeightsStore0[481];
			WeightsStore0[6] <= WeightsStore0[482];
			WeightsStore0[7] <= WeightsStore0[483];
			WeightsStore0[8] <= WeightsStore0[484];
			WeightsStore0[9] <= WeightsStore0[485];
			WeightsStore0[10] <= WeightsStore0[486];
			WeightsStore0[11] <= WeightsStore0[487];
			WeightsStore0[12] <= WeightsStore0[488];
			WeightsStore0[13] <= WeightsStore0[489];
			WeightsStore0[14] <= WeightsStore0[490];
			WeightsStore0[15] <= WeightsStore0[491];
			WeightsStore0[16] <= WeightsStore0[492];
			WeightsStore0[17] <= WeightsStore0[493];
			WeightsStore0[18] <= WeightsStore0[494];
			WeightsStore0[19] <= WeightsStore0[495];
			WeightsStore0[20] <= WeightsStore0[496];
			WeightsStore0[21] <= WeightsStore0[497];
			WeightsStore0[22] <= WeightsStore0[498];
			WeightsStore0[23] <= WeightsStore0[499];
			WeightsStore0[24] <= WeightsStore0[500];
			WeightsStore0[25] <= WeightsStore0[501];
			WeightsStore0[26] <= WeightsStore0[502];
			WeightsStore0[27] <= WeightsStore0[503];
			WeightsStore1[0] <= WeightsStore1[476];
			WeightsStore1[1] <= WeightsStore1[477];
			WeightsStore1[2] <= WeightsStore1[478];
			WeightsStore1[3] <= WeightsStore1[479];
			WeightsStore1[4] <= WeightsStore1[480];
			WeightsStore1[5] <= WeightsStore1[481];
			WeightsStore1[6] <= WeightsStore1[482];
			WeightsStore1[7] <= WeightsStore1[483];
			WeightsStore1[8] <= WeightsStore1[484];
			WeightsStore1[9] <= WeightsStore1[485];
			WeightsStore1[10] <= WeightsStore1[486];
			WeightsStore1[11] <= WeightsStore1[487];
			WeightsStore1[12] <= WeightsStore1[488];
			WeightsStore1[13] <= WeightsStore1[489];
			WeightsStore1[14] <= WeightsStore1[490];
			WeightsStore1[15] <= WeightsStore1[491];
			WeightsStore1[16] <= WeightsStore1[492];
			WeightsStore1[17] <= WeightsStore1[493];
			WeightsStore1[18] <= WeightsStore1[494];
			WeightsStore1[19] <= WeightsStore1[495];
			WeightsStore1[20] <= WeightsStore1[496];
			WeightsStore1[21] <= WeightsStore1[497];
			WeightsStore1[22] <= WeightsStore1[498];
			WeightsStore1[23] <= WeightsStore1[499];
			WeightsStore1[24] <= WeightsStore1[500];
			WeightsStore1[25] <= WeightsStore1[501];
			WeightsStore1[26] <= WeightsStore1[502];
			WeightsStore1[27] <= WeightsStore1[503];
			WeightsStore2[0] <= WeightsStore2[476];
			WeightsStore2[1] <= WeightsStore2[477];
			WeightsStore2[2] <= WeightsStore2[478];
			WeightsStore2[3] <= WeightsStore2[479];
			WeightsStore2[4] <= WeightsStore2[480];
			WeightsStore2[5] <= WeightsStore2[481];
			WeightsStore2[6] <= WeightsStore2[482];
			WeightsStore2[7] <= WeightsStore2[483];
			WeightsStore2[8] <= WeightsStore2[484];
			WeightsStore2[9] <= WeightsStore2[485];
			WeightsStore2[10] <= WeightsStore2[486];
			WeightsStore2[11] <= WeightsStore2[487];
			WeightsStore2[12] <= WeightsStore2[488];
			WeightsStore2[13] <= WeightsStore2[489];
			WeightsStore2[14] <= WeightsStore2[490];
			WeightsStore2[15] <= WeightsStore2[491];
			WeightsStore2[16] <= WeightsStore2[492];
			WeightsStore2[17] <= WeightsStore2[493];
			WeightsStore2[18] <= WeightsStore2[494];
			WeightsStore2[19] <= WeightsStore2[495];
			WeightsStore2[20] <= WeightsStore2[496];
			WeightsStore2[21] <= WeightsStore2[497];
			WeightsStore2[22] <= WeightsStore2[498];
			WeightsStore2[23] <= WeightsStore2[499];
			WeightsStore2[24] <= WeightsStore2[500];
			WeightsStore2[25] <= WeightsStore2[501];
			WeightsStore2[26] <= WeightsStore2[502];
			WeightsStore2[27] <= WeightsStore2[503];
			WeightsStore3[0] <= WeightsStore3[476];
			WeightsStore3[1] <= WeightsStore3[477];
			WeightsStore3[2] <= WeightsStore3[478];
			WeightsStore3[3] <= WeightsStore3[479];
			WeightsStore3[4] <= WeightsStore3[480];
			WeightsStore3[5] <= WeightsStore3[481];
			WeightsStore3[6] <= WeightsStore3[482];
			WeightsStore3[7] <= WeightsStore3[483];
			WeightsStore3[8] <= WeightsStore3[484];
			WeightsStore3[9] <= WeightsStore3[485];
			WeightsStore3[10] <= WeightsStore3[486];
			WeightsStore3[11] <= WeightsStore3[487];
			WeightsStore3[12] <= WeightsStore3[488];
			WeightsStore3[13] <= WeightsStore3[489];
			WeightsStore3[14] <= WeightsStore3[490];
			WeightsStore3[15] <= WeightsStore3[491];
			WeightsStore3[16] <= WeightsStore3[492];
			WeightsStore3[17] <= WeightsStore3[493];
			WeightsStore3[18] <= WeightsStore3[494];
			WeightsStore3[19] <= WeightsStore3[495];
			WeightsStore3[20] <= WeightsStore3[496];
			WeightsStore3[21] <= WeightsStore3[497];
			WeightsStore3[22] <= WeightsStore3[498];
			WeightsStore3[23] <= WeightsStore3[499];
			WeightsStore3[24] <= WeightsStore3[500];
			WeightsStore3[25] <= WeightsStore3[501];
			WeightsStore3[26] <= WeightsStore3[502];
			WeightsStore3[27] <= WeightsStore3[503];
			WeightsStore4[0] <= WeightsStore4[476];
			WeightsStore4[1] <= WeightsStore4[477];
			WeightsStore4[2] <= WeightsStore4[478];
			WeightsStore4[3] <= WeightsStore4[479];
			WeightsStore4[4] <= WeightsStore4[480];
			WeightsStore4[5] <= WeightsStore4[481];
			WeightsStore4[6] <= WeightsStore4[482];
			WeightsStore4[7] <= WeightsStore4[483];
			WeightsStore4[8] <= WeightsStore4[484];
			WeightsStore4[9] <= WeightsStore4[485];
			WeightsStore4[10] <= WeightsStore4[486];
			WeightsStore4[11] <= WeightsStore4[487];
			WeightsStore4[12] <= WeightsStore4[488];
			WeightsStore4[13] <= WeightsStore4[489];
			WeightsStore4[14] <= WeightsStore4[490];
			WeightsStore4[15] <= WeightsStore4[491];
			WeightsStore4[16] <= WeightsStore4[492];
			WeightsStore4[17] <= WeightsStore4[493];
			WeightsStore4[18] <= WeightsStore4[494];
			WeightsStore4[19] <= WeightsStore4[495];
			WeightsStore4[20] <= WeightsStore4[496];
			WeightsStore4[21] <= WeightsStore4[497];
			WeightsStore4[22] <= WeightsStore4[498];
			WeightsStore4[23] <= WeightsStore4[499];
			WeightsStore4[24] <= WeightsStore4[500];
			WeightsStore4[25] <= WeightsStore4[501];
			WeightsStore4[26] <= WeightsStore4[502];
			WeightsStore4[27] <= WeightsStore4[503];
			WeightsStore5[0] <= WeightsStore5[476];
			WeightsStore5[1] <= WeightsStore5[477];
			WeightsStore5[2] <= WeightsStore5[478];
			WeightsStore5[3] <= WeightsStore5[479];
			WeightsStore5[4] <= WeightsStore5[480];
			WeightsStore5[5] <= WeightsStore5[481];
			WeightsStore5[6] <= WeightsStore5[482];
			WeightsStore5[7] <= WeightsStore5[483];
			WeightsStore5[8] <= WeightsStore5[484];
			WeightsStore5[9] <= WeightsStore5[485];
			WeightsStore5[10] <= WeightsStore5[486];
			WeightsStore5[11] <= WeightsStore5[487];
			WeightsStore5[12] <= WeightsStore5[488];
			WeightsStore5[13] <= WeightsStore5[489];
			WeightsStore5[14] <= WeightsStore5[490];
			WeightsStore5[15] <= WeightsStore5[491];
			WeightsStore5[16] <= WeightsStore5[492];
			WeightsStore5[17] <= WeightsStore5[493];
			WeightsStore5[18] <= WeightsStore5[494];
			WeightsStore5[19] <= WeightsStore5[495];
			WeightsStore5[20] <= WeightsStore5[496];
			WeightsStore5[21] <= WeightsStore5[497];
			WeightsStore5[22] <= WeightsStore5[498];
			WeightsStore5[23] <= WeightsStore5[499];
			WeightsStore5[24] <= WeightsStore5[500];
			WeightsStore5[25] <= WeightsStore5[501];
			WeightsStore5[26] <= WeightsStore5[502];
			WeightsStore5[27] <= WeightsStore5[503];
			WeightsStore6[0] <= WeightsStore6[476];
			WeightsStore6[1] <= WeightsStore6[477];
			WeightsStore6[2] <= WeightsStore6[478];
			WeightsStore6[3] <= WeightsStore6[479];
			WeightsStore6[4] <= WeightsStore6[480];
			WeightsStore6[5] <= WeightsStore6[481];
			WeightsStore6[6] <= WeightsStore6[482];
			WeightsStore6[7] <= WeightsStore6[483];
			WeightsStore6[8] <= WeightsStore6[484];
			WeightsStore6[9] <= WeightsStore6[485];
			WeightsStore6[10] <= WeightsStore6[486];
			WeightsStore6[11] <= WeightsStore6[487];
			WeightsStore6[12] <= WeightsStore6[488];
			WeightsStore6[13] <= WeightsStore6[489];
			WeightsStore6[14] <= WeightsStore6[490];
			WeightsStore6[15] <= WeightsStore6[491];
			WeightsStore6[16] <= WeightsStore6[492];
			WeightsStore6[17] <= WeightsStore6[493];
			WeightsStore6[18] <= WeightsStore6[494];
			WeightsStore6[19] <= WeightsStore6[495];
			WeightsStore6[20] <= WeightsStore6[496];
			WeightsStore6[21] <= WeightsStore6[497];
			WeightsStore6[22] <= WeightsStore6[498];
			WeightsStore6[23] <= WeightsStore6[499];
			WeightsStore6[24] <= WeightsStore6[500];
			WeightsStore6[25] <= WeightsStore6[501];
			WeightsStore6[26] <= WeightsStore6[502];
			WeightsStore6[27] <= WeightsStore6[503];
			WeightsStore7[0] <= WeightsStore7[476];
			WeightsStore7[1] <= WeightsStore7[477];
			WeightsStore7[2] <= WeightsStore7[478];
			WeightsStore7[3] <= WeightsStore7[479];
			WeightsStore7[4] <= WeightsStore7[480];
			WeightsStore7[5] <= WeightsStore7[481];
			WeightsStore7[6] <= WeightsStore7[482];
			WeightsStore7[7] <= WeightsStore7[483];
			WeightsStore7[8] <= WeightsStore7[484];
			WeightsStore7[9] <= WeightsStore7[485];
			WeightsStore7[10] <= WeightsStore7[486];
			WeightsStore7[11] <= WeightsStore7[487];
			WeightsStore7[12] <= WeightsStore7[488];
			WeightsStore7[13] <= WeightsStore7[489];
			WeightsStore7[14] <= WeightsStore7[490];
			WeightsStore7[15] <= WeightsStore7[491];
			WeightsStore7[16] <= WeightsStore7[492];
			WeightsStore7[17] <= WeightsStore7[493];
			WeightsStore7[18] <= WeightsStore7[494];
			WeightsStore7[19] <= WeightsStore7[495];
			WeightsStore7[20] <= WeightsStore7[496];
			WeightsStore7[21] <= WeightsStore7[497];
			WeightsStore7[22] <= WeightsStore7[498];
			WeightsStore7[23] <= WeightsStore7[499];
			WeightsStore7[24] <= WeightsStore7[500];
			WeightsStore7[25] <= WeightsStore7[501];
			WeightsStore7[26] <= WeightsStore7[502];
			WeightsStore7[27] <= WeightsStore7[503];
			WeightsStore8[0] <= WeightsStore8[476];
			WeightsStore8[1] <= WeightsStore8[477];
			WeightsStore8[2] <= WeightsStore8[478];
			WeightsStore8[3] <= WeightsStore8[479];
			WeightsStore8[4] <= WeightsStore8[480];
			WeightsStore8[5] <= WeightsStore8[481];
			WeightsStore8[6] <= WeightsStore8[482];
			WeightsStore8[7] <= WeightsStore8[483];
			WeightsStore8[8] <= WeightsStore8[484];
			WeightsStore8[9] <= WeightsStore8[485];
			WeightsStore8[10] <= WeightsStore8[486];
			WeightsStore8[11] <= WeightsStore8[487];
			WeightsStore8[12] <= WeightsStore8[488];
			WeightsStore8[13] <= WeightsStore8[489];
			WeightsStore8[14] <= WeightsStore8[490];
			WeightsStore8[15] <= WeightsStore8[491];
			WeightsStore8[16] <= WeightsStore8[492];
			WeightsStore8[17] <= WeightsStore8[493];
			WeightsStore8[18] <= WeightsStore8[494];
			WeightsStore8[19] <= WeightsStore8[495];
			WeightsStore8[20] <= WeightsStore8[496];
			WeightsStore8[21] <= WeightsStore8[497];
			WeightsStore8[22] <= WeightsStore8[498];
			WeightsStore8[23] <= WeightsStore8[499];
			WeightsStore8[24] <= WeightsStore8[500];
			WeightsStore8[25] <= WeightsStore8[501];
			WeightsStore8[26] <= WeightsStore8[502];
			WeightsStore8[27] <= WeightsStore8[503];
			WeightsStore9[0] <= WeightsStore9[476];
			WeightsStore9[1] <= WeightsStore9[477];
			WeightsStore9[2] <= WeightsStore9[478];
			WeightsStore9[3] <= WeightsStore9[479];
			WeightsStore9[4] <= WeightsStore9[480];
			WeightsStore9[5] <= WeightsStore9[481];
			WeightsStore9[6] <= WeightsStore9[482];
			WeightsStore9[7] <= WeightsStore9[483];
			WeightsStore9[8] <= WeightsStore9[484];
			WeightsStore9[9] <= WeightsStore9[485];
			WeightsStore9[10] <= WeightsStore9[486];
			WeightsStore9[11] <= WeightsStore9[487];
			WeightsStore9[12] <= WeightsStore9[488];
			WeightsStore9[13] <= WeightsStore9[489];
			WeightsStore9[14] <= WeightsStore9[490];
			WeightsStore9[15] <= WeightsStore9[491];
			WeightsStore9[16] <= WeightsStore9[492];
			WeightsStore9[17] <= WeightsStore9[493];
			WeightsStore9[18] <= WeightsStore9[494];
			WeightsStore9[19] <= WeightsStore9[495];
			WeightsStore9[20] <= WeightsStore9[496];
			WeightsStore9[21] <= WeightsStore9[497];
			WeightsStore9[22] <= WeightsStore9[498];
			WeightsStore9[23] <= WeightsStore9[499];
			WeightsStore9[24] <= WeightsStore9[500];
			WeightsStore9[25] <= WeightsStore9[501];
			WeightsStore9[26] <= WeightsStore9[502];
			WeightsStore9[27] <= WeightsStore9[503];
		end else if(switchCounter == 32'd125)begin
			PixelsStore[0] <= PixelsStore[504];
			PixelsStore[1] <= PixelsStore[505];
			PixelsStore[2] <= PixelsStore[506];
			PixelsStore[3] <= PixelsStore[507];
			PixelsStore[4] <= PixelsStore[508];
			PixelsStore[5] <= PixelsStore[509];
			PixelsStore[6] <= PixelsStore[510];
			PixelsStore[7] <= PixelsStore[511];
			PixelsStore[8] <= PixelsStore[512];
			PixelsStore[9] <= PixelsStore[513];
			PixelsStore[10] <= PixelsStore[514];
			PixelsStore[11] <= PixelsStore[515];
			PixelsStore[12] <= PixelsStore[516];
			PixelsStore[13] <= PixelsStore[517];
			PixelsStore[14] <= PixelsStore[518];
			PixelsStore[15] <= PixelsStore[519];
			PixelsStore[16] <= PixelsStore[520];
			PixelsStore[17] <= PixelsStore[521];
			PixelsStore[18] <= PixelsStore[522];
			PixelsStore[19] <= PixelsStore[523];
			PixelsStore[20] <= PixelsStore[524];
			PixelsStore[21] <= PixelsStore[525];
			PixelsStore[22] <= PixelsStore[526];
			PixelsStore[23] <= PixelsStore[527];
			PixelsStore[24] <= PixelsStore[528];
			PixelsStore[25] <= PixelsStore[529];
			PixelsStore[26] <= PixelsStore[530];
			PixelsStore[27] <= PixelsStore[531];
			WeightsStore0[0] <= WeightsStore0[504];
			WeightsStore0[1] <= WeightsStore0[505];
			WeightsStore0[2] <= WeightsStore0[506];
			WeightsStore0[3] <= WeightsStore0[507];
			WeightsStore0[4] <= WeightsStore0[508];
			WeightsStore0[5] <= WeightsStore0[509];
			WeightsStore0[6] <= WeightsStore0[510];
			WeightsStore0[7] <= WeightsStore0[511];
			WeightsStore0[8] <= WeightsStore0[512];
			WeightsStore0[9] <= WeightsStore0[513];
			WeightsStore0[10] <= WeightsStore0[514];
			WeightsStore0[11] <= WeightsStore0[515];
			WeightsStore0[12] <= WeightsStore0[516];
			WeightsStore0[13] <= WeightsStore0[517];
			WeightsStore0[14] <= WeightsStore0[518];
			WeightsStore0[15] <= WeightsStore0[519];
			WeightsStore0[16] <= WeightsStore0[520];
			WeightsStore0[17] <= WeightsStore0[521];
			WeightsStore0[18] <= WeightsStore0[522];
			WeightsStore0[19] <= WeightsStore0[523];
			WeightsStore0[20] <= WeightsStore0[524];
			WeightsStore0[21] <= WeightsStore0[525];
			WeightsStore0[22] <= WeightsStore0[526];
			WeightsStore0[23] <= WeightsStore0[527];
			WeightsStore0[24] <= WeightsStore0[528];
			WeightsStore0[25] <= WeightsStore0[529];
			WeightsStore0[26] <= WeightsStore0[530];
			WeightsStore0[27] <= WeightsStore0[531];
			WeightsStore1[0] <= WeightsStore1[504];
			WeightsStore1[1] <= WeightsStore1[505];
			WeightsStore1[2] <= WeightsStore1[506];
			WeightsStore1[3] <= WeightsStore1[507];
			WeightsStore1[4] <= WeightsStore1[508];
			WeightsStore1[5] <= WeightsStore1[509];
			WeightsStore1[6] <= WeightsStore1[510];
			WeightsStore1[7] <= WeightsStore1[511];
			WeightsStore1[8] <= WeightsStore1[512];
			WeightsStore1[9] <= WeightsStore1[513];
			WeightsStore1[10] <= WeightsStore1[514];
			WeightsStore1[11] <= WeightsStore1[515];
			WeightsStore1[12] <= WeightsStore1[516];
			WeightsStore1[13] <= WeightsStore1[517];
			WeightsStore1[14] <= WeightsStore1[518];
			WeightsStore1[15] <= WeightsStore1[519];
			WeightsStore1[16] <= WeightsStore1[520];
			WeightsStore1[17] <= WeightsStore1[521];
			WeightsStore1[18] <= WeightsStore1[522];
			WeightsStore1[19] <= WeightsStore1[523];
			WeightsStore1[20] <= WeightsStore1[524];
			WeightsStore1[21] <= WeightsStore1[525];
			WeightsStore1[22] <= WeightsStore1[526];
			WeightsStore1[23] <= WeightsStore1[527];
			WeightsStore1[24] <= WeightsStore1[528];
			WeightsStore1[25] <= WeightsStore1[529];
			WeightsStore1[26] <= WeightsStore1[530];
			WeightsStore1[27] <= WeightsStore1[531];
			WeightsStore2[0] <= WeightsStore2[504];
			WeightsStore2[1] <= WeightsStore2[505];
			WeightsStore2[2] <= WeightsStore2[506];
			WeightsStore2[3] <= WeightsStore2[507];
			WeightsStore2[4] <= WeightsStore2[508];
			WeightsStore2[5] <= WeightsStore2[509];
			WeightsStore2[6] <= WeightsStore2[510];
			WeightsStore2[7] <= WeightsStore2[511];
			WeightsStore2[8] <= WeightsStore2[512];
			WeightsStore2[9] <= WeightsStore2[513];
			WeightsStore2[10] <= WeightsStore2[514];
			WeightsStore2[11] <= WeightsStore2[515];
			WeightsStore2[12] <= WeightsStore2[516];
			WeightsStore2[13] <= WeightsStore2[517];
			WeightsStore2[14] <= WeightsStore2[518];
			WeightsStore2[15] <= WeightsStore2[519];
			WeightsStore2[16] <= WeightsStore2[520];
			WeightsStore2[17] <= WeightsStore2[521];
			WeightsStore2[18] <= WeightsStore2[522];
			WeightsStore2[19] <= WeightsStore2[523];
			WeightsStore2[20] <= WeightsStore2[524];
			WeightsStore2[21] <= WeightsStore2[525];
			WeightsStore2[22] <= WeightsStore2[526];
			WeightsStore2[23] <= WeightsStore2[527];
			WeightsStore2[24] <= WeightsStore2[528];
			WeightsStore2[25] <= WeightsStore2[529];
			WeightsStore2[26] <= WeightsStore2[530];
			WeightsStore2[27] <= WeightsStore2[531];
			WeightsStore3[0] <= WeightsStore3[504];
			WeightsStore3[1] <= WeightsStore3[505];
			WeightsStore3[2] <= WeightsStore3[506];
			WeightsStore3[3] <= WeightsStore3[507];
			WeightsStore3[4] <= WeightsStore3[508];
			WeightsStore3[5] <= WeightsStore3[509];
			WeightsStore3[6] <= WeightsStore3[510];
			WeightsStore3[7] <= WeightsStore3[511];
			WeightsStore3[8] <= WeightsStore3[512];
			WeightsStore3[9] <= WeightsStore3[513];
			WeightsStore3[10] <= WeightsStore3[514];
			WeightsStore3[11] <= WeightsStore3[515];
			WeightsStore3[12] <= WeightsStore3[516];
			WeightsStore3[13] <= WeightsStore3[517];
			WeightsStore3[14] <= WeightsStore3[518];
			WeightsStore3[15] <= WeightsStore3[519];
			WeightsStore3[16] <= WeightsStore3[520];
			WeightsStore3[17] <= WeightsStore3[521];
			WeightsStore3[18] <= WeightsStore3[522];
			WeightsStore3[19] <= WeightsStore3[523];
			WeightsStore3[20] <= WeightsStore3[524];
			WeightsStore3[21] <= WeightsStore3[525];
			WeightsStore3[22] <= WeightsStore3[526];
			WeightsStore3[23] <= WeightsStore3[527];
			WeightsStore3[24] <= WeightsStore3[528];
			WeightsStore3[25] <= WeightsStore3[529];
			WeightsStore3[26] <= WeightsStore3[530];
			WeightsStore3[27] <= WeightsStore3[531];
			WeightsStore4[0] <= WeightsStore4[504];
			WeightsStore4[1] <= WeightsStore4[505];
			WeightsStore4[2] <= WeightsStore4[506];
			WeightsStore4[3] <= WeightsStore4[507];
			WeightsStore4[4] <= WeightsStore4[508];
			WeightsStore4[5] <= WeightsStore4[509];
			WeightsStore4[6] <= WeightsStore4[510];
			WeightsStore4[7] <= WeightsStore4[511];
			WeightsStore4[8] <= WeightsStore4[512];
			WeightsStore4[9] <= WeightsStore4[513];
			WeightsStore4[10] <= WeightsStore4[514];
			WeightsStore4[11] <= WeightsStore4[515];
			WeightsStore4[12] <= WeightsStore4[516];
			WeightsStore4[13] <= WeightsStore4[517];
			WeightsStore4[14] <= WeightsStore4[518];
			WeightsStore4[15] <= WeightsStore4[519];
			WeightsStore4[16] <= WeightsStore4[520];
			WeightsStore4[17] <= WeightsStore4[521];
			WeightsStore4[18] <= WeightsStore4[522];
			WeightsStore4[19] <= WeightsStore4[523];
			WeightsStore4[20] <= WeightsStore4[524];
			WeightsStore4[21] <= WeightsStore4[525];
			WeightsStore4[22] <= WeightsStore4[526];
			WeightsStore4[23] <= WeightsStore4[527];
			WeightsStore4[24] <= WeightsStore4[528];
			WeightsStore4[25] <= WeightsStore4[529];
			WeightsStore4[26] <= WeightsStore4[530];
			WeightsStore4[27] <= WeightsStore4[531];
			WeightsStore5[0] <= WeightsStore5[504];
			WeightsStore5[1] <= WeightsStore5[505];
			WeightsStore5[2] <= WeightsStore5[506];
			WeightsStore5[3] <= WeightsStore5[507];
			WeightsStore5[4] <= WeightsStore5[508];
			WeightsStore5[5] <= WeightsStore5[509];
			WeightsStore5[6] <= WeightsStore5[510];
			WeightsStore5[7] <= WeightsStore5[511];
			WeightsStore5[8] <= WeightsStore5[512];
			WeightsStore5[9] <= WeightsStore5[513];
			WeightsStore5[10] <= WeightsStore5[514];
			WeightsStore5[11] <= WeightsStore5[515];
			WeightsStore5[12] <= WeightsStore5[516];
			WeightsStore5[13] <= WeightsStore5[517];
			WeightsStore5[14] <= WeightsStore5[518];
			WeightsStore5[15] <= WeightsStore5[519];
			WeightsStore5[16] <= WeightsStore5[520];
			WeightsStore5[17] <= WeightsStore5[521];
			WeightsStore5[18] <= WeightsStore5[522];
			WeightsStore5[19] <= WeightsStore5[523];
			WeightsStore5[20] <= WeightsStore5[524];
			WeightsStore5[21] <= WeightsStore5[525];
			WeightsStore5[22] <= WeightsStore5[526];
			WeightsStore5[23] <= WeightsStore5[527];
			WeightsStore5[24] <= WeightsStore5[528];
			WeightsStore5[25] <= WeightsStore5[529];
			WeightsStore5[26] <= WeightsStore5[530];
			WeightsStore5[27] <= WeightsStore5[531];
			WeightsStore6[0] <= WeightsStore6[504];
			WeightsStore6[1] <= WeightsStore6[505];
			WeightsStore6[2] <= WeightsStore6[506];
			WeightsStore6[3] <= WeightsStore6[507];
			WeightsStore6[4] <= WeightsStore6[508];
			WeightsStore6[5] <= WeightsStore6[509];
			WeightsStore6[6] <= WeightsStore6[510];
			WeightsStore6[7] <= WeightsStore6[511];
			WeightsStore6[8] <= WeightsStore6[512];
			WeightsStore6[9] <= WeightsStore6[513];
			WeightsStore6[10] <= WeightsStore6[514];
			WeightsStore6[11] <= WeightsStore6[515];
			WeightsStore6[12] <= WeightsStore6[516];
			WeightsStore6[13] <= WeightsStore6[517];
			WeightsStore6[14] <= WeightsStore6[518];
			WeightsStore6[15] <= WeightsStore6[519];
			WeightsStore6[16] <= WeightsStore6[520];
			WeightsStore6[17] <= WeightsStore6[521];
			WeightsStore6[18] <= WeightsStore6[522];
			WeightsStore6[19] <= WeightsStore6[523];
			WeightsStore6[20] <= WeightsStore6[524];
			WeightsStore6[21] <= WeightsStore6[525];
			WeightsStore6[22] <= WeightsStore6[526];
			WeightsStore6[23] <= WeightsStore6[527];
			WeightsStore6[24] <= WeightsStore6[528];
			WeightsStore6[25] <= WeightsStore6[529];
			WeightsStore6[26] <= WeightsStore6[530];
			WeightsStore6[27] <= WeightsStore6[531];
			WeightsStore7[0] <= WeightsStore7[504];
			WeightsStore7[1] <= WeightsStore7[505];
			WeightsStore7[2] <= WeightsStore7[506];
			WeightsStore7[3] <= WeightsStore7[507];
			WeightsStore7[4] <= WeightsStore7[508];
			WeightsStore7[5] <= WeightsStore7[509];
			WeightsStore7[6] <= WeightsStore7[510];
			WeightsStore7[7] <= WeightsStore7[511];
			WeightsStore7[8] <= WeightsStore7[512];
			WeightsStore7[9] <= WeightsStore7[513];
			WeightsStore7[10] <= WeightsStore7[514];
			WeightsStore7[11] <= WeightsStore7[515];
			WeightsStore7[12] <= WeightsStore7[516];
			WeightsStore7[13] <= WeightsStore7[517];
			WeightsStore7[14] <= WeightsStore7[518];
			WeightsStore7[15] <= WeightsStore7[519];
			WeightsStore7[16] <= WeightsStore7[520];
			WeightsStore7[17] <= WeightsStore7[521];
			WeightsStore7[18] <= WeightsStore7[522];
			WeightsStore7[19] <= WeightsStore7[523];
			WeightsStore7[20] <= WeightsStore7[524];
			WeightsStore7[21] <= WeightsStore7[525];
			WeightsStore7[22] <= WeightsStore7[526];
			WeightsStore7[23] <= WeightsStore7[527];
			WeightsStore7[24] <= WeightsStore7[528];
			WeightsStore7[25] <= WeightsStore7[529];
			WeightsStore7[26] <= WeightsStore7[530];
			WeightsStore7[27] <= WeightsStore7[531];
			WeightsStore8[0] <= WeightsStore8[504];
			WeightsStore8[1] <= WeightsStore8[505];
			WeightsStore8[2] <= WeightsStore8[506];
			WeightsStore8[3] <= WeightsStore8[507];
			WeightsStore8[4] <= WeightsStore8[508];
			WeightsStore8[5] <= WeightsStore8[509];
			WeightsStore8[6] <= WeightsStore8[510];
			WeightsStore8[7] <= WeightsStore8[511];
			WeightsStore8[8] <= WeightsStore8[512];
			WeightsStore8[9] <= WeightsStore8[513];
			WeightsStore8[10] <= WeightsStore8[514];
			WeightsStore8[11] <= WeightsStore8[515];
			WeightsStore8[12] <= WeightsStore8[516];
			WeightsStore8[13] <= WeightsStore8[517];
			WeightsStore8[14] <= WeightsStore8[518];
			WeightsStore8[15] <= WeightsStore8[519];
			WeightsStore8[16] <= WeightsStore8[520];
			WeightsStore8[17] <= WeightsStore8[521];
			WeightsStore8[18] <= WeightsStore8[522];
			WeightsStore8[19] <= WeightsStore8[523];
			WeightsStore8[20] <= WeightsStore8[524];
			WeightsStore8[21] <= WeightsStore8[525];
			WeightsStore8[22] <= WeightsStore8[526];
			WeightsStore8[23] <= WeightsStore8[527];
			WeightsStore8[24] <= WeightsStore8[528];
			WeightsStore8[25] <= WeightsStore8[529];
			WeightsStore8[26] <= WeightsStore8[530];
			WeightsStore8[27] <= WeightsStore8[531];
			WeightsStore9[0] <= WeightsStore9[504];
			WeightsStore9[1] <= WeightsStore9[505];
			WeightsStore9[2] <= WeightsStore9[506];
			WeightsStore9[3] <= WeightsStore9[507];
			WeightsStore9[4] <= WeightsStore9[508];
			WeightsStore9[5] <= WeightsStore9[509];
			WeightsStore9[6] <= WeightsStore9[510];
			WeightsStore9[7] <= WeightsStore9[511];
			WeightsStore9[8] <= WeightsStore9[512];
			WeightsStore9[9] <= WeightsStore9[513];
			WeightsStore9[10] <= WeightsStore9[514];
			WeightsStore9[11] <= WeightsStore9[515];
			WeightsStore9[12] <= WeightsStore9[516];
			WeightsStore9[13] <= WeightsStore9[517];
			WeightsStore9[14] <= WeightsStore9[518];
			WeightsStore9[15] <= WeightsStore9[519];
			WeightsStore9[16] <= WeightsStore9[520];
			WeightsStore9[17] <= WeightsStore9[521];
			WeightsStore9[18] <= WeightsStore9[522];
			WeightsStore9[19] <= WeightsStore9[523];
			WeightsStore9[20] <= WeightsStore9[524];
			WeightsStore9[21] <= WeightsStore9[525];
			WeightsStore9[22] <= WeightsStore9[526];
			WeightsStore9[23] <= WeightsStore9[527];
			WeightsStore9[24] <= WeightsStore9[528];
			WeightsStore9[25] <= WeightsStore9[529];
			WeightsStore9[26] <= WeightsStore9[530];
			WeightsStore9[27] <= WeightsStore9[531];
		end else if(switchCounter == 32'd132)begin
			PixelsStore[0] <= PixelsStore[532];
			PixelsStore[1] <= PixelsStore[533];
			PixelsStore[2] <= PixelsStore[534];
			PixelsStore[3] <= PixelsStore[535];
			PixelsStore[4] <= PixelsStore[536];
			PixelsStore[5] <= PixelsStore[537];
			PixelsStore[6] <= PixelsStore[538];
			PixelsStore[7] <= PixelsStore[539];
			PixelsStore[8] <= PixelsStore[540];
			PixelsStore[9] <= PixelsStore[541];
			PixelsStore[10] <= PixelsStore[542];
			PixelsStore[11] <= PixelsStore[543];
			PixelsStore[12] <= PixelsStore[544];
			PixelsStore[13] <= PixelsStore[545];
			PixelsStore[14] <= PixelsStore[546];
			PixelsStore[15] <= PixelsStore[547];
			PixelsStore[16] <= PixelsStore[548];
			PixelsStore[17] <= PixelsStore[549];
			PixelsStore[18] <= PixelsStore[550];
			PixelsStore[19] <= PixelsStore[551];
			PixelsStore[20] <= PixelsStore[552];
			PixelsStore[21] <= PixelsStore[553];
			PixelsStore[22] <= PixelsStore[554];
			PixelsStore[23] <= PixelsStore[555];
			PixelsStore[24] <= PixelsStore[556];
			PixelsStore[25] <= PixelsStore[557];
			PixelsStore[26] <= PixelsStore[558];
			PixelsStore[27] <= PixelsStore[559];
			WeightsStore0[0] <= WeightsStore0[532];
			WeightsStore0[1] <= WeightsStore0[533];
			WeightsStore0[2] <= WeightsStore0[534];
			WeightsStore0[3] <= WeightsStore0[535];
			WeightsStore0[4] <= WeightsStore0[536];
			WeightsStore0[5] <= WeightsStore0[537];
			WeightsStore0[6] <= WeightsStore0[538];
			WeightsStore0[7] <= WeightsStore0[539];
			WeightsStore0[8] <= WeightsStore0[540];
			WeightsStore0[9] <= WeightsStore0[541];
			WeightsStore0[10] <= WeightsStore0[542];
			WeightsStore0[11] <= WeightsStore0[543];
			WeightsStore0[12] <= WeightsStore0[544];
			WeightsStore0[13] <= WeightsStore0[545];
			WeightsStore0[14] <= WeightsStore0[546];
			WeightsStore0[15] <= WeightsStore0[547];
			WeightsStore0[16] <= WeightsStore0[548];
			WeightsStore0[17] <= WeightsStore0[549];
			WeightsStore0[18] <= WeightsStore0[550];
			WeightsStore0[19] <= WeightsStore0[551];
			WeightsStore0[20] <= WeightsStore0[552];
			WeightsStore0[21] <= WeightsStore0[553];
			WeightsStore0[22] <= WeightsStore0[554];
			WeightsStore0[23] <= WeightsStore0[555];
			WeightsStore0[24] <= WeightsStore0[556];
			WeightsStore0[25] <= WeightsStore0[557];
			WeightsStore0[26] <= WeightsStore0[558];
			WeightsStore0[27] <= WeightsStore0[559];
			WeightsStore1[0] <= WeightsStore1[532];
			WeightsStore1[1] <= WeightsStore1[533];
			WeightsStore1[2] <= WeightsStore1[534];
			WeightsStore1[3] <= WeightsStore1[535];
			WeightsStore1[4] <= WeightsStore1[536];
			WeightsStore1[5] <= WeightsStore1[537];
			WeightsStore1[6] <= WeightsStore1[538];
			WeightsStore1[7] <= WeightsStore1[539];
			WeightsStore1[8] <= WeightsStore1[540];
			WeightsStore1[9] <= WeightsStore1[541];
			WeightsStore1[10] <= WeightsStore1[542];
			WeightsStore1[11] <= WeightsStore1[543];
			WeightsStore1[12] <= WeightsStore1[544];
			WeightsStore1[13] <= WeightsStore1[545];
			WeightsStore1[14] <= WeightsStore1[546];
			WeightsStore1[15] <= WeightsStore1[547];
			WeightsStore1[16] <= WeightsStore1[548];
			WeightsStore1[17] <= WeightsStore1[549];
			WeightsStore1[18] <= WeightsStore1[550];
			WeightsStore1[19] <= WeightsStore1[551];
			WeightsStore1[20] <= WeightsStore1[552];
			WeightsStore1[21] <= WeightsStore1[553];
			WeightsStore1[22] <= WeightsStore1[554];
			WeightsStore1[23] <= WeightsStore1[555];
			WeightsStore1[24] <= WeightsStore1[556];
			WeightsStore1[25] <= WeightsStore1[557];
			WeightsStore1[26] <= WeightsStore1[558];
			WeightsStore1[27] <= WeightsStore1[559];
			WeightsStore2[0] <= WeightsStore2[532];
			WeightsStore2[1] <= WeightsStore2[533];
			WeightsStore2[2] <= WeightsStore2[534];
			WeightsStore2[3] <= WeightsStore2[535];
			WeightsStore2[4] <= WeightsStore2[536];
			WeightsStore2[5] <= WeightsStore2[537];
			WeightsStore2[6] <= WeightsStore2[538];
			WeightsStore2[7] <= WeightsStore2[539];
			WeightsStore2[8] <= WeightsStore2[540];
			WeightsStore2[9] <= WeightsStore2[541];
			WeightsStore2[10] <= WeightsStore2[542];
			WeightsStore2[11] <= WeightsStore2[543];
			WeightsStore2[12] <= WeightsStore2[544];
			WeightsStore2[13] <= WeightsStore2[545];
			WeightsStore2[14] <= WeightsStore2[546];
			WeightsStore2[15] <= WeightsStore2[547];
			WeightsStore2[16] <= WeightsStore2[548];
			WeightsStore2[17] <= WeightsStore2[549];
			WeightsStore2[18] <= WeightsStore2[550];
			WeightsStore2[19] <= WeightsStore2[551];
			WeightsStore2[20] <= WeightsStore2[552];
			WeightsStore2[21] <= WeightsStore2[553];
			WeightsStore2[22] <= WeightsStore2[554];
			WeightsStore2[23] <= WeightsStore2[555];
			WeightsStore2[24] <= WeightsStore2[556];
			WeightsStore2[25] <= WeightsStore2[557];
			WeightsStore2[26] <= WeightsStore2[558];
			WeightsStore2[27] <= WeightsStore2[559];
			WeightsStore3[0] <= WeightsStore3[532];
			WeightsStore3[1] <= WeightsStore3[533];
			WeightsStore3[2] <= WeightsStore3[534];
			WeightsStore3[3] <= WeightsStore3[535];
			WeightsStore3[4] <= WeightsStore3[536];
			WeightsStore3[5] <= WeightsStore3[537];
			WeightsStore3[6] <= WeightsStore3[538];
			WeightsStore3[7] <= WeightsStore3[539];
			WeightsStore3[8] <= WeightsStore3[540];
			WeightsStore3[9] <= WeightsStore3[541];
			WeightsStore3[10] <= WeightsStore3[542];
			WeightsStore3[11] <= WeightsStore3[543];
			WeightsStore3[12] <= WeightsStore3[544];
			WeightsStore3[13] <= WeightsStore3[545];
			WeightsStore3[14] <= WeightsStore3[546];
			WeightsStore3[15] <= WeightsStore3[547];
			WeightsStore3[16] <= WeightsStore3[548];
			WeightsStore3[17] <= WeightsStore3[549];
			WeightsStore3[18] <= WeightsStore3[550];
			WeightsStore3[19] <= WeightsStore3[551];
			WeightsStore3[20] <= WeightsStore3[552];
			WeightsStore3[21] <= WeightsStore3[553];
			WeightsStore3[22] <= WeightsStore3[554];
			WeightsStore3[23] <= WeightsStore3[555];
			WeightsStore3[24] <= WeightsStore3[556];
			WeightsStore3[25] <= WeightsStore3[557];
			WeightsStore3[26] <= WeightsStore3[558];
			WeightsStore3[27] <= WeightsStore3[559];
			WeightsStore4[0] <= WeightsStore4[532];
			WeightsStore4[1] <= WeightsStore4[533];
			WeightsStore4[2] <= WeightsStore4[534];
			WeightsStore4[3] <= WeightsStore4[535];
			WeightsStore4[4] <= WeightsStore4[536];
			WeightsStore4[5] <= WeightsStore4[537];
			WeightsStore4[6] <= WeightsStore4[538];
			WeightsStore4[7] <= WeightsStore4[539];
			WeightsStore4[8] <= WeightsStore4[540];
			WeightsStore4[9] <= WeightsStore4[541];
			WeightsStore4[10] <= WeightsStore4[542];
			WeightsStore4[11] <= WeightsStore4[543];
			WeightsStore4[12] <= WeightsStore4[544];
			WeightsStore4[13] <= WeightsStore4[545];
			WeightsStore4[14] <= WeightsStore4[546];
			WeightsStore4[15] <= WeightsStore4[547];
			WeightsStore4[16] <= WeightsStore4[548];
			WeightsStore4[17] <= WeightsStore4[549];
			WeightsStore4[18] <= WeightsStore4[550];
			WeightsStore4[19] <= WeightsStore4[551];
			WeightsStore4[20] <= WeightsStore4[552];
			WeightsStore4[21] <= WeightsStore4[553];
			WeightsStore4[22] <= WeightsStore4[554];
			WeightsStore4[23] <= WeightsStore4[555];
			WeightsStore4[24] <= WeightsStore4[556];
			WeightsStore4[25] <= WeightsStore4[557];
			WeightsStore4[26] <= WeightsStore4[558];
			WeightsStore4[27] <= WeightsStore4[559];
			WeightsStore5[0] <= WeightsStore5[532];
			WeightsStore5[1] <= WeightsStore5[533];
			WeightsStore5[2] <= WeightsStore5[534];
			WeightsStore5[3] <= WeightsStore5[535];
			WeightsStore5[4] <= WeightsStore5[536];
			WeightsStore5[5] <= WeightsStore5[537];
			WeightsStore5[6] <= WeightsStore5[538];
			WeightsStore5[7] <= WeightsStore5[539];
			WeightsStore5[8] <= WeightsStore5[540];
			WeightsStore5[9] <= WeightsStore5[541];
			WeightsStore5[10] <= WeightsStore5[542];
			WeightsStore5[11] <= WeightsStore5[543];
			WeightsStore5[12] <= WeightsStore5[544];
			WeightsStore5[13] <= WeightsStore5[545];
			WeightsStore5[14] <= WeightsStore5[546];
			WeightsStore5[15] <= WeightsStore5[547];
			WeightsStore5[16] <= WeightsStore5[548];
			WeightsStore5[17] <= WeightsStore5[549];
			WeightsStore5[18] <= WeightsStore5[550];
			WeightsStore5[19] <= WeightsStore5[551];
			WeightsStore5[20] <= WeightsStore5[552];
			WeightsStore5[21] <= WeightsStore5[553];
			WeightsStore5[22] <= WeightsStore5[554];
			WeightsStore5[23] <= WeightsStore5[555];
			WeightsStore5[24] <= WeightsStore5[556];
			WeightsStore5[25] <= WeightsStore5[557];
			WeightsStore5[26] <= WeightsStore5[558];
			WeightsStore5[27] <= WeightsStore5[559];
			WeightsStore6[0] <= WeightsStore6[532];
			WeightsStore6[1] <= WeightsStore6[533];
			WeightsStore6[2] <= WeightsStore6[534];
			WeightsStore6[3] <= WeightsStore6[535];
			WeightsStore6[4] <= WeightsStore6[536];
			WeightsStore6[5] <= WeightsStore6[537];
			WeightsStore6[6] <= WeightsStore6[538];
			WeightsStore6[7] <= WeightsStore6[539];
			WeightsStore6[8] <= WeightsStore6[540];
			WeightsStore6[9] <= WeightsStore6[541];
			WeightsStore6[10] <= WeightsStore6[542];
			WeightsStore6[11] <= WeightsStore6[543];
			WeightsStore6[12] <= WeightsStore6[544];
			WeightsStore6[13] <= WeightsStore6[545];
			WeightsStore6[14] <= WeightsStore6[546];
			WeightsStore6[15] <= WeightsStore6[547];
			WeightsStore6[16] <= WeightsStore6[548];
			WeightsStore6[17] <= WeightsStore6[549];
			WeightsStore6[18] <= WeightsStore6[550];
			WeightsStore6[19] <= WeightsStore6[551];
			WeightsStore6[20] <= WeightsStore6[552];
			WeightsStore6[21] <= WeightsStore6[553];
			WeightsStore6[22] <= WeightsStore6[554];
			WeightsStore6[23] <= WeightsStore6[555];
			WeightsStore6[24] <= WeightsStore6[556];
			WeightsStore6[25] <= WeightsStore6[557];
			WeightsStore6[26] <= WeightsStore6[558];
			WeightsStore6[27] <= WeightsStore6[559];
			WeightsStore7[0] <= WeightsStore7[532];
			WeightsStore7[1] <= WeightsStore7[533];
			WeightsStore7[2] <= WeightsStore7[534];
			WeightsStore7[3] <= WeightsStore7[535];
			WeightsStore7[4] <= WeightsStore7[536];
			WeightsStore7[5] <= WeightsStore7[537];
			WeightsStore7[6] <= WeightsStore7[538];
			WeightsStore7[7] <= WeightsStore7[539];
			WeightsStore7[8] <= WeightsStore7[540];
			WeightsStore7[9] <= WeightsStore7[541];
			WeightsStore7[10] <= WeightsStore7[542];
			WeightsStore7[11] <= WeightsStore7[543];
			WeightsStore7[12] <= WeightsStore7[544];
			WeightsStore7[13] <= WeightsStore7[545];
			WeightsStore7[14] <= WeightsStore7[546];
			WeightsStore7[15] <= WeightsStore7[547];
			WeightsStore7[16] <= WeightsStore7[548];
			WeightsStore7[17] <= WeightsStore7[549];
			WeightsStore7[18] <= WeightsStore7[550];
			WeightsStore7[19] <= WeightsStore7[551];
			WeightsStore7[20] <= WeightsStore7[552];
			WeightsStore7[21] <= WeightsStore7[553];
			WeightsStore7[22] <= WeightsStore7[554];
			WeightsStore7[23] <= WeightsStore7[555];
			WeightsStore7[24] <= WeightsStore7[556];
			WeightsStore7[25] <= WeightsStore7[557];
			WeightsStore7[26] <= WeightsStore7[558];
			WeightsStore7[27] <= WeightsStore7[559];
			WeightsStore8[0] <= WeightsStore8[532];
			WeightsStore8[1] <= WeightsStore8[533];
			WeightsStore8[2] <= WeightsStore8[534];
			WeightsStore8[3] <= WeightsStore8[535];
			WeightsStore8[4] <= WeightsStore8[536];
			WeightsStore8[5] <= WeightsStore8[537];
			WeightsStore8[6] <= WeightsStore8[538];
			WeightsStore8[7] <= WeightsStore8[539];
			WeightsStore8[8] <= WeightsStore8[540];
			WeightsStore8[9] <= WeightsStore8[541];
			WeightsStore8[10] <= WeightsStore8[542];
			WeightsStore8[11] <= WeightsStore8[543];
			WeightsStore8[12] <= WeightsStore8[544];
			WeightsStore8[13] <= WeightsStore8[545];
			WeightsStore8[14] <= WeightsStore8[546];
			WeightsStore8[15] <= WeightsStore8[547];
			WeightsStore8[16] <= WeightsStore8[548];
			WeightsStore8[17] <= WeightsStore8[549];
			WeightsStore8[18] <= WeightsStore8[550];
			WeightsStore8[19] <= WeightsStore8[551];
			WeightsStore8[20] <= WeightsStore8[552];
			WeightsStore8[21] <= WeightsStore8[553];
			WeightsStore8[22] <= WeightsStore8[554];
			WeightsStore8[23] <= WeightsStore8[555];
			WeightsStore8[24] <= WeightsStore8[556];
			WeightsStore8[25] <= WeightsStore8[557];
			WeightsStore8[26] <= WeightsStore8[558];
			WeightsStore8[27] <= WeightsStore8[559];
			WeightsStore9[0] <= WeightsStore9[532];
			WeightsStore9[1] <= WeightsStore9[533];
			WeightsStore9[2] <= WeightsStore9[534];
			WeightsStore9[3] <= WeightsStore9[535];
			WeightsStore9[4] <= WeightsStore9[536];
			WeightsStore9[5] <= WeightsStore9[537];
			WeightsStore9[6] <= WeightsStore9[538];
			WeightsStore9[7] <= WeightsStore9[539];
			WeightsStore9[8] <= WeightsStore9[540];
			WeightsStore9[9] <= WeightsStore9[541];
			WeightsStore9[10] <= WeightsStore9[542];
			WeightsStore9[11] <= WeightsStore9[543];
			WeightsStore9[12] <= WeightsStore9[544];
			WeightsStore9[13] <= WeightsStore9[545];
			WeightsStore9[14] <= WeightsStore9[546];
			WeightsStore9[15] <= WeightsStore9[547];
			WeightsStore9[16] <= WeightsStore9[548];
			WeightsStore9[17] <= WeightsStore9[549];
			WeightsStore9[18] <= WeightsStore9[550];
			WeightsStore9[19] <= WeightsStore9[551];
			WeightsStore9[20] <= WeightsStore9[552];
			WeightsStore9[21] <= WeightsStore9[553];
			WeightsStore9[22] <= WeightsStore9[554];
			WeightsStore9[23] <= WeightsStore9[555];
			WeightsStore9[24] <= WeightsStore9[556];
			WeightsStore9[25] <= WeightsStore9[557];
			WeightsStore9[26] <= WeightsStore9[558];
			WeightsStore9[27] <= WeightsStore9[559];
		end else if(switchCounter == 32'd139)begin
			PixelsStore[0] <= PixelsStore[560];
			PixelsStore[1] <= PixelsStore[561];
			PixelsStore[2] <= PixelsStore[562];
			PixelsStore[3] <= PixelsStore[563];
			PixelsStore[4] <= PixelsStore[564];
			PixelsStore[5] <= PixelsStore[565];
			PixelsStore[6] <= PixelsStore[566];
			PixelsStore[7] <= PixelsStore[567];
			PixelsStore[8] <= PixelsStore[568];
			PixelsStore[9] <= PixelsStore[569];
			PixelsStore[10] <= PixelsStore[570];
			PixelsStore[11] <= PixelsStore[571];
			PixelsStore[12] <= PixelsStore[572];
			PixelsStore[13] <= PixelsStore[573];
			PixelsStore[14] <= PixelsStore[574];
			PixelsStore[15] <= PixelsStore[575];
			PixelsStore[16] <= PixelsStore[576];
			PixelsStore[17] <= PixelsStore[577];
			PixelsStore[18] <= PixelsStore[578];
			PixelsStore[19] <= PixelsStore[579];
			PixelsStore[20] <= PixelsStore[580];
			PixelsStore[21] <= PixelsStore[581];
			PixelsStore[22] <= PixelsStore[582];
			PixelsStore[23] <= PixelsStore[583];
			PixelsStore[24] <= PixelsStore[584];
			PixelsStore[25] <= PixelsStore[585];
			PixelsStore[26] <= PixelsStore[586];
			PixelsStore[27] <= PixelsStore[587];
			WeightsStore0[0] <= WeightsStore0[560];
			WeightsStore0[1] <= WeightsStore0[561];
			WeightsStore0[2] <= WeightsStore0[562];
			WeightsStore0[3] <= WeightsStore0[563];
			WeightsStore0[4] <= WeightsStore0[564];
			WeightsStore0[5] <= WeightsStore0[565];
			WeightsStore0[6] <= WeightsStore0[566];
			WeightsStore0[7] <= WeightsStore0[567];
			WeightsStore0[8] <= WeightsStore0[568];
			WeightsStore0[9] <= WeightsStore0[569];
			WeightsStore0[10] <= WeightsStore0[570];
			WeightsStore0[11] <= WeightsStore0[571];
			WeightsStore0[12] <= WeightsStore0[572];
			WeightsStore0[13] <= WeightsStore0[573];
			WeightsStore0[14] <= WeightsStore0[574];
			WeightsStore0[15] <= WeightsStore0[575];
			WeightsStore0[16] <= WeightsStore0[576];
			WeightsStore0[17] <= WeightsStore0[577];
			WeightsStore0[18] <= WeightsStore0[578];
			WeightsStore0[19] <= WeightsStore0[579];
			WeightsStore0[20] <= WeightsStore0[580];
			WeightsStore0[21] <= WeightsStore0[581];
			WeightsStore0[22] <= WeightsStore0[582];
			WeightsStore0[23] <= WeightsStore0[583];
			WeightsStore0[24] <= WeightsStore0[584];
			WeightsStore0[25] <= WeightsStore0[585];
			WeightsStore0[26] <= WeightsStore0[586];
			WeightsStore0[27] <= WeightsStore0[587];
			WeightsStore1[0] <= WeightsStore1[560];
			WeightsStore1[1] <= WeightsStore1[561];
			WeightsStore1[2] <= WeightsStore1[562];
			WeightsStore1[3] <= WeightsStore1[563];
			WeightsStore1[4] <= WeightsStore1[564];
			WeightsStore1[5] <= WeightsStore1[565];
			WeightsStore1[6] <= WeightsStore1[566];
			WeightsStore1[7] <= WeightsStore1[567];
			WeightsStore1[8] <= WeightsStore1[568];
			WeightsStore1[9] <= WeightsStore1[569];
			WeightsStore1[10] <= WeightsStore1[570];
			WeightsStore1[11] <= WeightsStore1[571];
			WeightsStore1[12] <= WeightsStore1[572];
			WeightsStore1[13] <= WeightsStore1[573];
			WeightsStore1[14] <= WeightsStore1[574];
			WeightsStore1[15] <= WeightsStore1[575];
			WeightsStore1[16] <= WeightsStore1[576];
			WeightsStore1[17] <= WeightsStore1[577];
			WeightsStore1[18] <= WeightsStore1[578];
			WeightsStore1[19] <= WeightsStore1[579];
			WeightsStore1[20] <= WeightsStore1[580];
			WeightsStore1[21] <= WeightsStore1[581];
			WeightsStore1[22] <= WeightsStore1[582];
			WeightsStore1[23] <= WeightsStore1[583];
			WeightsStore1[24] <= WeightsStore1[584];
			WeightsStore1[25] <= WeightsStore1[585];
			WeightsStore1[26] <= WeightsStore1[586];
			WeightsStore1[27] <= WeightsStore1[587];
			WeightsStore2[0] <= WeightsStore2[560];
			WeightsStore2[1] <= WeightsStore2[561];
			WeightsStore2[2] <= WeightsStore2[562];
			WeightsStore2[3] <= WeightsStore2[563];
			WeightsStore2[4] <= WeightsStore2[564];
			WeightsStore2[5] <= WeightsStore2[565];
			WeightsStore2[6] <= WeightsStore2[566];
			WeightsStore2[7] <= WeightsStore2[567];
			WeightsStore2[8] <= WeightsStore2[568];
			WeightsStore2[9] <= WeightsStore2[569];
			WeightsStore2[10] <= WeightsStore2[570];
			WeightsStore2[11] <= WeightsStore2[571];
			WeightsStore2[12] <= WeightsStore2[572];
			WeightsStore2[13] <= WeightsStore2[573];
			WeightsStore2[14] <= WeightsStore2[574];
			WeightsStore2[15] <= WeightsStore2[575];
			WeightsStore2[16] <= WeightsStore2[576];
			WeightsStore2[17] <= WeightsStore2[577];
			WeightsStore2[18] <= WeightsStore2[578];
			WeightsStore2[19] <= WeightsStore2[579];
			WeightsStore2[20] <= WeightsStore2[580];
			WeightsStore2[21] <= WeightsStore2[581];
			WeightsStore2[22] <= WeightsStore2[582];
			WeightsStore2[23] <= WeightsStore2[583];
			WeightsStore2[24] <= WeightsStore2[584];
			WeightsStore2[25] <= WeightsStore2[585];
			WeightsStore2[26] <= WeightsStore2[586];
			WeightsStore2[27] <= WeightsStore2[587];
			WeightsStore3[0] <= WeightsStore3[560];
			WeightsStore3[1] <= WeightsStore3[561];
			WeightsStore3[2] <= WeightsStore3[562];
			WeightsStore3[3] <= WeightsStore3[563];
			WeightsStore3[4] <= WeightsStore3[564];
			WeightsStore3[5] <= WeightsStore3[565];
			WeightsStore3[6] <= WeightsStore3[566];
			WeightsStore3[7] <= WeightsStore3[567];
			WeightsStore3[8] <= WeightsStore3[568];
			WeightsStore3[9] <= WeightsStore3[569];
			WeightsStore3[10] <= WeightsStore3[570];
			WeightsStore3[11] <= WeightsStore3[571];
			WeightsStore3[12] <= WeightsStore3[572];
			WeightsStore3[13] <= WeightsStore3[573];
			WeightsStore3[14] <= WeightsStore3[574];
			WeightsStore3[15] <= WeightsStore3[575];
			WeightsStore3[16] <= WeightsStore3[576];
			WeightsStore3[17] <= WeightsStore3[577];
			WeightsStore3[18] <= WeightsStore3[578];
			WeightsStore3[19] <= WeightsStore3[579];
			WeightsStore3[20] <= WeightsStore3[580];
			WeightsStore3[21] <= WeightsStore3[581];
			WeightsStore3[22] <= WeightsStore3[582];
			WeightsStore3[23] <= WeightsStore3[583];
			WeightsStore3[24] <= WeightsStore3[584];
			WeightsStore3[25] <= WeightsStore3[585];
			WeightsStore3[26] <= WeightsStore3[586];
			WeightsStore3[27] <= WeightsStore3[587];
			WeightsStore4[0] <= WeightsStore4[560];
			WeightsStore4[1] <= WeightsStore4[561];
			WeightsStore4[2] <= WeightsStore4[562];
			WeightsStore4[3] <= WeightsStore4[563];
			WeightsStore4[4] <= WeightsStore4[564];
			WeightsStore4[5] <= WeightsStore4[565];
			WeightsStore4[6] <= WeightsStore4[566];
			WeightsStore4[7] <= WeightsStore4[567];
			WeightsStore4[8] <= WeightsStore4[568];
			WeightsStore4[9] <= WeightsStore4[569];
			WeightsStore4[10] <= WeightsStore4[570];
			WeightsStore4[11] <= WeightsStore4[571];
			WeightsStore4[12] <= WeightsStore4[572];
			WeightsStore4[13] <= WeightsStore4[573];
			WeightsStore4[14] <= WeightsStore4[574];
			WeightsStore4[15] <= WeightsStore4[575];
			WeightsStore4[16] <= WeightsStore4[576];
			WeightsStore4[17] <= WeightsStore4[577];
			WeightsStore4[18] <= WeightsStore4[578];
			WeightsStore4[19] <= WeightsStore4[579];
			WeightsStore4[20] <= WeightsStore4[580];
			WeightsStore4[21] <= WeightsStore4[581];
			WeightsStore4[22] <= WeightsStore4[582];
			WeightsStore4[23] <= WeightsStore4[583];
			WeightsStore4[24] <= WeightsStore4[584];
			WeightsStore4[25] <= WeightsStore4[585];
			WeightsStore4[26] <= WeightsStore4[586];
			WeightsStore4[27] <= WeightsStore4[587];
			WeightsStore5[0] <= WeightsStore5[560];
			WeightsStore5[1] <= WeightsStore5[561];
			WeightsStore5[2] <= WeightsStore5[562];
			WeightsStore5[3] <= WeightsStore5[563];
			WeightsStore5[4] <= WeightsStore5[564];
			WeightsStore5[5] <= WeightsStore5[565];
			WeightsStore5[6] <= WeightsStore5[566];
			WeightsStore5[7] <= WeightsStore5[567];
			WeightsStore5[8] <= WeightsStore5[568];
			WeightsStore5[9] <= WeightsStore5[569];
			WeightsStore5[10] <= WeightsStore5[570];
			WeightsStore5[11] <= WeightsStore5[571];
			WeightsStore5[12] <= WeightsStore5[572];
			WeightsStore5[13] <= WeightsStore5[573];
			WeightsStore5[14] <= WeightsStore5[574];
			WeightsStore5[15] <= WeightsStore5[575];
			WeightsStore5[16] <= WeightsStore5[576];
			WeightsStore5[17] <= WeightsStore5[577];
			WeightsStore5[18] <= WeightsStore5[578];
			WeightsStore5[19] <= WeightsStore5[579];
			WeightsStore5[20] <= WeightsStore5[580];
			WeightsStore5[21] <= WeightsStore5[581];
			WeightsStore5[22] <= WeightsStore5[582];
			WeightsStore5[23] <= WeightsStore5[583];
			WeightsStore5[24] <= WeightsStore5[584];
			WeightsStore5[25] <= WeightsStore5[585];
			WeightsStore5[26] <= WeightsStore5[586];
			WeightsStore5[27] <= WeightsStore5[587];
			WeightsStore6[0] <= WeightsStore6[560];
			WeightsStore6[1] <= WeightsStore6[561];
			WeightsStore6[2] <= WeightsStore6[562];
			WeightsStore6[3] <= WeightsStore6[563];
			WeightsStore6[4] <= WeightsStore6[564];
			WeightsStore6[5] <= WeightsStore6[565];
			WeightsStore6[6] <= WeightsStore6[566];
			WeightsStore6[7] <= WeightsStore6[567];
			WeightsStore6[8] <= WeightsStore6[568];
			WeightsStore6[9] <= WeightsStore6[569];
			WeightsStore6[10] <= WeightsStore6[570];
			WeightsStore6[11] <= WeightsStore6[571];
			WeightsStore6[12] <= WeightsStore6[572];
			WeightsStore6[13] <= WeightsStore6[573];
			WeightsStore6[14] <= WeightsStore6[574];
			WeightsStore6[15] <= WeightsStore6[575];
			WeightsStore6[16] <= WeightsStore6[576];
			WeightsStore6[17] <= WeightsStore6[577];
			WeightsStore6[18] <= WeightsStore6[578];
			WeightsStore6[19] <= WeightsStore6[579];
			WeightsStore6[20] <= WeightsStore6[580];
			WeightsStore6[21] <= WeightsStore6[581];
			WeightsStore6[22] <= WeightsStore6[582];
			WeightsStore6[23] <= WeightsStore6[583];
			WeightsStore6[24] <= WeightsStore6[584];
			WeightsStore6[25] <= WeightsStore6[585];
			WeightsStore6[26] <= WeightsStore6[586];
			WeightsStore6[27] <= WeightsStore6[587];
			WeightsStore7[0] <= WeightsStore7[560];
			WeightsStore7[1] <= WeightsStore7[561];
			WeightsStore7[2] <= WeightsStore7[562];
			WeightsStore7[3] <= WeightsStore7[563];
			WeightsStore7[4] <= WeightsStore7[564];
			WeightsStore7[5] <= WeightsStore7[565];
			WeightsStore7[6] <= WeightsStore7[566];
			WeightsStore7[7] <= WeightsStore7[567];
			WeightsStore7[8] <= WeightsStore7[568];
			WeightsStore7[9] <= WeightsStore7[569];
			WeightsStore7[10] <= WeightsStore7[570];
			WeightsStore7[11] <= WeightsStore7[571];
			WeightsStore7[12] <= WeightsStore7[572];
			WeightsStore7[13] <= WeightsStore7[573];
			WeightsStore7[14] <= WeightsStore7[574];
			WeightsStore7[15] <= WeightsStore7[575];
			WeightsStore7[16] <= WeightsStore7[576];
			WeightsStore7[17] <= WeightsStore7[577];
			WeightsStore7[18] <= WeightsStore7[578];
			WeightsStore7[19] <= WeightsStore7[579];
			WeightsStore7[20] <= WeightsStore7[580];
			WeightsStore7[21] <= WeightsStore7[581];
			WeightsStore7[22] <= WeightsStore7[582];
			WeightsStore7[23] <= WeightsStore7[583];
			WeightsStore7[24] <= WeightsStore7[584];
			WeightsStore7[25] <= WeightsStore7[585];
			WeightsStore7[26] <= WeightsStore7[586];
			WeightsStore7[27] <= WeightsStore7[587];
			WeightsStore8[0] <= WeightsStore8[560];
			WeightsStore8[1] <= WeightsStore8[561];
			WeightsStore8[2] <= WeightsStore8[562];
			WeightsStore8[3] <= WeightsStore8[563];
			WeightsStore8[4] <= WeightsStore8[564];
			WeightsStore8[5] <= WeightsStore8[565];
			WeightsStore8[6] <= WeightsStore8[566];
			WeightsStore8[7] <= WeightsStore8[567];
			WeightsStore8[8] <= WeightsStore8[568];
			WeightsStore8[9] <= WeightsStore8[569];
			WeightsStore8[10] <= WeightsStore8[570];
			WeightsStore8[11] <= WeightsStore8[571];
			WeightsStore8[12] <= WeightsStore8[572];
			WeightsStore8[13] <= WeightsStore8[573];
			WeightsStore8[14] <= WeightsStore8[574];
			WeightsStore8[15] <= WeightsStore8[575];
			WeightsStore8[16] <= WeightsStore8[576];
			WeightsStore8[17] <= WeightsStore8[577];
			WeightsStore8[18] <= WeightsStore8[578];
			WeightsStore8[19] <= WeightsStore8[579];
			WeightsStore8[20] <= WeightsStore8[580];
			WeightsStore8[21] <= WeightsStore8[581];
			WeightsStore8[22] <= WeightsStore8[582];
			WeightsStore8[23] <= WeightsStore8[583];
			WeightsStore8[24] <= WeightsStore8[584];
			WeightsStore8[25] <= WeightsStore8[585];
			WeightsStore8[26] <= WeightsStore8[586];
			WeightsStore8[27] <= WeightsStore8[587];
			WeightsStore9[0] <= WeightsStore9[560];
			WeightsStore9[1] <= WeightsStore9[561];
			WeightsStore9[2] <= WeightsStore9[562];
			WeightsStore9[3] <= WeightsStore9[563];
			WeightsStore9[4] <= WeightsStore9[564];
			WeightsStore9[5] <= WeightsStore9[565];
			WeightsStore9[6] <= WeightsStore9[566];
			WeightsStore9[7] <= WeightsStore9[567];
			WeightsStore9[8] <= WeightsStore9[568];
			WeightsStore9[9] <= WeightsStore9[569];
			WeightsStore9[10] <= WeightsStore9[570];
			WeightsStore9[11] <= WeightsStore9[571];
			WeightsStore9[12] <= WeightsStore9[572];
			WeightsStore9[13] <= WeightsStore9[573];
			WeightsStore9[14] <= WeightsStore9[574];
			WeightsStore9[15] <= WeightsStore9[575];
			WeightsStore9[16] <= WeightsStore9[576];
			WeightsStore9[17] <= WeightsStore9[577];
			WeightsStore9[18] <= WeightsStore9[578];
			WeightsStore9[19] <= WeightsStore9[579];
			WeightsStore9[20] <= WeightsStore9[580];
			WeightsStore9[21] <= WeightsStore9[581];
			WeightsStore9[22] <= WeightsStore9[582];
			WeightsStore9[23] <= WeightsStore9[583];
			WeightsStore9[24] <= WeightsStore9[584];
			WeightsStore9[25] <= WeightsStore9[585];
			WeightsStore9[26] <= WeightsStore9[586];
			WeightsStore9[27] <= WeightsStore9[587];
		end else if(switchCounter == 32'd146)begin
			PixelsStore[0] <= PixelsStore[588];
			PixelsStore[1] <= PixelsStore[589];
			PixelsStore[2] <= PixelsStore[590];
			PixelsStore[3] <= PixelsStore[591];
			PixelsStore[4] <= PixelsStore[592];
			PixelsStore[5] <= PixelsStore[593];
			PixelsStore[6] <= PixelsStore[594];
			PixelsStore[7] <= PixelsStore[595];
			PixelsStore[8] <= PixelsStore[596];
			PixelsStore[9] <= PixelsStore[597];
			PixelsStore[10] <= PixelsStore[598];
			PixelsStore[11] <= PixelsStore[599];
			PixelsStore[12] <= PixelsStore[600];
			PixelsStore[13] <= PixelsStore[601];
			PixelsStore[14] <= PixelsStore[602];
			PixelsStore[15] <= PixelsStore[603];
			PixelsStore[16] <= PixelsStore[604];
			PixelsStore[17] <= PixelsStore[605];
			PixelsStore[18] <= PixelsStore[606];
			PixelsStore[19] <= PixelsStore[607];
			PixelsStore[20] <= PixelsStore[608];
			PixelsStore[21] <= PixelsStore[609];
			PixelsStore[22] <= PixelsStore[610];
			PixelsStore[23] <= PixelsStore[611];
			PixelsStore[24] <= PixelsStore[612];
			PixelsStore[25] <= PixelsStore[613];
			PixelsStore[26] <= PixelsStore[614];
			PixelsStore[27] <= PixelsStore[615];
			WeightsStore0[0] <= WeightsStore0[588];
			WeightsStore0[1] <= WeightsStore0[589];
			WeightsStore0[2] <= WeightsStore0[590];
			WeightsStore0[3] <= WeightsStore0[591];
			WeightsStore0[4] <= WeightsStore0[592];
			WeightsStore0[5] <= WeightsStore0[593];
			WeightsStore0[6] <= WeightsStore0[594];
			WeightsStore0[7] <= WeightsStore0[595];
			WeightsStore0[8] <= WeightsStore0[596];
			WeightsStore0[9] <= WeightsStore0[597];
			WeightsStore0[10] <= WeightsStore0[598];
			WeightsStore0[11] <= WeightsStore0[599];
			WeightsStore0[12] <= WeightsStore0[600];
			WeightsStore0[13] <= WeightsStore0[601];
			WeightsStore0[14] <= WeightsStore0[602];
			WeightsStore0[15] <= WeightsStore0[603];
			WeightsStore0[16] <= WeightsStore0[604];
			WeightsStore0[17] <= WeightsStore0[605];
			WeightsStore0[18] <= WeightsStore0[606];
			WeightsStore0[19] <= WeightsStore0[607];
			WeightsStore0[20] <= WeightsStore0[608];
			WeightsStore0[21] <= WeightsStore0[609];
			WeightsStore0[22] <= WeightsStore0[610];
			WeightsStore0[23] <= WeightsStore0[611];
			WeightsStore0[24] <= WeightsStore0[612];
			WeightsStore0[25] <= WeightsStore0[613];
			WeightsStore0[26] <= WeightsStore0[614];
			WeightsStore0[27] <= WeightsStore0[615];
			WeightsStore1[0] <= WeightsStore1[588];
			WeightsStore1[1] <= WeightsStore1[589];
			WeightsStore1[2] <= WeightsStore1[590];
			WeightsStore1[3] <= WeightsStore1[591];
			WeightsStore1[4] <= WeightsStore1[592];
			WeightsStore1[5] <= WeightsStore1[593];
			WeightsStore1[6] <= WeightsStore1[594];
			WeightsStore1[7] <= WeightsStore1[595];
			WeightsStore1[8] <= WeightsStore1[596];
			WeightsStore1[9] <= WeightsStore1[597];
			WeightsStore1[10] <= WeightsStore1[598];
			WeightsStore1[11] <= WeightsStore1[599];
			WeightsStore1[12] <= WeightsStore1[600];
			WeightsStore1[13] <= WeightsStore1[601];
			WeightsStore1[14] <= WeightsStore1[602];
			WeightsStore1[15] <= WeightsStore1[603];
			WeightsStore1[16] <= WeightsStore1[604];
			WeightsStore1[17] <= WeightsStore1[605];
			WeightsStore1[18] <= WeightsStore1[606];
			WeightsStore1[19] <= WeightsStore1[607];
			WeightsStore1[20] <= WeightsStore1[608];
			WeightsStore1[21] <= WeightsStore1[609];
			WeightsStore1[22] <= WeightsStore1[610];
			WeightsStore1[23] <= WeightsStore1[611];
			WeightsStore1[24] <= WeightsStore1[612];
			WeightsStore1[25] <= WeightsStore1[613];
			WeightsStore1[26] <= WeightsStore1[614];
			WeightsStore1[27] <= WeightsStore1[615];
			WeightsStore2[0] <= WeightsStore2[588];
			WeightsStore2[1] <= WeightsStore2[589];
			WeightsStore2[2] <= WeightsStore2[590];
			WeightsStore2[3] <= WeightsStore2[591];
			WeightsStore2[4] <= WeightsStore2[592];
			WeightsStore2[5] <= WeightsStore2[593];
			WeightsStore2[6] <= WeightsStore2[594];
			WeightsStore2[7] <= WeightsStore2[595];
			WeightsStore2[8] <= WeightsStore2[596];
			WeightsStore2[9] <= WeightsStore2[597];
			WeightsStore2[10] <= WeightsStore2[598];
			WeightsStore2[11] <= WeightsStore2[599];
			WeightsStore2[12] <= WeightsStore2[600];
			WeightsStore2[13] <= WeightsStore2[601];
			WeightsStore2[14] <= WeightsStore2[602];
			WeightsStore2[15] <= WeightsStore2[603];
			WeightsStore2[16] <= WeightsStore2[604];
			WeightsStore2[17] <= WeightsStore2[605];
			WeightsStore2[18] <= WeightsStore2[606];
			WeightsStore2[19] <= WeightsStore2[607];
			WeightsStore2[20] <= WeightsStore2[608];
			WeightsStore2[21] <= WeightsStore2[609];
			WeightsStore2[22] <= WeightsStore2[610];
			WeightsStore2[23] <= WeightsStore2[611];
			WeightsStore2[24] <= WeightsStore2[612];
			WeightsStore2[25] <= WeightsStore2[613];
			WeightsStore2[26] <= WeightsStore2[614];
			WeightsStore2[27] <= WeightsStore2[615];
			WeightsStore3[0] <= WeightsStore3[588];
			WeightsStore3[1] <= WeightsStore3[589];
			WeightsStore3[2] <= WeightsStore3[590];
			WeightsStore3[3] <= WeightsStore3[591];
			WeightsStore3[4] <= WeightsStore3[592];
			WeightsStore3[5] <= WeightsStore3[593];
			WeightsStore3[6] <= WeightsStore3[594];
			WeightsStore3[7] <= WeightsStore3[595];
			WeightsStore3[8] <= WeightsStore3[596];
			WeightsStore3[9] <= WeightsStore3[597];
			WeightsStore3[10] <= WeightsStore3[598];
			WeightsStore3[11] <= WeightsStore3[599];
			WeightsStore3[12] <= WeightsStore3[600];
			WeightsStore3[13] <= WeightsStore3[601];
			WeightsStore3[14] <= WeightsStore3[602];
			WeightsStore3[15] <= WeightsStore3[603];
			WeightsStore3[16] <= WeightsStore3[604];
			WeightsStore3[17] <= WeightsStore3[605];
			WeightsStore3[18] <= WeightsStore3[606];
			WeightsStore3[19] <= WeightsStore3[607];
			WeightsStore3[20] <= WeightsStore3[608];
			WeightsStore3[21] <= WeightsStore3[609];
			WeightsStore3[22] <= WeightsStore3[610];
			WeightsStore3[23] <= WeightsStore3[611];
			WeightsStore3[24] <= WeightsStore3[612];
			WeightsStore3[25] <= WeightsStore3[613];
			WeightsStore3[26] <= WeightsStore3[614];
			WeightsStore3[27] <= WeightsStore3[615];
			WeightsStore4[0] <= WeightsStore4[588];
			WeightsStore4[1] <= WeightsStore4[589];
			WeightsStore4[2] <= WeightsStore4[590];
			WeightsStore4[3] <= WeightsStore4[591];
			WeightsStore4[4] <= WeightsStore4[592];
			WeightsStore4[5] <= WeightsStore4[593];
			WeightsStore4[6] <= WeightsStore4[594];
			WeightsStore4[7] <= WeightsStore4[595];
			WeightsStore4[8] <= WeightsStore4[596];
			WeightsStore4[9] <= WeightsStore4[597];
			WeightsStore4[10] <= WeightsStore4[598];
			WeightsStore4[11] <= WeightsStore4[599];
			WeightsStore4[12] <= WeightsStore4[600];
			WeightsStore4[13] <= WeightsStore4[601];
			WeightsStore4[14] <= WeightsStore4[602];
			WeightsStore4[15] <= WeightsStore4[603];
			WeightsStore4[16] <= WeightsStore4[604];
			WeightsStore4[17] <= WeightsStore4[605];
			WeightsStore4[18] <= WeightsStore4[606];
			WeightsStore4[19] <= WeightsStore4[607];
			WeightsStore4[20] <= WeightsStore4[608];
			WeightsStore4[21] <= WeightsStore4[609];
			WeightsStore4[22] <= WeightsStore4[610];
			WeightsStore4[23] <= WeightsStore4[611];
			WeightsStore4[24] <= WeightsStore4[612];
			WeightsStore4[25] <= WeightsStore4[613];
			WeightsStore4[26] <= WeightsStore4[614];
			WeightsStore4[27] <= WeightsStore4[615];
			WeightsStore5[0] <= WeightsStore5[588];
			WeightsStore5[1] <= WeightsStore5[589];
			WeightsStore5[2] <= WeightsStore5[590];
			WeightsStore5[3] <= WeightsStore5[591];
			WeightsStore5[4] <= WeightsStore5[592];
			WeightsStore5[5] <= WeightsStore5[593];
			WeightsStore5[6] <= WeightsStore5[594];
			WeightsStore5[7] <= WeightsStore5[595];
			WeightsStore5[8] <= WeightsStore5[596];
			WeightsStore5[9] <= WeightsStore5[597];
			WeightsStore5[10] <= WeightsStore5[598];
			WeightsStore5[11] <= WeightsStore5[599];
			WeightsStore5[12] <= WeightsStore5[600];
			WeightsStore5[13] <= WeightsStore5[601];
			WeightsStore5[14] <= WeightsStore5[602];
			WeightsStore5[15] <= WeightsStore5[603];
			WeightsStore5[16] <= WeightsStore5[604];
			WeightsStore5[17] <= WeightsStore5[605];
			WeightsStore5[18] <= WeightsStore5[606];
			WeightsStore5[19] <= WeightsStore5[607];
			WeightsStore5[20] <= WeightsStore5[608];
			WeightsStore5[21] <= WeightsStore5[609];
			WeightsStore5[22] <= WeightsStore5[610];
			WeightsStore5[23] <= WeightsStore5[611];
			WeightsStore5[24] <= WeightsStore5[612];
			WeightsStore5[25] <= WeightsStore5[613];
			WeightsStore5[26] <= WeightsStore5[614];
			WeightsStore5[27] <= WeightsStore5[615];
			WeightsStore6[0] <= WeightsStore6[588];
			WeightsStore6[1] <= WeightsStore6[589];
			WeightsStore6[2] <= WeightsStore6[590];
			WeightsStore6[3] <= WeightsStore6[591];
			WeightsStore6[4] <= WeightsStore6[592];
			WeightsStore6[5] <= WeightsStore6[593];
			WeightsStore6[6] <= WeightsStore6[594];
			WeightsStore6[7] <= WeightsStore6[595];
			WeightsStore6[8] <= WeightsStore6[596];
			WeightsStore6[9] <= WeightsStore6[597];
			WeightsStore6[10] <= WeightsStore6[598];
			WeightsStore6[11] <= WeightsStore6[599];
			WeightsStore6[12] <= WeightsStore6[600];
			WeightsStore6[13] <= WeightsStore6[601];
			WeightsStore6[14] <= WeightsStore6[602];
			WeightsStore6[15] <= WeightsStore6[603];
			WeightsStore6[16] <= WeightsStore6[604];
			WeightsStore6[17] <= WeightsStore6[605];
			WeightsStore6[18] <= WeightsStore6[606];
			WeightsStore6[19] <= WeightsStore6[607];
			WeightsStore6[20] <= WeightsStore6[608];
			WeightsStore6[21] <= WeightsStore6[609];
			WeightsStore6[22] <= WeightsStore6[610];
			WeightsStore6[23] <= WeightsStore6[611];
			WeightsStore6[24] <= WeightsStore6[612];
			WeightsStore6[25] <= WeightsStore6[613];
			WeightsStore6[26] <= WeightsStore6[614];
			WeightsStore6[27] <= WeightsStore6[615];
			WeightsStore7[0] <= WeightsStore7[588];
			WeightsStore7[1] <= WeightsStore7[589];
			WeightsStore7[2] <= WeightsStore7[590];
			WeightsStore7[3] <= WeightsStore7[591];
			WeightsStore7[4] <= WeightsStore7[592];
			WeightsStore7[5] <= WeightsStore7[593];
			WeightsStore7[6] <= WeightsStore7[594];
			WeightsStore7[7] <= WeightsStore7[595];
			WeightsStore7[8] <= WeightsStore7[596];
			WeightsStore7[9] <= WeightsStore7[597];
			WeightsStore7[10] <= WeightsStore7[598];
			WeightsStore7[11] <= WeightsStore7[599];
			WeightsStore7[12] <= WeightsStore7[600];
			WeightsStore7[13] <= WeightsStore7[601];
			WeightsStore7[14] <= WeightsStore7[602];
			WeightsStore7[15] <= WeightsStore7[603];
			WeightsStore7[16] <= WeightsStore7[604];
			WeightsStore7[17] <= WeightsStore7[605];
			WeightsStore7[18] <= WeightsStore7[606];
			WeightsStore7[19] <= WeightsStore7[607];
			WeightsStore7[20] <= WeightsStore7[608];
			WeightsStore7[21] <= WeightsStore7[609];
			WeightsStore7[22] <= WeightsStore7[610];
			WeightsStore7[23] <= WeightsStore7[611];
			WeightsStore7[24] <= WeightsStore7[612];
			WeightsStore7[25] <= WeightsStore7[613];
			WeightsStore7[26] <= WeightsStore7[614];
			WeightsStore7[27] <= WeightsStore7[615];
			WeightsStore8[0] <= WeightsStore8[588];
			WeightsStore8[1] <= WeightsStore8[589];
			WeightsStore8[2] <= WeightsStore8[590];
			WeightsStore8[3] <= WeightsStore8[591];
			WeightsStore8[4] <= WeightsStore8[592];
			WeightsStore8[5] <= WeightsStore8[593];
			WeightsStore8[6] <= WeightsStore8[594];
			WeightsStore8[7] <= WeightsStore8[595];
			WeightsStore8[8] <= WeightsStore8[596];
			WeightsStore8[9] <= WeightsStore8[597];
			WeightsStore8[10] <= WeightsStore8[598];
			WeightsStore8[11] <= WeightsStore8[599];
			WeightsStore8[12] <= WeightsStore8[600];
			WeightsStore8[13] <= WeightsStore8[601];
			WeightsStore8[14] <= WeightsStore8[602];
			WeightsStore8[15] <= WeightsStore8[603];
			WeightsStore8[16] <= WeightsStore8[604];
			WeightsStore8[17] <= WeightsStore8[605];
			WeightsStore8[18] <= WeightsStore8[606];
			WeightsStore8[19] <= WeightsStore8[607];
			WeightsStore8[20] <= WeightsStore8[608];
			WeightsStore8[21] <= WeightsStore8[609];
			WeightsStore8[22] <= WeightsStore8[610];
			WeightsStore8[23] <= WeightsStore8[611];
			WeightsStore8[24] <= WeightsStore8[612];
			WeightsStore8[25] <= WeightsStore8[613];
			WeightsStore8[26] <= WeightsStore8[614];
			WeightsStore8[27] <= WeightsStore8[615];
			WeightsStore9[0] <= WeightsStore9[588];
			WeightsStore9[1] <= WeightsStore9[589];
			WeightsStore9[2] <= WeightsStore9[590];
			WeightsStore9[3] <= WeightsStore9[591];
			WeightsStore9[4] <= WeightsStore9[592];
			WeightsStore9[5] <= WeightsStore9[593];
			WeightsStore9[6] <= WeightsStore9[594];
			WeightsStore9[7] <= WeightsStore9[595];
			WeightsStore9[8] <= WeightsStore9[596];
			WeightsStore9[9] <= WeightsStore9[597];
			WeightsStore9[10] <= WeightsStore9[598];
			WeightsStore9[11] <= WeightsStore9[599];
			WeightsStore9[12] <= WeightsStore9[600];
			WeightsStore9[13] <= WeightsStore9[601];
			WeightsStore9[14] <= WeightsStore9[602];
			WeightsStore9[15] <= WeightsStore9[603];
			WeightsStore9[16] <= WeightsStore9[604];
			WeightsStore9[17] <= WeightsStore9[605];
			WeightsStore9[18] <= WeightsStore9[606];
			WeightsStore9[19] <= WeightsStore9[607];
			WeightsStore9[20] <= WeightsStore9[608];
			WeightsStore9[21] <= WeightsStore9[609];
			WeightsStore9[22] <= WeightsStore9[610];
			WeightsStore9[23] <= WeightsStore9[611];
			WeightsStore9[24] <= WeightsStore9[612];
			WeightsStore9[25] <= WeightsStore9[613];
			WeightsStore9[26] <= WeightsStore9[614];
			WeightsStore9[27] <= WeightsStore9[615];
		end else if(switchCounter == 32'd153)begin
			PixelsStore[0] <= PixelsStore[616];
			PixelsStore[1] <= PixelsStore[617];
			PixelsStore[2] <= PixelsStore[618];
			PixelsStore[3] <= PixelsStore[619];
			PixelsStore[4] <= PixelsStore[620];
			PixelsStore[5] <= PixelsStore[621];
			PixelsStore[6] <= PixelsStore[622];
			PixelsStore[7] <= PixelsStore[623];
			PixelsStore[8] <= PixelsStore[624];
			PixelsStore[9] <= PixelsStore[625];
			PixelsStore[10] <= PixelsStore[626];
			PixelsStore[11] <= PixelsStore[627];
			PixelsStore[12] <= PixelsStore[628];
			PixelsStore[13] <= PixelsStore[629];
			PixelsStore[14] <= PixelsStore[630];
			PixelsStore[15] <= PixelsStore[631];
			PixelsStore[16] <= PixelsStore[632];
			PixelsStore[17] <= PixelsStore[633];
			PixelsStore[18] <= PixelsStore[634];
			PixelsStore[19] <= PixelsStore[635];
			PixelsStore[20] <= PixelsStore[636];
			PixelsStore[21] <= PixelsStore[637];
			PixelsStore[22] <= PixelsStore[638];
			PixelsStore[23] <= PixelsStore[639];
			PixelsStore[24] <= PixelsStore[640];
			PixelsStore[25] <= PixelsStore[641];
			PixelsStore[26] <= PixelsStore[642];
			PixelsStore[27] <= PixelsStore[643];
			WeightsStore0[0] <= WeightsStore0[616];
			WeightsStore0[1] <= WeightsStore0[617];
			WeightsStore0[2] <= WeightsStore0[618];
			WeightsStore0[3] <= WeightsStore0[619];
			WeightsStore0[4] <= WeightsStore0[620];
			WeightsStore0[5] <= WeightsStore0[621];
			WeightsStore0[6] <= WeightsStore0[622];
			WeightsStore0[7] <= WeightsStore0[623];
			WeightsStore0[8] <= WeightsStore0[624];
			WeightsStore0[9] <= WeightsStore0[625];
			WeightsStore0[10] <= WeightsStore0[626];
			WeightsStore0[11] <= WeightsStore0[627];
			WeightsStore0[12] <= WeightsStore0[628];
			WeightsStore0[13] <= WeightsStore0[629];
			WeightsStore0[14] <= WeightsStore0[630];
			WeightsStore0[15] <= WeightsStore0[631];
			WeightsStore0[16] <= WeightsStore0[632];
			WeightsStore0[17] <= WeightsStore0[633];
			WeightsStore0[18] <= WeightsStore0[634];
			WeightsStore0[19] <= WeightsStore0[635];
			WeightsStore0[20] <= WeightsStore0[636];
			WeightsStore0[21] <= WeightsStore0[637];
			WeightsStore0[22] <= WeightsStore0[638];
			WeightsStore0[23] <= WeightsStore0[639];
			WeightsStore0[24] <= WeightsStore0[640];
			WeightsStore0[25] <= WeightsStore0[641];
			WeightsStore0[26] <= WeightsStore0[642];
			WeightsStore0[27] <= WeightsStore0[643];
			WeightsStore1[0] <= WeightsStore1[616];
			WeightsStore1[1] <= WeightsStore1[617];
			WeightsStore1[2] <= WeightsStore1[618];
			WeightsStore1[3] <= WeightsStore1[619];
			WeightsStore1[4] <= WeightsStore1[620];
			WeightsStore1[5] <= WeightsStore1[621];
			WeightsStore1[6] <= WeightsStore1[622];
			WeightsStore1[7] <= WeightsStore1[623];
			WeightsStore1[8] <= WeightsStore1[624];
			WeightsStore1[9] <= WeightsStore1[625];
			WeightsStore1[10] <= WeightsStore1[626];
			WeightsStore1[11] <= WeightsStore1[627];
			WeightsStore1[12] <= WeightsStore1[628];
			WeightsStore1[13] <= WeightsStore1[629];
			WeightsStore1[14] <= WeightsStore1[630];
			WeightsStore1[15] <= WeightsStore1[631];
			WeightsStore1[16] <= WeightsStore1[632];
			WeightsStore1[17] <= WeightsStore1[633];
			WeightsStore1[18] <= WeightsStore1[634];
			WeightsStore1[19] <= WeightsStore1[635];
			WeightsStore1[20] <= WeightsStore1[636];
			WeightsStore1[21] <= WeightsStore1[637];
			WeightsStore1[22] <= WeightsStore1[638];
			WeightsStore1[23] <= WeightsStore1[639];
			WeightsStore1[24] <= WeightsStore1[640];
			WeightsStore1[25] <= WeightsStore1[641];
			WeightsStore1[26] <= WeightsStore1[642];
			WeightsStore1[27] <= WeightsStore1[643];
			WeightsStore2[0] <= WeightsStore2[616];
			WeightsStore2[1] <= WeightsStore2[617];
			WeightsStore2[2] <= WeightsStore2[618];
			WeightsStore2[3] <= WeightsStore2[619];
			WeightsStore2[4] <= WeightsStore2[620];
			WeightsStore2[5] <= WeightsStore2[621];
			WeightsStore2[6] <= WeightsStore2[622];
			WeightsStore2[7] <= WeightsStore2[623];
			WeightsStore2[8] <= WeightsStore2[624];
			WeightsStore2[9] <= WeightsStore2[625];
			WeightsStore2[10] <= WeightsStore2[626];
			WeightsStore2[11] <= WeightsStore2[627];
			WeightsStore2[12] <= WeightsStore2[628];
			WeightsStore2[13] <= WeightsStore2[629];
			WeightsStore2[14] <= WeightsStore2[630];
			WeightsStore2[15] <= WeightsStore2[631];
			WeightsStore2[16] <= WeightsStore2[632];
			WeightsStore2[17] <= WeightsStore2[633];
			WeightsStore2[18] <= WeightsStore2[634];
			WeightsStore2[19] <= WeightsStore2[635];
			WeightsStore2[20] <= WeightsStore2[636];
			WeightsStore2[21] <= WeightsStore2[637];
			WeightsStore2[22] <= WeightsStore2[638];
			WeightsStore2[23] <= WeightsStore2[639];
			WeightsStore2[24] <= WeightsStore2[640];
			WeightsStore2[25] <= WeightsStore2[641];
			WeightsStore2[26] <= WeightsStore2[642];
			WeightsStore2[27] <= WeightsStore2[643];
			WeightsStore3[0] <= WeightsStore3[616];
			WeightsStore3[1] <= WeightsStore3[617];
			WeightsStore3[2] <= WeightsStore3[618];
			WeightsStore3[3] <= WeightsStore3[619];
			WeightsStore3[4] <= WeightsStore3[620];
			WeightsStore3[5] <= WeightsStore3[621];
			WeightsStore3[6] <= WeightsStore3[622];
			WeightsStore3[7] <= WeightsStore3[623];
			WeightsStore3[8] <= WeightsStore3[624];
			WeightsStore3[9] <= WeightsStore3[625];
			WeightsStore3[10] <= WeightsStore3[626];
			WeightsStore3[11] <= WeightsStore3[627];
			WeightsStore3[12] <= WeightsStore3[628];
			WeightsStore3[13] <= WeightsStore3[629];
			WeightsStore3[14] <= WeightsStore3[630];
			WeightsStore3[15] <= WeightsStore3[631];
			WeightsStore3[16] <= WeightsStore3[632];
			WeightsStore3[17] <= WeightsStore3[633];
			WeightsStore3[18] <= WeightsStore3[634];
			WeightsStore3[19] <= WeightsStore3[635];
			WeightsStore3[20] <= WeightsStore3[636];
			WeightsStore3[21] <= WeightsStore3[637];
			WeightsStore3[22] <= WeightsStore3[638];
			WeightsStore3[23] <= WeightsStore3[639];
			WeightsStore3[24] <= WeightsStore3[640];
			WeightsStore3[25] <= WeightsStore3[641];
			WeightsStore3[26] <= WeightsStore3[642];
			WeightsStore3[27] <= WeightsStore3[643];
			WeightsStore4[0] <= WeightsStore4[616];
			WeightsStore4[1] <= WeightsStore4[617];
			WeightsStore4[2] <= WeightsStore4[618];
			WeightsStore4[3] <= WeightsStore4[619];
			WeightsStore4[4] <= WeightsStore4[620];
			WeightsStore4[5] <= WeightsStore4[621];
			WeightsStore4[6] <= WeightsStore4[622];
			WeightsStore4[7] <= WeightsStore4[623];
			WeightsStore4[8] <= WeightsStore4[624];
			WeightsStore4[9] <= WeightsStore4[625];
			WeightsStore4[10] <= WeightsStore4[626];
			WeightsStore4[11] <= WeightsStore4[627];
			WeightsStore4[12] <= WeightsStore4[628];
			WeightsStore4[13] <= WeightsStore4[629];
			WeightsStore4[14] <= WeightsStore4[630];
			WeightsStore4[15] <= WeightsStore4[631];
			WeightsStore4[16] <= WeightsStore4[632];
			WeightsStore4[17] <= WeightsStore4[633];
			WeightsStore4[18] <= WeightsStore4[634];
			WeightsStore4[19] <= WeightsStore4[635];
			WeightsStore4[20] <= WeightsStore4[636];
			WeightsStore4[21] <= WeightsStore4[637];
			WeightsStore4[22] <= WeightsStore4[638];
			WeightsStore4[23] <= WeightsStore4[639];
			WeightsStore4[24] <= WeightsStore4[640];
			WeightsStore4[25] <= WeightsStore4[641];
			WeightsStore4[26] <= WeightsStore4[642];
			WeightsStore4[27] <= WeightsStore4[643];
			WeightsStore5[0] <= WeightsStore5[616];
			WeightsStore5[1] <= WeightsStore5[617];
			WeightsStore5[2] <= WeightsStore5[618];
			WeightsStore5[3] <= WeightsStore5[619];
			WeightsStore5[4] <= WeightsStore5[620];
			WeightsStore5[5] <= WeightsStore5[621];
			WeightsStore5[6] <= WeightsStore5[622];
			WeightsStore5[7] <= WeightsStore5[623];
			WeightsStore5[8] <= WeightsStore5[624];
			WeightsStore5[9] <= WeightsStore5[625];
			WeightsStore5[10] <= WeightsStore5[626];
			WeightsStore5[11] <= WeightsStore5[627];
			WeightsStore5[12] <= WeightsStore5[628];
			WeightsStore5[13] <= WeightsStore5[629];
			WeightsStore5[14] <= WeightsStore5[630];
			WeightsStore5[15] <= WeightsStore5[631];
			WeightsStore5[16] <= WeightsStore5[632];
			WeightsStore5[17] <= WeightsStore5[633];
			WeightsStore5[18] <= WeightsStore5[634];
			WeightsStore5[19] <= WeightsStore5[635];
			WeightsStore5[20] <= WeightsStore5[636];
			WeightsStore5[21] <= WeightsStore5[637];
			WeightsStore5[22] <= WeightsStore5[638];
			WeightsStore5[23] <= WeightsStore5[639];
			WeightsStore5[24] <= WeightsStore5[640];
			WeightsStore5[25] <= WeightsStore5[641];
			WeightsStore5[26] <= WeightsStore5[642];
			WeightsStore5[27] <= WeightsStore5[643];
			WeightsStore6[0] <= WeightsStore6[616];
			WeightsStore6[1] <= WeightsStore6[617];
			WeightsStore6[2] <= WeightsStore6[618];
			WeightsStore6[3] <= WeightsStore6[619];
			WeightsStore6[4] <= WeightsStore6[620];
			WeightsStore6[5] <= WeightsStore6[621];
			WeightsStore6[6] <= WeightsStore6[622];
			WeightsStore6[7] <= WeightsStore6[623];
			WeightsStore6[8] <= WeightsStore6[624];
			WeightsStore6[9] <= WeightsStore6[625];
			WeightsStore6[10] <= WeightsStore6[626];
			WeightsStore6[11] <= WeightsStore6[627];
			WeightsStore6[12] <= WeightsStore6[628];
			WeightsStore6[13] <= WeightsStore6[629];
			WeightsStore6[14] <= WeightsStore6[630];
			WeightsStore6[15] <= WeightsStore6[631];
			WeightsStore6[16] <= WeightsStore6[632];
			WeightsStore6[17] <= WeightsStore6[633];
			WeightsStore6[18] <= WeightsStore6[634];
			WeightsStore6[19] <= WeightsStore6[635];
			WeightsStore6[20] <= WeightsStore6[636];
			WeightsStore6[21] <= WeightsStore6[637];
			WeightsStore6[22] <= WeightsStore6[638];
			WeightsStore6[23] <= WeightsStore6[639];
			WeightsStore6[24] <= WeightsStore6[640];
			WeightsStore6[25] <= WeightsStore6[641];
			WeightsStore6[26] <= WeightsStore6[642];
			WeightsStore6[27] <= WeightsStore6[643];
			WeightsStore7[0] <= WeightsStore7[616];
			WeightsStore7[1] <= WeightsStore7[617];
			WeightsStore7[2] <= WeightsStore7[618];
			WeightsStore7[3] <= WeightsStore7[619];
			WeightsStore7[4] <= WeightsStore7[620];
			WeightsStore7[5] <= WeightsStore7[621];
			WeightsStore7[6] <= WeightsStore7[622];
			WeightsStore7[7] <= WeightsStore7[623];
			WeightsStore7[8] <= WeightsStore7[624];
			WeightsStore7[9] <= WeightsStore7[625];
			WeightsStore7[10] <= WeightsStore7[626];
			WeightsStore7[11] <= WeightsStore7[627];
			WeightsStore7[12] <= WeightsStore7[628];
			WeightsStore7[13] <= WeightsStore7[629];
			WeightsStore7[14] <= WeightsStore7[630];
			WeightsStore7[15] <= WeightsStore7[631];
			WeightsStore7[16] <= WeightsStore7[632];
			WeightsStore7[17] <= WeightsStore7[633];
			WeightsStore7[18] <= WeightsStore7[634];
			WeightsStore7[19] <= WeightsStore7[635];
			WeightsStore7[20] <= WeightsStore7[636];
			WeightsStore7[21] <= WeightsStore7[637];
			WeightsStore7[22] <= WeightsStore7[638];
			WeightsStore7[23] <= WeightsStore7[639];
			WeightsStore7[24] <= WeightsStore7[640];
			WeightsStore7[25] <= WeightsStore7[641];
			WeightsStore7[26] <= WeightsStore7[642];
			WeightsStore7[27] <= WeightsStore7[643];
			WeightsStore8[0] <= WeightsStore8[616];
			WeightsStore8[1] <= WeightsStore8[617];
			WeightsStore8[2] <= WeightsStore8[618];
			WeightsStore8[3] <= WeightsStore8[619];
			WeightsStore8[4] <= WeightsStore8[620];
			WeightsStore8[5] <= WeightsStore8[621];
			WeightsStore8[6] <= WeightsStore8[622];
			WeightsStore8[7] <= WeightsStore8[623];
			WeightsStore8[8] <= WeightsStore8[624];
			WeightsStore8[9] <= WeightsStore8[625];
			WeightsStore8[10] <= WeightsStore8[626];
			WeightsStore8[11] <= WeightsStore8[627];
			WeightsStore8[12] <= WeightsStore8[628];
			WeightsStore8[13] <= WeightsStore8[629];
			WeightsStore8[14] <= WeightsStore8[630];
			WeightsStore8[15] <= WeightsStore8[631];
			WeightsStore8[16] <= WeightsStore8[632];
			WeightsStore8[17] <= WeightsStore8[633];
			WeightsStore8[18] <= WeightsStore8[634];
			WeightsStore8[19] <= WeightsStore8[635];
			WeightsStore8[20] <= WeightsStore8[636];
			WeightsStore8[21] <= WeightsStore8[637];
			WeightsStore8[22] <= WeightsStore8[638];
			WeightsStore8[23] <= WeightsStore8[639];
			WeightsStore8[24] <= WeightsStore8[640];
			WeightsStore8[25] <= WeightsStore8[641];
			WeightsStore8[26] <= WeightsStore8[642];
			WeightsStore8[27] <= WeightsStore8[643];
			WeightsStore9[0] <= WeightsStore9[616];
			WeightsStore9[1] <= WeightsStore9[617];
			WeightsStore9[2] <= WeightsStore9[618];
			WeightsStore9[3] <= WeightsStore9[619];
			WeightsStore9[4] <= WeightsStore9[620];
			WeightsStore9[5] <= WeightsStore9[621];
			WeightsStore9[6] <= WeightsStore9[622];
			WeightsStore9[7] <= WeightsStore9[623];
			WeightsStore9[8] <= WeightsStore9[624];
			WeightsStore9[9] <= WeightsStore9[625];
			WeightsStore9[10] <= WeightsStore9[626];
			WeightsStore9[11] <= WeightsStore9[627];
			WeightsStore9[12] <= WeightsStore9[628];
			WeightsStore9[13] <= WeightsStore9[629];
			WeightsStore9[14] <= WeightsStore9[630];
			WeightsStore9[15] <= WeightsStore9[631];
			WeightsStore9[16] <= WeightsStore9[632];
			WeightsStore9[17] <= WeightsStore9[633];
			WeightsStore9[18] <= WeightsStore9[634];
			WeightsStore9[19] <= WeightsStore9[635];
			WeightsStore9[20] <= WeightsStore9[636];
			WeightsStore9[21] <= WeightsStore9[637];
			WeightsStore9[22] <= WeightsStore9[638];
			WeightsStore9[23] <= WeightsStore9[639];
			WeightsStore9[24] <= WeightsStore9[640];
			WeightsStore9[25] <= WeightsStore9[641];
			WeightsStore9[26] <= WeightsStore9[642];
			WeightsStore9[27] <= WeightsStore9[643];
		end else if(switchCounter == 32'd160)begin
			PixelsStore[0] <= PixelsStore[644];
			PixelsStore[1] <= PixelsStore[645];
			PixelsStore[2] <= PixelsStore[646];
			PixelsStore[3] <= PixelsStore[647];
			PixelsStore[4] <= PixelsStore[648];
			PixelsStore[5] <= PixelsStore[649];
			PixelsStore[6] <= PixelsStore[650];
			PixelsStore[7] <= PixelsStore[651];
			PixelsStore[8] <= PixelsStore[652];
			PixelsStore[9] <= PixelsStore[653];
			PixelsStore[10] <= PixelsStore[654];
			PixelsStore[11] <= PixelsStore[655];
			PixelsStore[12] <= PixelsStore[656];
			PixelsStore[13] <= PixelsStore[657];
			PixelsStore[14] <= PixelsStore[658];
			PixelsStore[15] <= PixelsStore[659];
			PixelsStore[16] <= PixelsStore[660];
			PixelsStore[17] <= PixelsStore[661];
			PixelsStore[18] <= PixelsStore[662];
			PixelsStore[19] <= PixelsStore[663];
			PixelsStore[20] <= PixelsStore[664];
			PixelsStore[21] <= PixelsStore[665];
			PixelsStore[22] <= PixelsStore[666];
			PixelsStore[23] <= PixelsStore[667];
			PixelsStore[24] <= PixelsStore[668];
			PixelsStore[25] <= PixelsStore[669];
			PixelsStore[26] <= PixelsStore[670];
			PixelsStore[27] <= PixelsStore[671];
			WeightsStore0[0] <= WeightsStore0[644];
			WeightsStore0[1] <= WeightsStore0[645];
			WeightsStore0[2] <= WeightsStore0[646];
			WeightsStore0[3] <= WeightsStore0[647];
			WeightsStore0[4] <= WeightsStore0[648];
			WeightsStore0[5] <= WeightsStore0[649];
			WeightsStore0[6] <= WeightsStore0[650];
			WeightsStore0[7] <= WeightsStore0[651];
			WeightsStore0[8] <= WeightsStore0[652];
			WeightsStore0[9] <= WeightsStore0[653];
			WeightsStore0[10] <= WeightsStore0[654];
			WeightsStore0[11] <= WeightsStore0[655];
			WeightsStore0[12] <= WeightsStore0[656];
			WeightsStore0[13] <= WeightsStore0[657];
			WeightsStore0[14] <= WeightsStore0[658];
			WeightsStore0[15] <= WeightsStore0[659];
			WeightsStore0[16] <= WeightsStore0[660];
			WeightsStore0[17] <= WeightsStore0[661];
			WeightsStore0[18] <= WeightsStore0[662];
			WeightsStore0[19] <= WeightsStore0[663];
			WeightsStore0[20] <= WeightsStore0[664];
			WeightsStore0[21] <= WeightsStore0[665];
			WeightsStore0[22] <= WeightsStore0[666];
			WeightsStore0[23] <= WeightsStore0[667];
			WeightsStore0[24] <= WeightsStore0[668];
			WeightsStore0[25] <= WeightsStore0[669];
			WeightsStore0[26] <= WeightsStore0[670];
			WeightsStore0[27] <= WeightsStore0[671];
			WeightsStore1[0] <= WeightsStore1[644];
			WeightsStore1[1] <= WeightsStore1[645];
			WeightsStore1[2] <= WeightsStore1[646];
			WeightsStore1[3] <= WeightsStore1[647];
			WeightsStore1[4] <= WeightsStore1[648];
			WeightsStore1[5] <= WeightsStore1[649];
			WeightsStore1[6] <= WeightsStore1[650];
			WeightsStore1[7] <= WeightsStore1[651];
			WeightsStore1[8] <= WeightsStore1[652];
			WeightsStore1[9] <= WeightsStore1[653];
			WeightsStore1[10] <= WeightsStore1[654];
			WeightsStore1[11] <= WeightsStore1[655];
			WeightsStore1[12] <= WeightsStore1[656];
			WeightsStore1[13] <= WeightsStore1[657];
			WeightsStore1[14] <= WeightsStore1[658];
			WeightsStore1[15] <= WeightsStore1[659];
			WeightsStore1[16] <= WeightsStore1[660];
			WeightsStore1[17] <= WeightsStore1[661];
			WeightsStore1[18] <= WeightsStore1[662];
			WeightsStore1[19] <= WeightsStore1[663];
			WeightsStore1[20] <= WeightsStore1[664];
			WeightsStore1[21] <= WeightsStore1[665];
			WeightsStore1[22] <= WeightsStore1[666];
			WeightsStore1[23] <= WeightsStore1[667];
			WeightsStore1[24] <= WeightsStore1[668];
			WeightsStore1[25] <= WeightsStore1[669];
			WeightsStore1[26] <= WeightsStore1[670];
			WeightsStore1[27] <= WeightsStore1[671];
			WeightsStore2[0] <= WeightsStore2[644];
			WeightsStore2[1] <= WeightsStore2[645];
			WeightsStore2[2] <= WeightsStore2[646];
			WeightsStore2[3] <= WeightsStore2[647];
			WeightsStore2[4] <= WeightsStore2[648];
			WeightsStore2[5] <= WeightsStore2[649];
			WeightsStore2[6] <= WeightsStore2[650];
			WeightsStore2[7] <= WeightsStore2[651];
			WeightsStore2[8] <= WeightsStore2[652];
			WeightsStore2[9] <= WeightsStore2[653];
			WeightsStore2[10] <= WeightsStore2[654];
			WeightsStore2[11] <= WeightsStore2[655];
			WeightsStore2[12] <= WeightsStore2[656];
			WeightsStore2[13] <= WeightsStore2[657];
			WeightsStore2[14] <= WeightsStore2[658];
			WeightsStore2[15] <= WeightsStore2[659];
			WeightsStore2[16] <= WeightsStore2[660];
			WeightsStore2[17] <= WeightsStore2[661];
			WeightsStore2[18] <= WeightsStore2[662];
			WeightsStore2[19] <= WeightsStore2[663];
			WeightsStore2[20] <= WeightsStore2[664];
			WeightsStore2[21] <= WeightsStore2[665];
			WeightsStore2[22] <= WeightsStore2[666];
			WeightsStore2[23] <= WeightsStore2[667];
			WeightsStore2[24] <= WeightsStore2[668];
			WeightsStore2[25] <= WeightsStore2[669];
			WeightsStore2[26] <= WeightsStore2[670];
			WeightsStore2[27] <= WeightsStore2[671];
			WeightsStore3[0] <= WeightsStore3[644];
			WeightsStore3[1] <= WeightsStore3[645];
			WeightsStore3[2] <= WeightsStore3[646];
			WeightsStore3[3] <= WeightsStore3[647];
			WeightsStore3[4] <= WeightsStore3[648];
			WeightsStore3[5] <= WeightsStore3[649];
			WeightsStore3[6] <= WeightsStore3[650];
			WeightsStore3[7] <= WeightsStore3[651];
			WeightsStore3[8] <= WeightsStore3[652];
			WeightsStore3[9] <= WeightsStore3[653];
			WeightsStore3[10] <= WeightsStore3[654];
			WeightsStore3[11] <= WeightsStore3[655];
			WeightsStore3[12] <= WeightsStore3[656];
			WeightsStore3[13] <= WeightsStore3[657];
			WeightsStore3[14] <= WeightsStore3[658];
			WeightsStore3[15] <= WeightsStore3[659];
			WeightsStore3[16] <= WeightsStore3[660];
			WeightsStore3[17] <= WeightsStore3[661];
			WeightsStore3[18] <= WeightsStore3[662];
			WeightsStore3[19] <= WeightsStore3[663];
			WeightsStore3[20] <= WeightsStore3[664];
			WeightsStore3[21] <= WeightsStore3[665];
			WeightsStore3[22] <= WeightsStore3[666];
			WeightsStore3[23] <= WeightsStore3[667];
			WeightsStore3[24] <= WeightsStore3[668];
			WeightsStore3[25] <= WeightsStore3[669];
			WeightsStore3[26] <= WeightsStore3[670];
			WeightsStore3[27] <= WeightsStore3[671];
			WeightsStore4[0] <= WeightsStore4[644];
			WeightsStore4[1] <= WeightsStore4[645];
			WeightsStore4[2] <= WeightsStore4[646];
			WeightsStore4[3] <= WeightsStore4[647];
			WeightsStore4[4] <= WeightsStore4[648];
			WeightsStore4[5] <= WeightsStore4[649];
			WeightsStore4[6] <= WeightsStore4[650];
			WeightsStore4[7] <= WeightsStore4[651];
			WeightsStore4[8] <= WeightsStore4[652];
			WeightsStore4[9] <= WeightsStore4[653];
			WeightsStore4[10] <= WeightsStore4[654];
			WeightsStore4[11] <= WeightsStore4[655];
			WeightsStore4[12] <= WeightsStore4[656];
			WeightsStore4[13] <= WeightsStore4[657];
			WeightsStore4[14] <= WeightsStore4[658];
			WeightsStore4[15] <= WeightsStore4[659];
			WeightsStore4[16] <= WeightsStore4[660];
			WeightsStore4[17] <= WeightsStore4[661];
			WeightsStore4[18] <= WeightsStore4[662];
			WeightsStore4[19] <= WeightsStore4[663];
			WeightsStore4[20] <= WeightsStore4[664];
			WeightsStore4[21] <= WeightsStore4[665];
			WeightsStore4[22] <= WeightsStore4[666];
			WeightsStore4[23] <= WeightsStore4[667];
			WeightsStore4[24] <= WeightsStore4[668];
			WeightsStore4[25] <= WeightsStore4[669];
			WeightsStore4[26] <= WeightsStore4[670];
			WeightsStore4[27] <= WeightsStore4[671];
			WeightsStore5[0] <= WeightsStore5[644];
			WeightsStore5[1] <= WeightsStore5[645];
			WeightsStore5[2] <= WeightsStore5[646];
			WeightsStore5[3] <= WeightsStore5[647];
			WeightsStore5[4] <= WeightsStore5[648];
			WeightsStore5[5] <= WeightsStore5[649];
			WeightsStore5[6] <= WeightsStore5[650];
			WeightsStore5[7] <= WeightsStore5[651];
			WeightsStore5[8] <= WeightsStore5[652];
			WeightsStore5[9] <= WeightsStore5[653];
			WeightsStore5[10] <= WeightsStore5[654];
			WeightsStore5[11] <= WeightsStore5[655];
			WeightsStore5[12] <= WeightsStore5[656];
			WeightsStore5[13] <= WeightsStore5[657];
			WeightsStore5[14] <= WeightsStore5[658];
			WeightsStore5[15] <= WeightsStore5[659];
			WeightsStore5[16] <= WeightsStore5[660];
			WeightsStore5[17] <= WeightsStore5[661];
			WeightsStore5[18] <= WeightsStore5[662];
			WeightsStore5[19] <= WeightsStore5[663];
			WeightsStore5[20] <= WeightsStore5[664];
			WeightsStore5[21] <= WeightsStore5[665];
			WeightsStore5[22] <= WeightsStore5[666];
			WeightsStore5[23] <= WeightsStore5[667];
			WeightsStore5[24] <= WeightsStore5[668];
			WeightsStore5[25] <= WeightsStore5[669];
			WeightsStore5[26] <= WeightsStore5[670];
			WeightsStore5[27] <= WeightsStore5[671];
			WeightsStore6[0] <= WeightsStore6[644];
			WeightsStore6[1] <= WeightsStore6[645];
			WeightsStore6[2] <= WeightsStore6[646];
			WeightsStore6[3] <= WeightsStore6[647];
			WeightsStore6[4] <= WeightsStore6[648];
			WeightsStore6[5] <= WeightsStore6[649];
			WeightsStore6[6] <= WeightsStore6[650];
			WeightsStore6[7] <= WeightsStore6[651];
			WeightsStore6[8] <= WeightsStore6[652];
			WeightsStore6[9] <= WeightsStore6[653];
			WeightsStore6[10] <= WeightsStore6[654];
			WeightsStore6[11] <= WeightsStore6[655];
			WeightsStore6[12] <= WeightsStore6[656];
			WeightsStore6[13] <= WeightsStore6[657];
			WeightsStore6[14] <= WeightsStore6[658];
			WeightsStore6[15] <= WeightsStore6[659];
			WeightsStore6[16] <= WeightsStore6[660];
			WeightsStore6[17] <= WeightsStore6[661];
			WeightsStore6[18] <= WeightsStore6[662];
			WeightsStore6[19] <= WeightsStore6[663];
			WeightsStore6[20] <= WeightsStore6[664];
			WeightsStore6[21] <= WeightsStore6[665];
			WeightsStore6[22] <= WeightsStore6[666];
			WeightsStore6[23] <= WeightsStore6[667];
			WeightsStore6[24] <= WeightsStore6[668];
			WeightsStore6[25] <= WeightsStore6[669];
			WeightsStore6[26] <= WeightsStore6[670];
			WeightsStore6[27] <= WeightsStore6[671];
			WeightsStore7[0] <= WeightsStore7[644];
			WeightsStore7[1] <= WeightsStore7[645];
			WeightsStore7[2] <= WeightsStore7[646];
			WeightsStore7[3] <= WeightsStore7[647];
			WeightsStore7[4] <= WeightsStore7[648];
			WeightsStore7[5] <= WeightsStore7[649];
			WeightsStore7[6] <= WeightsStore7[650];
			WeightsStore7[7] <= WeightsStore7[651];
			WeightsStore7[8] <= WeightsStore7[652];
			WeightsStore7[9] <= WeightsStore7[653];
			WeightsStore7[10] <= WeightsStore7[654];
			WeightsStore7[11] <= WeightsStore7[655];
			WeightsStore7[12] <= WeightsStore7[656];
			WeightsStore7[13] <= WeightsStore7[657];
			WeightsStore7[14] <= WeightsStore7[658];
			WeightsStore7[15] <= WeightsStore7[659];
			WeightsStore7[16] <= WeightsStore7[660];
			WeightsStore7[17] <= WeightsStore7[661];
			WeightsStore7[18] <= WeightsStore7[662];
			WeightsStore7[19] <= WeightsStore7[663];
			WeightsStore7[20] <= WeightsStore7[664];
			WeightsStore7[21] <= WeightsStore7[665];
			WeightsStore7[22] <= WeightsStore7[666];
			WeightsStore7[23] <= WeightsStore7[667];
			WeightsStore7[24] <= WeightsStore7[668];
			WeightsStore7[25] <= WeightsStore7[669];
			WeightsStore7[26] <= WeightsStore7[670];
			WeightsStore7[27] <= WeightsStore7[671];
			WeightsStore8[0] <= WeightsStore8[644];
			WeightsStore8[1] <= WeightsStore8[645];
			WeightsStore8[2] <= WeightsStore8[646];
			WeightsStore8[3] <= WeightsStore8[647];
			WeightsStore8[4] <= WeightsStore8[648];
			WeightsStore8[5] <= WeightsStore8[649];
			WeightsStore8[6] <= WeightsStore8[650];
			WeightsStore8[7] <= WeightsStore8[651];
			WeightsStore8[8] <= WeightsStore8[652];
			WeightsStore8[9] <= WeightsStore8[653];
			WeightsStore8[10] <= WeightsStore8[654];
			WeightsStore8[11] <= WeightsStore8[655];
			WeightsStore8[12] <= WeightsStore8[656];
			WeightsStore8[13] <= WeightsStore8[657];
			WeightsStore8[14] <= WeightsStore8[658];
			WeightsStore8[15] <= WeightsStore8[659];
			WeightsStore8[16] <= WeightsStore8[660];
			WeightsStore8[17] <= WeightsStore8[661];
			WeightsStore8[18] <= WeightsStore8[662];
			WeightsStore8[19] <= WeightsStore8[663];
			WeightsStore8[20] <= WeightsStore8[664];
			WeightsStore8[21] <= WeightsStore8[665];
			WeightsStore8[22] <= WeightsStore8[666];
			WeightsStore8[23] <= WeightsStore8[667];
			WeightsStore8[24] <= WeightsStore8[668];
			WeightsStore8[25] <= WeightsStore8[669];
			WeightsStore8[26] <= WeightsStore8[670];
			WeightsStore8[27] <= WeightsStore8[671];
			WeightsStore9[0] <= WeightsStore9[644];
			WeightsStore9[1] <= WeightsStore9[645];
			WeightsStore9[2] <= WeightsStore9[646];
			WeightsStore9[3] <= WeightsStore9[647];
			WeightsStore9[4] <= WeightsStore9[648];
			WeightsStore9[5] <= WeightsStore9[649];
			WeightsStore9[6] <= WeightsStore9[650];
			WeightsStore9[7] <= WeightsStore9[651];
			WeightsStore9[8] <= WeightsStore9[652];
			WeightsStore9[9] <= WeightsStore9[653];
			WeightsStore9[10] <= WeightsStore9[654];
			WeightsStore9[11] <= WeightsStore9[655];
			WeightsStore9[12] <= WeightsStore9[656];
			WeightsStore9[13] <= WeightsStore9[657];
			WeightsStore9[14] <= WeightsStore9[658];
			WeightsStore9[15] <= WeightsStore9[659];
			WeightsStore9[16] <= WeightsStore9[660];
			WeightsStore9[17] <= WeightsStore9[661];
			WeightsStore9[18] <= WeightsStore9[662];
			WeightsStore9[19] <= WeightsStore9[663];
			WeightsStore9[20] <= WeightsStore9[664];
			WeightsStore9[21] <= WeightsStore9[665];
			WeightsStore9[22] <= WeightsStore9[666];
			WeightsStore9[23] <= WeightsStore9[667];
			WeightsStore9[24] <= WeightsStore9[668];
			WeightsStore9[25] <= WeightsStore9[669];
			WeightsStore9[26] <= WeightsStore9[670];
			WeightsStore9[27] <= WeightsStore9[671];
		end else if(switchCounter == 32'd167)begin
			PixelsStore[0] <= PixelsStore[672];
			PixelsStore[1] <= PixelsStore[673];
			PixelsStore[2] <= PixelsStore[674];
			PixelsStore[3] <= PixelsStore[675];
			PixelsStore[4] <= PixelsStore[676];
			PixelsStore[5] <= PixelsStore[677];
			PixelsStore[6] <= PixelsStore[678];
			PixelsStore[7] <= PixelsStore[679];
			PixelsStore[8] <= PixelsStore[680];
			PixelsStore[9] <= PixelsStore[681];
			PixelsStore[10] <= PixelsStore[682];
			PixelsStore[11] <= PixelsStore[683];
			PixelsStore[12] <= PixelsStore[684];
			PixelsStore[13] <= PixelsStore[685];
			PixelsStore[14] <= PixelsStore[686];
			PixelsStore[15] <= PixelsStore[687];
			PixelsStore[16] <= PixelsStore[688];
			PixelsStore[17] <= PixelsStore[689];
			PixelsStore[18] <= PixelsStore[690];
			PixelsStore[19] <= PixelsStore[691];
			PixelsStore[20] <= PixelsStore[692];
			PixelsStore[21] <= PixelsStore[693];
			PixelsStore[22] <= PixelsStore[694];
			PixelsStore[23] <= PixelsStore[695];
			PixelsStore[24] <= PixelsStore[696];
			PixelsStore[25] <= PixelsStore[697];
			PixelsStore[26] <= PixelsStore[698];
			PixelsStore[27] <= PixelsStore[699];
			WeightsStore0[0] <= WeightsStore0[672];
			WeightsStore0[1] <= WeightsStore0[673];
			WeightsStore0[2] <= WeightsStore0[674];
			WeightsStore0[3] <= WeightsStore0[675];
			WeightsStore0[4] <= WeightsStore0[676];
			WeightsStore0[5] <= WeightsStore0[677];
			WeightsStore0[6] <= WeightsStore0[678];
			WeightsStore0[7] <= WeightsStore0[679];
			WeightsStore0[8] <= WeightsStore0[680];
			WeightsStore0[9] <= WeightsStore0[681];
			WeightsStore0[10] <= WeightsStore0[682];
			WeightsStore0[11] <= WeightsStore0[683];
			WeightsStore0[12] <= WeightsStore0[684];
			WeightsStore0[13] <= WeightsStore0[685];
			WeightsStore0[14] <= WeightsStore0[686];
			WeightsStore0[15] <= WeightsStore0[687];
			WeightsStore0[16] <= WeightsStore0[688];
			WeightsStore0[17] <= WeightsStore0[689];
			WeightsStore0[18] <= WeightsStore0[690];
			WeightsStore0[19] <= WeightsStore0[691];
			WeightsStore0[20] <= WeightsStore0[692];
			WeightsStore0[21] <= WeightsStore0[693];
			WeightsStore0[22] <= WeightsStore0[694];
			WeightsStore0[23] <= WeightsStore0[695];
			WeightsStore0[24] <= WeightsStore0[696];
			WeightsStore0[25] <= WeightsStore0[697];
			WeightsStore0[26] <= WeightsStore0[698];
			WeightsStore0[27] <= WeightsStore0[699];
			WeightsStore1[0] <= WeightsStore1[672];
			WeightsStore1[1] <= WeightsStore1[673];
			WeightsStore1[2] <= WeightsStore1[674];
			WeightsStore1[3] <= WeightsStore1[675];
			WeightsStore1[4] <= WeightsStore1[676];
			WeightsStore1[5] <= WeightsStore1[677];
			WeightsStore1[6] <= WeightsStore1[678];
			WeightsStore1[7] <= WeightsStore1[679];
			WeightsStore1[8] <= WeightsStore1[680];
			WeightsStore1[9] <= WeightsStore1[681];
			WeightsStore1[10] <= WeightsStore1[682];
			WeightsStore1[11] <= WeightsStore1[683];
			WeightsStore1[12] <= WeightsStore1[684];
			WeightsStore1[13] <= WeightsStore1[685];
			WeightsStore1[14] <= WeightsStore1[686];
			WeightsStore1[15] <= WeightsStore1[687];
			WeightsStore1[16] <= WeightsStore1[688];
			WeightsStore1[17] <= WeightsStore1[689];
			WeightsStore1[18] <= WeightsStore1[690];
			WeightsStore1[19] <= WeightsStore1[691];
			WeightsStore1[20] <= WeightsStore1[692];
			WeightsStore1[21] <= WeightsStore1[693];
			WeightsStore1[22] <= WeightsStore1[694];
			WeightsStore1[23] <= WeightsStore1[695];
			WeightsStore1[24] <= WeightsStore1[696];
			WeightsStore1[25] <= WeightsStore1[697];
			WeightsStore1[26] <= WeightsStore1[698];
			WeightsStore1[27] <= WeightsStore1[699];
			WeightsStore2[0] <= WeightsStore2[672];
			WeightsStore2[1] <= WeightsStore2[673];
			WeightsStore2[2] <= WeightsStore2[674];
			WeightsStore2[3] <= WeightsStore2[675];
			WeightsStore2[4] <= WeightsStore2[676];
			WeightsStore2[5] <= WeightsStore2[677];
			WeightsStore2[6] <= WeightsStore2[678];
			WeightsStore2[7] <= WeightsStore2[679];
			WeightsStore2[8] <= WeightsStore2[680];
			WeightsStore2[9] <= WeightsStore2[681];
			WeightsStore2[10] <= WeightsStore2[682];
			WeightsStore2[11] <= WeightsStore2[683];
			WeightsStore2[12] <= WeightsStore2[684];
			WeightsStore2[13] <= WeightsStore2[685];
			WeightsStore2[14] <= WeightsStore2[686];
			WeightsStore2[15] <= WeightsStore2[687];
			WeightsStore2[16] <= WeightsStore2[688];
			WeightsStore2[17] <= WeightsStore2[689];
			WeightsStore2[18] <= WeightsStore2[690];
			WeightsStore2[19] <= WeightsStore2[691];
			WeightsStore2[20] <= WeightsStore2[692];
			WeightsStore2[21] <= WeightsStore2[693];
			WeightsStore2[22] <= WeightsStore2[694];
			WeightsStore2[23] <= WeightsStore2[695];
			WeightsStore2[24] <= WeightsStore2[696];
			WeightsStore2[25] <= WeightsStore2[697];
			WeightsStore2[26] <= WeightsStore2[698];
			WeightsStore2[27] <= WeightsStore2[699];
			WeightsStore3[0] <= WeightsStore3[672];
			WeightsStore3[1] <= WeightsStore3[673];
			WeightsStore3[2] <= WeightsStore3[674];
			WeightsStore3[3] <= WeightsStore3[675];
			WeightsStore3[4] <= WeightsStore3[676];
			WeightsStore3[5] <= WeightsStore3[677];
			WeightsStore3[6] <= WeightsStore3[678];
			WeightsStore3[7] <= WeightsStore3[679];
			WeightsStore3[8] <= WeightsStore3[680];
			WeightsStore3[9] <= WeightsStore3[681];
			WeightsStore3[10] <= WeightsStore3[682];
			WeightsStore3[11] <= WeightsStore3[683];
			WeightsStore3[12] <= WeightsStore3[684];
			WeightsStore3[13] <= WeightsStore3[685];
			WeightsStore3[14] <= WeightsStore3[686];
			WeightsStore3[15] <= WeightsStore3[687];
			WeightsStore3[16] <= WeightsStore3[688];
			WeightsStore3[17] <= WeightsStore3[689];
			WeightsStore3[18] <= WeightsStore3[690];
			WeightsStore3[19] <= WeightsStore3[691];
			WeightsStore3[20] <= WeightsStore3[692];
			WeightsStore3[21] <= WeightsStore3[693];
			WeightsStore3[22] <= WeightsStore3[694];
			WeightsStore3[23] <= WeightsStore3[695];
			WeightsStore3[24] <= WeightsStore3[696];
			WeightsStore3[25] <= WeightsStore3[697];
			WeightsStore3[26] <= WeightsStore3[698];
			WeightsStore3[27] <= WeightsStore3[699];
			WeightsStore4[0] <= WeightsStore4[672];
			WeightsStore4[1] <= WeightsStore4[673];
			WeightsStore4[2] <= WeightsStore4[674];
			WeightsStore4[3] <= WeightsStore4[675];
			WeightsStore4[4] <= WeightsStore4[676];
			WeightsStore4[5] <= WeightsStore4[677];
			WeightsStore4[6] <= WeightsStore4[678];
			WeightsStore4[7] <= WeightsStore4[679];
			WeightsStore4[8] <= WeightsStore4[680];
			WeightsStore4[9] <= WeightsStore4[681];
			WeightsStore4[10] <= WeightsStore4[682];
			WeightsStore4[11] <= WeightsStore4[683];
			WeightsStore4[12] <= WeightsStore4[684];
			WeightsStore4[13] <= WeightsStore4[685];
			WeightsStore4[14] <= WeightsStore4[686];
			WeightsStore4[15] <= WeightsStore4[687];
			WeightsStore4[16] <= WeightsStore4[688];
			WeightsStore4[17] <= WeightsStore4[689];
			WeightsStore4[18] <= WeightsStore4[690];
			WeightsStore4[19] <= WeightsStore4[691];
			WeightsStore4[20] <= WeightsStore4[692];
			WeightsStore4[21] <= WeightsStore4[693];
			WeightsStore4[22] <= WeightsStore4[694];
			WeightsStore4[23] <= WeightsStore4[695];
			WeightsStore4[24] <= WeightsStore4[696];
			WeightsStore4[25] <= WeightsStore4[697];
			WeightsStore4[26] <= WeightsStore4[698];
			WeightsStore4[27] <= WeightsStore4[699];
			WeightsStore5[0] <= WeightsStore5[672];
			WeightsStore5[1] <= WeightsStore5[673];
			WeightsStore5[2] <= WeightsStore5[674];
			WeightsStore5[3] <= WeightsStore5[675];
			WeightsStore5[4] <= WeightsStore5[676];
			WeightsStore5[5] <= WeightsStore5[677];
			WeightsStore5[6] <= WeightsStore5[678];
			WeightsStore5[7] <= WeightsStore5[679];
			WeightsStore5[8] <= WeightsStore5[680];
			WeightsStore5[9] <= WeightsStore5[681];
			WeightsStore5[10] <= WeightsStore5[682];
			WeightsStore5[11] <= WeightsStore5[683];
			WeightsStore5[12] <= WeightsStore5[684];
			WeightsStore5[13] <= WeightsStore5[685];
			WeightsStore5[14] <= WeightsStore5[686];
			WeightsStore5[15] <= WeightsStore5[687];
			WeightsStore5[16] <= WeightsStore5[688];
			WeightsStore5[17] <= WeightsStore5[689];
			WeightsStore5[18] <= WeightsStore5[690];
			WeightsStore5[19] <= WeightsStore5[691];
			WeightsStore5[20] <= WeightsStore5[692];
			WeightsStore5[21] <= WeightsStore5[693];
			WeightsStore5[22] <= WeightsStore5[694];
			WeightsStore5[23] <= WeightsStore5[695];
			WeightsStore5[24] <= WeightsStore5[696];
			WeightsStore5[25] <= WeightsStore5[697];
			WeightsStore5[26] <= WeightsStore5[698];
			WeightsStore5[27] <= WeightsStore5[699];
			WeightsStore6[0] <= WeightsStore6[672];
			WeightsStore6[1] <= WeightsStore6[673];
			WeightsStore6[2] <= WeightsStore6[674];
			WeightsStore6[3] <= WeightsStore6[675];
			WeightsStore6[4] <= WeightsStore6[676];
			WeightsStore6[5] <= WeightsStore6[677];
			WeightsStore6[6] <= WeightsStore6[678];
			WeightsStore6[7] <= WeightsStore6[679];
			WeightsStore6[8] <= WeightsStore6[680];
			WeightsStore6[9] <= WeightsStore6[681];
			WeightsStore6[10] <= WeightsStore6[682];
			WeightsStore6[11] <= WeightsStore6[683];
			WeightsStore6[12] <= WeightsStore6[684];
			WeightsStore6[13] <= WeightsStore6[685];
			WeightsStore6[14] <= WeightsStore6[686];
			WeightsStore6[15] <= WeightsStore6[687];
			WeightsStore6[16] <= WeightsStore6[688];
			WeightsStore6[17] <= WeightsStore6[689];
			WeightsStore6[18] <= WeightsStore6[690];
			WeightsStore6[19] <= WeightsStore6[691];
			WeightsStore6[20] <= WeightsStore6[692];
			WeightsStore6[21] <= WeightsStore6[693];
			WeightsStore6[22] <= WeightsStore6[694];
			WeightsStore6[23] <= WeightsStore6[695];
			WeightsStore6[24] <= WeightsStore6[696];
			WeightsStore6[25] <= WeightsStore6[697];
			WeightsStore6[26] <= WeightsStore6[698];
			WeightsStore6[27] <= WeightsStore6[699];
			WeightsStore7[0] <= WeightsStore7[672];
			WeightsStore7[1] <= WeightsStore7[673];
			WeightsStore7[2] <= WeightsStore7[674];
			WeightsStore7[3] <= WeightsStore7[675];
			WeightsStore7[4] <= WeightsStore7[676];
			WeightsStore7[5] <= WeightsStore7[677];
			WeightsStore7[6] <= WeightsStore7[678];
			WeightsStore7[7] <= WeightsStore7[679];
			WeightsStore7[8] <= WeightsStore7[680];
			WeightsStore7[9] <= WeightsStore7[681];
			WeightsStore7[10] <= WeightsStore7[682];
			WeightsStore7[11] <= WeightsStore7[683];
			WeightsStore7[12] <= WeightsStore7[684];
			WeightsStore7[13] <= WeightsStore7[685];
			WeightsStore7[14] <= WeightsStore7[686];
			WeightsStore7[15] <= WeightsStore7[687];
			WeightsStore7[16] <= WeightsStore7[688];
			WeightsStore7[17] <= WeightsStore7[689];
			WeightsStore7[18] <= WeightsStore7[690];
			WeightsStore7[19] <= WeightsStore7[691];
			WeightsStore7[20] <= WeightsStore7[692];
			WeightsStore7[21] <= WeightsStore7[693];
			WeightsStore7[22] <= WeightsStore7[694];
			WeightsStore7[23] <= WeightsStore7[695];
			WeightsStore7[24] <= WeightsStore7[696];
			WeightsStore7[25] <= WeightsStore7[697];
			WeightsStore7[26] <= WeightsStore7[698];
			WeightsStore7[27] <= WeightsStore7[699];
			WeightsStore8[0] <= WeightsStore8[672];
			WeightsStore8[1] <= WeightsStore8[673];
			WeightsStore8[2] <= WeightsStore8[674];
			WeightsStore8[3] <= WeightsStore8[675];
			WeightsStore8[4] <= WeightsStore8[676];
			WeightsStore8[5] <= WeightsStore8[677];
			WeightsStore8[6] <= WeightsStore8[678];
			WeightsStore8[7] <= WeightsStore8[679];
			WeightsStore8[8] <= WeightsStore8[680];
			WeightsStore8[9] <= WeightsStore8[681];
			WeightsStore8[10] <= WeightsStore8[682];
			WeightsStore8[11] <= WeightsStore8[683];
			WeightsStore8[12] <= WeightsStore8[684];
			WeightsStore8[13] <= WeightsStore8[685];
			WeightsStore8[14] <= WeightsStore8[686];
			WeightsStore8[15] <= WeightsStore8[687];
			WeightsStore8[16] <= WeightsStore8[688];
			WeightsStore8[17] <= WeightsStore8[689];
			WeightsStore8[18] <= WeightsStore8[690];
			WeightsStore8[19] <= WeightsStore8[691];
			WeightsStore8[20] <= WeightsStore8[692];
			WeightsStore8[21] <= WeightsStore8[693];
			WeightsStore8[22] <= WeightsStore8[694];
			WeightsStore8[23] <= WeightsStore8[695];
			WeightsStore8[24] <= WeightsStore8[696];
			WeightsStore8[25] <= WeightsStore8[697];
			WeightsStore8[26] <= WeightsStore8[698];
			WeightsStore8[27] <= WeightsStore8[699];
			WeightsStore9[0] <= WeightsStore9[672];
			WeightsStore9[1] <= WeightsStore9[673];
			WeightsStore9[2] <= WeightsStore9[674];
			WeightsStore9[3] <= WeightsStore9[675];
			WeightsStore9[4] <= WeightsStore9[676];
			WeightsStore9[5] <= WeightsStore9[677];
			WeightsStore9[6] <= WeightsStore9[678];
			WeightsStore9[7] <= WeightsStore9[679];
			WeightsStore9[8] <= WeightsStore9[680];
			WeightsStore9[9] <= WeightsStore9[681];
			WeightsStore9[10] <= WeightsStore9[682];
			WeightsStore9[11] <= WeightsStore9[683];
			WeightsStore9[12] <= WeightsStore9[684];
			WeightsStore9[13] <= WeightsStore9[685];
			WeightsStore9[14] <= WeightsStore9[686];
			WeightsStore9[15] <= WeightsStore9[687];
			WeightsStore9[16] <= WeightsStore9[688];
			WeightsStore9[17] <= WeightsStore9[689];
			WeightsStore9[18] <= WeightsStore9[690];
			WeightsStore9[19] <= WeightsStore9[691];
			WeightsStore9[20] <= WeightsStore9[692];
			WeightsStore9[21] <= WeightsStore9[693];
			WeightsStore9[22] <= WeightsStore9[694];
			WeightsStore9[23] <= WeightsStore9[695];
			WeightsStore9[24] <= WeightsStore9[696];
			WeightsStore9[25] <= WeightsStore9[697];
			WeightsStore9[26] <= WeightsStore9[698];
			WeightsStore9[27] <= WeightsStore9[699];
		end else if(switchCounter == 32'd174)begin
			PixelsStore[0] <= PixelsStore[700];
			PixelsStore[1] <= PixelsStore[701];
			PixelsStore[2] <= PixelsStore[702];
			PixelsStore[3] <= PixelsStore[703];
			PixelsStore[4] <= PixelsStore[704];
			PixelsStore[5] <= PixelsStore[705];
			PixelsStore[6] <= PixelsStore[706];
			PixelsStore[7] <= PixelsStore[707];
			PixelsStore[8] <= PixelsStore[708];
			PixelsStore[9] <= PixelsStore[709];
			PixelsStore[10] <= PixelsStore[710];
			PixelsStore[11] <= PixelsStore[711];
			PixelsStore[12] <= PixelsStore[712];
			PixelsStore[13] <= PixelsStore[713];
			PixelsStore[14] <= PixelsStore[714];
			PixelsStore[15] <= PixelsStore[715];
			PixelsStore[16] <= PixelsStore[716];
			PixelsStore[17] <= PixelsStore[717];
			PixelsStore[18] <= PixelsStore[718];
			PixelsStore[19] <= PixelsStore[719];
			PixelsStore[20] <= PixelsStore[720];
			PixelsStore[21] <= PixelsStore[721];
			PixelsStore[22] <= PixelsStore[722];
			PixelsStore[23] <= PixelsStore[723];
			PixelsStore[24] <= PixelsStore[724];
			PixelsStore[25] <= PixelsStore[725];
			PixelsStore[26] <= PixelsStore[726];
			PixelsStore[27] <= PixelsStore[727];
			WeightsStore0[0] <= WeightsStore0[700];
			WeightsStore0[1] <= WeightsStore0[701];
			WeightsStore0[2] <= WeightsStore0[702];
			WeightsStore0[3] <= WeightsStore0[703];
			WeightsStore0[4] <= WeightsStore0[704];
			WeightsStore0[5] <= WeightsStore0[705];
			WeightsStore0[6] <= WeightsStore0[706];
			WeightsStore0[7] <= WeightsStore0[707];
			WeightsStore0[8] <= WeightsStore0[708];
			WeightsStore0[9] <= WeightsStore0[709];
			WeightsStore0[10] <= WeightsStore0[710];
			WeightsStore0[11] <= WeightsStore0[711];
			WeightsStore0[12] <= WeightsStore0[712];
			WeightsStore0[13] <= WeightsStore0[713];
			WeightsStore0[14] <= WeightsStore0[714];
			WeightsStore0[15] <= WeightsStore0[715];
			WeightsStore0[16] <= WeightsStore0[716];
			WeightsStore0[17] <= WeightsStore0[717];
			WeightsStore0[18] <= WeightsStore0[718];
			WeightsStore0[19] <= WeightsStore0[719];
			WeightsStore0[20] <= WeightsStore0[720];
			WeightsStore0[21] <= WeightsStore0[721];
			WeightsStore0[22] <= WeightsStore0[722];
			WeightsStore0[23] <= WeightsStore0[723];
			WeightsStore0[24] <= WeightsStore0[724];
			WeightsStore0[25] <= WeightsStore0[725];
			WeightsStore0[26] <= WeightsStore0[726];
			WeightsStore0[27] <= WeightsStore0[727];
			WeightsStore1[0] <= WeightsStore1[700];
			WeightsStore1[1] <= WeightsStore1[701];
			WeightsStore1[2] <= WeightsStore1[702];
			WeightsStore1[3] <= WeightsStore1[703];
			WeightsStore1[4] <= WeightsStore1[704];
			WeightsStore1[5] <= WeightsStore1[705];
			WeightsStore1[6] <= WeightsStore1[706];
			WeightsStore1[7] <= WeightsStore1[707];
			WeightsStore1[8] <= WeightsStore1[708];
			WeightsStore1[9] <= WeightsStore1[709];
			WeightsStore1[10] <= WeightsStore1[710];
			WeightsStore1[11] <= WeightsStore1[711];
			WeightsStore1[12] <= WeightsStore1[712];
			WeightsStore1[13] <= WeightsStore1[713];
			WeightsStore1[14] <= WeightsStore1[714];
			WeightsStore1[15] <= WeightsStore1[715];
			WeightsStore1[16] <= WeightsStore1[716];
			WeightsStore1[17] <= WeightsStore1[717];
			WeightsStore1[18] <= WeightsStore1[718];
			WeightsStore1[19] <= WeightsStore1[719];
			WeightsStore1[20] <= WeightsStore1[720];
			WeightsStore1[21] <= WeightsStore1[721];
			WeightsStore1[22] <= WeightsStore1[722];
			WeightsStore1[23] <= WeightsStore1[723];
			WeightsStore1[24] <= WeightsStore1[724];
			WeightsStore1[25] <= WeightsStore1[725];
			WeightsStore1[26] <= WeightsStore1[726];
			WeightsStore1[27] <= WeightsStore1[727];
			WeightsStore2[0] <= WeightsStore2[700];
			WeightsStore2[1] <= WeightsStore2[701];
			WeightsStore2[2] <= WeightsStore2[702];
			WeightsStore2[3] <= WeightsStore2[703];
			WeightsStore2[4] <= WeightsStore2[704];
			WeightsStore2[5] <= WeightsStore2[705];
			WeightsStore2[6] <= WeightsStore2[706];
			WeightsStore2[7] <= WeightsStore2[707];
			WeightsStore2[8] <= WeightsStore2[708];
			WeightsStore2[9] <= WeightsStore2[709];
			WeightsStore2[10] <= WeightsStore2[710];
			WeightsStore2[11] <= WeightsStore2[711];
			WeightsStore2[12] <= WeightsStore2[712];
			WeightsStore2[13] <= WeightsStore2[713];
			WeightsStore2[14] <= WeightsStore2[714];
			WeightsStore2[15] <= WeightsStore2[715];
			WeightsStore2[16] <= WeightsStore2[716];
			WeightsStore2[17] <= WeightsStore2[717];
			WeightsStore2[18] <= WeightsStore2[718];
			WeightsStore2[19] <= WeightsStore2[719];
			WeightsStore2[20] <= WeightsStore2[720];
			WeightsStore2[21] <= WeightsStore2[721];
			WeightsStore2[22] <= WeightsStore2[722];
			WeightsStore2[23] <= WeightsStore2[723];
			WeightsStore2[24] <= WeightsStore2[724];
			WeightsStore2[25] <= WeightsStore2[725];
			WeightsStore2[26] <= WeightsStore2[726];
			WeightsStore2[27] <= WeightsStore2[727];
			WeightsStore3[0] <= WeightsStore3[700];
			WeightsStore3[1] <= WeightsStore3[701];
			WeightsStore3[2] <= WeightsStore3[702];
			WeightsStore3[3] <= WeightsStore3[703];
			WeightsStore3[4] <= WeightsStore3[704];
			WeightsStore3[5] <= WeightsStore3[705];
			WeightsStore3[6] <= WeightsStore3[706];
			WeightsStore3[7] <= WeightsStore3[707];
			WeightsStore3[8] <= WeightsStore3[708];
			WeightsStore3[9] <= WeightsStore3[709];
			WeightsStore3[10] <= WeightsStore3[710];
			WeightsStore3[11] <= WeightsStore3[711];
			WeightsStore3[12] <= WeightsStore3[712];
			WeightsStore3[13] <= WeightsStore3[713];
			WeightsStore3[14] <= WeightsStore3[714];
			WeightsStore3[15] <= WeightsStore3[715];
			WeightsStore3[16] <= WeightsStore3[716];
			WeightsStore3[17] <= WeightsStore3[717];
			WeightsStore3[18] <= WeightsStore3[718];
			WeightsStore3[19] <= WeightsStore3[719];
			WeightsStore3[20] <= WeightsStore3[720];
			WeightsStore3[21] <= WeightsStore3[721];
			WeightsStore3[22] <= WeightsStore3[722];
			WeightsStore3[23] <= WeightsStore3[723];
			WeightsStore3[24] <= WeightsStore3[724];
			WeightsStore3[25] <= WeightsStore3[725];
			WeightsStore3[26] <= WeightsStore3[726];
			WeightsStore3[27] <= WeightsStore3[727];
			WeightsStore4[0] <= WeightsStore4[700];
			WeightsStore4[1] <= WeightsStore4[701];
			WeightsStore4[2] <= WeightsStore4[702];
			WeightsStore4[3] <= WeightsStore4[703];
			WeightsStore4[4] <= WeightsStore4[704];
			WeightsStore4[5] <= WeightsStore4[705];
			WeightsStore4[6] <= WeightsStore4[706];
			WeightsStore4[7] <= WeightsStore4[707];
			WeightsStore4[8] <= WeightsStore4[708];
			WeightsStore4[9] <= WeightsStore4[709];
			WeightsStore4[10] <= WeightsStore4[710];
			WeightsStore4[11] <= WeightsStore4[711];
			WeightsStore4[12] <= WeightsStore4[712];
			WeightsStore4[13] <= WeightsStore4[713];
			WeightsStore4[14] <= WeightsStore4[714];
			WeightsStore4[15] <= WeightsStore4[715];
			WeightsStore4[16] <= WeightsStore4[716];
			WeightsStore4[17] <= WeightsStore4[717];
			WeightsStore4[18] <= WeightsStore4[718];
			WeightsStore4[19] <= WeightsStore4[719];
			WeightsStore4[20] <= WeightsStore4[720];
			WeightsStore4[21] <= WeightsStore4[721];
			WeightsStore4[22] <= WeightsStore4[722];
			WeightsStore4[23] <= WeightsStore4[723];
			WeightsStore4[24] <= WeightsStore4[724];
			WeightsStore4[25] <= WeightsStore4[725];
			WeightsStore4[26] <= WeightsStore4[726];
			WeightsStore4[27] <= WeightsStore4[727];
			WeightsStore5[0] <= WeightsStore5[700];
			WeightsStore5[1] <= WeightsStore5[701];
			WeightsStore5[2] <= WeightsStore5[702];
			WeightsStore5[3] <= WeightsStore5[703];
			WeightsStore5[4] <= WeightsStore5[704];
			WeightsStore5[5] <= WeightsStore5[705];
			WeightsStore5[6] <= WeightsStore5[706];
			WeightsStore5[7] <= WeightsStore5[707];
			WeightsStore5[8] <= WeightsStore5[708];
			WeightsStore5[9] <= WeightsStore5[709];
			WeightsStore5[10] <= WeightsStore5[710];
			WeightsStore5[11] <= WeightsStore5[711];
			WeightsStore5[12] <= WeightsStore5[712];
			WeightsStore5[13] <= WeightsStore5[713];
			WeightsStore5[14] <= WeightsStore5[714];
			WeightsStore5[15] <= WeightsStore5[715];
			WeightsStore5[16] <= WeightsStore5[716];
			WeightsStore5[17] <= WeightsStore5[717];
			WeightsStore5[18] <= WeightsStore5[718];
			WeightsStore5[19] <= WeightsStore5[719];
			WeightsStore5[20] <= WeightsStore5[720];
			WeightsStore5[21] <= WeightsStore5[721];
			WeightsStore5[22] <= WeightsStore5[722];
			WeightsStore5[23] <= WeightsStore5[723];
			WeightsStore5[24] <= WeightsStore5[724];
			WeightsStore5[25] <= WeightsStore5[725];
			WeightsStore5[26] <= WeightsStore5[726];
			WeightsStore5[27] <= WeightsStore5[727];
			WeightsStore6[0] <= WeightsStore6[700];
			WeightsStore6[1] <= WeightsStore6[701];
			WeightsStore6[2] <= WeightsStore6[702];
			WeightsStore6[3] <= WeightsStore6[703];
			WeightsStore6[4] <= WeightsStore6[704];
			WeightsStore6[5] <= WeightsStore6[705];
			WeightsStore6[6] <= WeightsStore6[706];
			WeightsStore6[7] <= WeightsStore6[707];
			WeightsStore6[8] <= WeightsStore6[708];
			WeightsStore6[9] <= WeightsStore6[709];
			WeightsStore6[10] <= WeightsStore6[710];
			WeightsStore6[11] <= WeightsStore6[711];
			WeightsStore6[12] <= WeightsStore6[712];
			WeightsStore6[13] <= WeightsStore6[713];
			WeightsStore6[14] <= WeightsStore6[714];
			WeightsStore6[15] <= WeightsStore6[715];
			WeightsStore6[16] <= WeightsStore6[716];
			WeightsStore6[17] <= WeightsStore6[717];
			WeightsStore6[18] <= WeightsStore6[718];
			WeightsStore6[19] <= WeightsStore6[719];
			WeightsStore6[20] <= WeightsStore6[720];
			WeightsStore6[21] <= WeightsStore6[721];
			WeightsStore6[22] <= WeightsStore6[722];
			WeightsStore6[23] <= WeightsStore6[723];
			WeightsStore6[24] <= WeightsStore6[724];
			WeightsStore6[25] <= WeightsStore6[725];
			WeightsStore6[26] <= WeightsStore6[726];
			WeightsStore6[27] <= WeightsStore6[727];
			WeightsStore7[0] <= WeightsStore7[700];
			WeightsStore7[1] <= WeightsStore7[701];
			WeightsStore7[2] <= WeightsStore7[702];
			WeightsStore7[3] <= WeightsStore7[703];
			WeightsStore7[4] <= WeightsStore7[704];
			WeightsStore7[5] <= WeightsStore7[705];
			WeightsStore7[6] <= WeightsStore7[706];
			WeightsStore7[7] <= WeightsStore7[707];
			WeightsStore7[8] <= WeightsStore7[708];
			WeightsStore7[9] <= WeightsStore7[709];
			WeightsStore7[10] <= WeightsStore7[710];
			WeightsStore7[11] <= WeightsStore7[711];
			WeightsStore7[12] <= WeightsStore7[712];
			WeightsStore7[13] <= WeightsStore7[713];
			WeightsStore7[14] <= WeightsStore7[714];
			WeightsStore7[15] <= WeightsStore7[715];
			WeightsStore7[16] <= WeightsStore7[716];
			WeightsStore7[17] <= WeightsStore7[717];
			WeightsStore7[18] <= WeightsStore7[718];
			WeightsStore7[19] <= WeightsStore7[719];
			WeightsStore7[20] <= WeightsStore7[720];
			WeightsStore7[21] <= WeightsStore7[721];
			WeightsStore7[22] <= WeightsStore7[722];
			WeightsStore7[23] <= WeightsStore7[723];
			WeightsStore7[24] <= WeightsStore7[724];
			WeightsStore7[25] <= WeightsStore7[725];
			WeightsStore7[26] <= WeightsStore7[726];
			WeightsStore7[27] <= WeightsStore7[727];
			WeightsStore8[0] <= WeightsStore8[700];
			WeightsStore8[1] <= WeightsStore8[701];
			WeightsStore8[2] <= WeightsStore8[702];
			WeightsStore8[3] <= WeightsStore8[703];
			WeightsStore8[4] <= WeightsStore8[704];
			WeightsStore8[5] <= WeightsStore8[705];
			WeightsStore8[6] <= WeightsStore8[706];
			WeightsStore8[7] <= WeightsStore8[707];
			WeightsStore8[8] <= WeightsStore8[708];
			WeightsStore8[9] <= WeightsStore8[709];
			WeightsStore8[10] <= WeightsStore8[710];
			WeightsStore8[11] <= WeightsStore8[711];
			WeightsStore8[12] <= WeightsStore8[712];
			WeightsStore8[13] <= WeightsStore8[713];
			WeightsStore8[14] <= WeightsStore8[714];
			WeightsStore8[15] <= WeightsStore8[715];
			WeightsStore8[16] <= WeightsStore8[716];
			WeightsStore8[17] <= WeightsStore8[717];
			WeightsStore8[18] <= WeightsStore8[718];
			WeightsStore8[19] <= WeightsStore8[719];
			WeightsStore8[20] <= WeightsStore8[720];
			WeightsStore8[21] <= WeightsStore8[721];
			WeightsStore8[22] <= WeightsStore8[722];
			WeightsStore8[23] <= WeightsStore8[723];
			WeightsStore8[24] <= WeightsStore8[724];
			WeightsStore8[25] <= WeightsStore8[725];
			WeightsStore8[26] <= WeightsStore8[726];
			WeightsStore8[27] <= WeightsStore8[727];
			WeightsStore9[0] <= WeightsStore9[700];
			WeightsStore9[1] <= WeightsStore9[701];
			WeightsStore9[2] <= WeightsStore9[702];
			WeightsStore9[3] <= WeightsStore9[703];
			WeightsStore9[4] <= WeightsStore9[704];
			WeightsStore9[5] <= WeightsStore9[705];
			WeightsStore9[6] <= WeightsStore9[706];
			WeightsStore9[7] <= WeightsStore9[707];
			WeightsStore9[8] <= WeightsStore9[708];
			WeightsStore9[9] <= WeightsStore9[709];
			WeightsStore9[10] <= WeightsStore9[710];
			WeightsStore9[11] <= WeightsStore9[711];
			WeightsStore9[12] <= WeightsStore9[712];
			WeightsStore9[13] <= WeightsStore9[713];
			WeightsStore9[14] <= WeightsStore9[714];
			WeightsStore9[15] <= WeightsStore9[715];
			WeightsStore9[16] <= WeightsStore9[716];
			WeightsStore9[17] <= WeightsStore9[717];
			WeightsStore9[18] <= WeightsStore9[718];
			WeightsStore9[19] <= WeightsStore9[719];
			WeightsStore9[20] <= WeightsStore9[720];
			WeightsStore9[21] <= WeightsStore9[721];
			WeightsStore9[22] <= WeightsStore9[722];
			WeightsStore9[23] <= WeightsStore9[723];
			WeightsStore9[24] <= WeightsStore9[724];
			WeightsStore9[25] <= WeightsStore9[725];
			WeightsStore9[26] <= WeightsStore9[726];
			WeightsStore9[27] <= WeightsStore9[727];
		end else if(switchCounter == 32'd181)begin
			PixelsStore[0] <= PixelsStore[728];
			PixelsStore[1] <= PixelsStore[729];
			PixelsStore[2] <= PixelsStore[730];
			PixelsStore[3] <= PixelsStore[731];
			PixelsStore[4] <= PixelsStore[732];
			PixelsStore[5] <= PixelsStore[733];
			PixelsStore[6] <= PixelsStore[734];
			PixelsStore[7] <= PixelsStore[735];
			PixelsStore[8] <= PixelsStore[736];
			PixelsStore[9] <= PixelsStore[737];
			PixelsStore[10] <= PixelsStore[738];
			PixelsStore[11] <= PixelsStore[739];
			PixelsStore[12] <= PixelsStore[740];
			PixelsStore[13] <= PixelsStore[741];
			PixelsStore[14] <= PixelsStore[742];
			PixelsStore[15] <= PixelsStore[743];
			PixelsStore[16] <= PixelsStore[744];
			PixelsStore[17] <= PixelsStore[745];
			PixelsStore[18] <= PixelsStore[746];
			PixelsStore[19] <= PixelsStore[747];
			PixelsStore[20] <= PixelsStore[748];
			PixelsStore[21] <= PixelsStore[749];
			PixelsStore[22] <= PixelsStore[750];
			PixelsStore[23] <= PixelsStore[751];
			PixelsStore[24] <= PixelsStore[752];
			PixelsStore[25] <= PixelsStore[753];
			PixelsStore[26] <= PixelsStore[754];
			PixelsStore[27] <= PixelsStore[755];
			WeightsStore0[0] <= WeightsStore0[728];
			WeightsStore0[1] <= WeightsStore0[729];
			WeightsStore0[2] <= WeightsStore0[730];
			WeightsStore0[3] <= WeightsStore0[731];
			WeightsStore0[4] <= WeightsStore0[732];
			WeightsStore0[5] <= WeightsStore0[733];
			WeightsStore0[6] <= WeightsStore0[734];
			WeightsStore0[7] <= WeightsStore0[735];
			WeightsStore0[8] <= WeightsStore0[736];
			WeightsStore0[9] <= WeightsStore0[737];
			WeightsStore0[10] <= WeightsStore0[738];
			WeightsStore0[11] <= WeightsStore0[739];
			WeightsStore0[12] <= WeightsStore0[740];
			WeightsStore0[13] <= WeightsStore0[741];
			WeightsStore0[14] <= WeightsStore0[742];
			WeightsStore0[15] <= WeightsStore0[743];
			WeightsStore0[16] <= WeightsStore0[744];
			WeightsStore0[17] <= WeightsStore0[745];
			WeightsStore0[18] <= WeightsStore0[746];
			WeightsStore0[19] <= WeightsStore0[747];
			WeightsStore0[20] <= WeightsStore0[748];
			WeightsStore0[21] <= WeightsStore0[749];
			WeightsStore0[22] <= WeightsStore0[750];
			WeightsStore0[23] <= WeightsStore0[751];
			WeightsStore0[24] <= WeightsStore0[752];
			WeightsStore0[25] <= WeightsStore0[753];
			WeightsStore0[26] <= WeightsStore0[754];
			WeightsStore0[27] <= WeightsStore0[755];
			WeightsStore1[0] <= WeightsStore1[728];
			WeightsStore1[1] <= WeightsStore1[729];
			WeightsStore1[2] <= WeightsStore1[730];
			WeightsStore1[3] <= WeightsStore1[731];
			WeightsStore1[4] <= WeightsStore1[732];
			WeightsStore1[5] <= WeightsStore1[733];
			WeightsStore1[6] <= WeightsStore1[734];
			WeightsStore1[7] <= WeightsStore1[735];
			WeightsStore1[8] <= WeightsStore1[736];
			WeightsStore1[9] <= WeightsStore1[737];
			WeightsStore1[10] <= WeightsStore1[738];
			WeightsStore1[11] <= WeightsStore1[739];
			WeightsStore1[12] <= WeightsStore1[740];
			WeightsStore1[13] <= WeightsStore1[741];
			WeightsStore1[14] <= WeightsStore1[742];
			WeightsStore1[15] <= WeightsStore1[743];
			WeightsStore1[16] <= WeightsStore1[744];
			WeightsStore1[17] <= WeightsStore1[745];
			WeightsStore1[18] <= WeightsStore1[746];
			WeightsStore1[19] <= WeightsStore1[747];
			WeightsStore1[20] <= WeightsStore1[748];
			WeightsStore1[21] <= WeightsStore1[749];
			WeightsStore1[22] <= WeightsStore1[750];
			WeightsStore1[23] <= WeightsStore1[751];
			WeightsStore1[24] <= WeightsStore1[752];
			WeightsStore1[25] <= WeightsStore1[753];
			WeightsStore1[26] <= WeightsStore1[754];
			WeightsStore1[27] <= WeightsStore1[755];
			WeightsStore2[0] <= WeightsStore2[728];
			WeightsStore2[1] <= WeightsStore2[729];
			WeightsStore2[2] <= WeightsStore2[730];
			WeightsStore2[3] <= WeightsStore2[731];
			WeightsStore2[4] <= WeightsStore2[732];
			WeightsStore2[5] <= WeightsStore2[733];
			WeightsStore2[6] <= WeightsStore2[734];
			WeightsStore2[7] <= WeightsStore2[735];
			WeightsStore2[8] <= WeightsStore2[736];
			WeightsStore2[9] <= WeightsStore2[737];
			WeightsStore2[10] <= WeightsStore2[738];
			WeightsStore2[11] <= WeightsStore2[739];
			WeightsStore2[12] <= WeightsStore2[740];
			WeightsStore2[13] <= WeightsStore2[741];
			WeightsStore2[14] <= WeightsStore2[742];
			WeightsStore2[15] <= WeightsStore2[743];
			WeightsStore2[16] <= WeightsStore2[744];
			WeightsStore2[17] <= WeightsStore2[745];
			WeightsStore2[18] <= WeightsStore2[746];
			WeightsStore2[19] <= WeightsStore2[747];
			WeightsStore2[20] <= WeightsStore2[748];
			WeightsStore2[21] <= WeightsStore2[749];
			WeightsStore2[22] <= WeightsStore2[750];
			WeightsStore2[23] <= WeightsStore2[751];
			WeightsStore2[24] <= WeightsStore2[752];
			WeightsStore2[25] <= WeightsStore2[753];
			WeightsStore2[26] <= WeightsStore2[754];
			WeightsStore2[27] <= WeightsStore2[755];
			WeightsStore3[0] <= WeightsStore3[728];
			WeightsStore3[1] <= WeightsStore3[729];
			WeightsStore3[2] <= WeightsStore3[730];
			WeightsStore3[3] <= WeightsStore3[731];
			WeightsStore3[4] <= WeightsStore3[732];
			WeightsStore3[5] <= WeightsStore3[733];
			WeightsStore3[6] <= WeightsStore3[734];
			WeightsStore3[7] <= WeightsStore3[735];
			WeightsStore3[8] <= WeightsStore3[736];
			WeightsStore3[9] <= WeightsStore3[737];
			WeightsStore3[10] <= WeightsStore3[738];
			WeightsStore3[11] <= WeightsStore3[739];
			WeightsStore3[12] <= WeightsStore3[740];
			WeightsStore3[13] <= WeightsStore3[741];
			WeightsStore3[14] <= WeightsStore3[742];
			WeightsStore3[15] <= WeightsStore3[743];
			WeightsStore3[16] <= WeightsStore3[744];
			WeightsStore3[17] <= WeightsStore3[745];
			WeightsStore3[18] <= WeightsStore3[746];
			WeightsStore3[19] <= WeightsStore3[747];
			WeightsStore3[20] <= WeightsStore3[748];
			WeightsStore3[21] <= WeightsStore3[749];
			WeightsStore3[22] <= WeightsStore3[750];
			WeightsStore3[23] <= WeightsStore3[751];
			WeightsStore3[24] <= WeightsStore3[752];
			WeightsStore3[25] <= WeightsStore3[753];
			WeightsStore3[26] <= WeightsStore3[754];
			WeightsStore3[27] <= WeightsStore3[755];
			WeightsStore4[0] <= WeightsStore4[728];
			WeightsStore4[1] <= WeightsStore4[729];
			WeightsStore4[2] <= WeightsStore4[730];
			WeightsStore4[3] <= WeightsStore4[731];
			WeightsStore4[4] <= WeightsStore4[732];
			WeightsStore4[5] <= WeightsStore4[733];
			WeightsStore4[6] <= WeightsStore4[734];
			WeightsStore4[7] <= WeightsStore4[735];
			WeightsStore4[8] <= WeightsStore4[736];
			WeightsStore4[9] <= WeightsStore4[737];
			WeightsStore4[10] <= WeightsStore4[738];
			WeightsStore4[11] <= WeightsStore4[739];
			WeightsStore4[12] <= WeightsStore4[740];
			WeightsStore4[13] <= WeightsStore4[741];
			WeightsStore4[14] <= WeightsStore4[742];
			WeightsStore4[15] <= WeightsStore4[743];
			WeightsStore4[16] <= WeightsStore4[744];
			WeightsStore4[17] <= WeightsStore4[745];
			WeightsStore4[18] <= WeightsStore4[746];
			WeightsStore4[19] <= WeightsStore4[747];
			WeightsStore4[20] <= WeightsStore4[748];
			WeightsStore4[21] <= WeightsStore4[749];
			WeightsStore4[22] <= WeightsStore4[750];
			WeightsStore4[23] <= WeightsStore4[751];
			WeightsStore4[24] <= WeightsStore4[752];
			WeightsStore4[25] <= WeightsStore4[753];
			WeightsStore4[26] <= WeightsStore4[754];
			WeightsStore4[27] <= WeightsStore4[755];
			WeightsStore5[0] <= WeightsStore5[728];
			WeightsStore5[1] <= WeightsStore5[729];
			WeightsStore5[2] <= WeightsStore5[730];
			WeightsStore5[3] <= WeightsStore5[731];
			WeightsStore5[4] <= WeightsStore5[732];
			WeightsStore5[5] <= WeightsStore5[733];
			WeightsStore5[6] <= WeightsStore5[734];
			WeightsStore5[7] <= WeightsStore5[735];
			WeightsStore5[8] <= WeightsStore5[736];
			WeightsStore5[9] <= WeightsStore5[737];
			WeightsStore5[10] <= WeightsStore5[738];
			WeightsStore5[11] <= WeightsStore5[739];
			WeightsStore5[12] <= WeightsStore5[740];
			WeightsStore5[13] <= WeightsStore5[741];
			WeightsStore5[14] <= WeightsStore5[742];
			WeightsStore5[15] <= WeightsStore5[743];
			WeightsStore5[16] <= WeightsStore5[744];
			WeightsStore5[17] <= WeightsStore5[745];
			WeightsStore5[18] <= WeightsStore5[746];
			WeightsStore5[19] <= WeightsStore5[747];
			WeightsStore5[20] <= WeightsStore5[748];
			WeightsStore5[21] <= WeightsStore5[749];
			WeightsStore5[22] <= WeightsStore5[750];
			WeightsStore5[23] <= WeightsStore5[751];
			WeightsStore5[24] <= WeightsStore5[752];
			WeightsStore5[25] <= WeightsStore5[753];
			WeightsStore5[26] <= WeightsStore5[754];
			WeightsStore5[27] <= WeightsStore5[755];
			WeightsStore6[0] <= WeightsStore6[728];
			WeightsStore6[1] <= WeightsStore6[729];
			WeightsStore6[2] <= WeightsStore6[730];
			WeightsStore6[3] <= WeightsStore6[731];
			WeightsStore6[4] <= WeightsStore6[732];
			WeightsStore6[5] <= WeightsStore6[733];
			WeightsStore6[6] <= WeightsStore6[734];
			WeightsStore6[7] <= WeightsStore6[735];
			WeightsStore6[8] <= WeightsStore6[736];
			WeightsStore6[9] <= WeightsStore6[737];
			WeightsStore6[10] <= WeightsStore6[738];
			WeightsStore6[11] <= WeightsStore6[739];
			WeightsStore6[12] <= WeightsStore6[740];
			WeightsStore6[13] <= WeightsStore6[741];
			WeightsStore6[14] <= WeightsStore6[742];
			WeightsStore6[15] <= WeightsStore6[743];
			WeightsStore6[16] <= WeightsStore6[744];
			WeightsStore6[17] <= WeightsStore6[745];
			WeightsStore6[18] <= WeightsStore6[746];
			WeightsStore6[19] <= WeightsStore6[747];
			WeightsStore6[20] <= WeightsStore6[748];
			WeightsStore6[21] <= WeightsStore6[749];
			WeightsStore6[22] <= WeightsStore6[750];
			WeightsStore6[23] <= WeightsStore6[751];
			WeightsStore6[24] <= WeightsStore6[752];
			WeightsStore6[25] <= WeightsStore6[753];
			WeightsStore6[26] <= WeightsStore6[754];
			WeightsStore6[27] <= WeightsStore6[755];
			WeightsStore7[0] <= WeightsStore7[728];
			WeightsStore7[1] <= WeightsStore7[729];
			WeightsStore7[2] <= WeightsStore7[730];
			WeightsStore7[3] <= WeightsStore7[731];
			WeightsStore7[4] <= WeightsStore7[732];
			WeightsStore7[5] <= WeightsStore7[733];
			WeightsStore7[6] <= WeightsStore7[734];
			WeightsStore7[7] <= WeightsStore7[735];
			WeightsStore7[8] <= WeightsStore7[736];
			WeightsStore7[9] <= WeightsStore7[737];
			WeightsStore7[10] <= WeightsStore7[738];
			WeightsStore7[11] <= WeightsStore7[739];
			WeightsStore7[12] <= WeightsStore7[740];
			WeightsStore7[13] <= WeightsStore7[741];
			WeightsStore7[14] <= WeightsStore7[742];
			WeightsStore7[15] <= WeightsStore7[743];
			WeightsStore7[16] <= WeightsStore7[744];
			WeightsStore7[17] <= WeightsStore7[745];
			WeightsStore7[18] <= WeightsStore7[746];
			WeightsStore7[19] <= WeightsStore7[747];
			WeightsStore7[20] <= WeightsStore7[748];
			WeightsStore7[21] <= WeightsStore7[749];
			WeightsStore7[22] <= WeightsStore7[750];
			WeightsStore7[23] <= WeightsStore7[751];
			WeightsStore7[24] <= WeightsStore7[752];
			WeightsStore7[25] <= WeightsStore7[753];
			WeightsStore7[26] <= WeightsStore7[754];
			WeightsStore7[27] <= WeightsStore7[755];
			WeightsStore8[0] <= WeightsStore8[728];
			WeightsStore8[1] <= WeightsStore8[729];
			WeightsStore8[2] <= WeightsStore8[730];
			WeightsStore8[3] <= WeightsStore8[731];
			WeightsStore8[4] <= WeightsStore8[732];
			WeightsStore8[5] <= WeightsStore8[733];
			WeightsStore8[6] <= WeightsStore8[734];
			WeightsStore8[7] <= WeightsStore8[735];
			WeightsStore8[8] <= WeightsStore8[736];
			WeightsStore8[9] <= WeightsStore8[737];
			WeightsStore8[10] <= WeightsStore8[738];
			WeightsStore8[11] <= WeightsStore8[739];
			WeightsStore8[12] <= WeightsStore8[740];
			WeightsStore8[13] <= WeightsStore8[741];
			WeightsStore8[14] <= WeightsStore8[742];
			WeightsStore8[15] <= WeightsStore8[743];
			WeightsStore8[16] <= WeightsStore8[744];
			WeightsStore8[17] <= WeightsStore8[745];
			WeightsStore8[18] <= WeightsStore8[746];
			WeightsStore8[19] <= WeightsStore8[747];
			WeightsStore8[20] <= WeightsStore8[748];
			WeightsStore8[21] <= WeightsStore8[749];
			WeightsStore8[22] <= WeightsStore8[750];
			WeightsStore8[23] <= WeightsStore8[751];
			WeightsStore8[24] <= WeightsStore8[752];
			WeightsStore8[25] <= WeightsStore8[753];
			WeightsStore8[26] <= WeightsStore8[754];
			WeightsStore8[27] <= WeightsStore8[755];
			WeightsStore9[0] <= WeightsStore9[728];
			WeightsStore9[1] <= WeightsStore9[729];
			WeightsStore9[2] <= WeightsStore9[730];
			WeightsStore9[3] <= WeightsStore9[731];
			WeightsStore9[4] <= WeightsStore9[732];
			WeightsStore9[5] <= WeightsStore9[733];
			WeightsStore9[6] <= WeightsStore9[734];
			WeightsStore9[7] <= WeightsStore9[735];
			WeightsStore9[8] <= WeightsStore9[736];
			WeightsStore9[9] <= WeightsStore9[737];
			WeightsStore9[10] <= WeightsStore9[738];
			WeightsStore9[11] <= WeightsStore9[739];
			WeightsStore9[12] <= WeightsStore9[740];
			WeightsStore9[13] <= WeightsStore9[741];
			WeightsStore9[14] <= WeightsStore9[742];
			WeightsStore9[15] <= WeightsStore9[743];
			WeightsStore9[16] <= WeightsStore9[744];
			WeightsStore9[17] <= WeightsStore9[745];
			WeightsStore9[18] <= WeightsStore9[746];
			WeightsStore9[19] <= WeightsStore9[747];
			WeightsStore9[20] <= WeightsStore9[748];
			WeightsStore9[21] <= WeightsStore9[749];
			WeightsStore9[22] <= WeightsStore9[750];
			WeightsStore9[23] <= WeightsStore9[751];
			WeightsStore9[24] <= WeightsStore9[752];
			WeightsStore9[25] <= WeightsStore9[753];
			WeightsStore9[26] <= WeightsStore9[754];
			WeightsStore9[27] <= WeightsStore9[755];
		end else if(switchCounter == 32'd188)begin
			PixelsStore[0] <= PixelsStore[756];
			PixelsStore[1] <= PixelsStore[757];
			PixelsStore[2] <= PixelsStore[758];
			PixelsStore[3] <= PixelsStore[759];
			PixelsStore[4] <= PixelsStore[760];
			PixelsStore[5] <= PixelsStore[761];
			PixelsStore[6] <= PixelsStore[762];
			PixelsStore[7] <= PixelsStore[763];
			PixelsStore[8] <= PixelsStore[764];
			PixelsStore[9] <= PixelsStore[765];
			PixelsStore[10] <= PixelsStore[766];
			PixelsStore[11] <= PixelsStore[767];
			PixelsStore[12] <= PixelsStore[768];
			PixelsStore[13] <= PixelsStore[769];
			PixelsStore[14] <= PixelsStore[770];
			PixelsStore[15] <= PixelsStore[771];
			PixelsStore[16] <= PixelsStore[772];
			PixelsStore[17] <= PixelsStore[773];
			PixelsStore[18] <= PixelsStore[774];
			PixelsStore[19] <= PixelsStore[775];
			PixelsStore[20] <= PixelsStore[776];
			PixelsStore[21] <= PixelsStore[777];
			PixelsStore[22] <= PixelsStore[778];
			PixelsStore[23] <= PixelsStore[779];
			PixelsStore[24] <= PixelsStore[780];
			PixelsStore[25] <= PixelsStore[781];
			PixelsStore[26] <= PixelsStore[782];
			PixelsStore[27] <= PixelsStore[783];
			WeightsStore0[0] <= WeightsStore0[756];
			WeightsStore0[1] <= WeightsStore0[757];
			WeightsStore0[2] <= WeightsStore0[758];
			WeightsStore0[3] <= WeightsStore0[759];
			WeightsStore0[4] <= WeightsStore0[760];
			WeightsStore0[5] <= WeightsStore0[761];
			WeightsStore0[6] <= WeightsStore0[762];
			WeightsStore0[7] <= WeightsStore0[763];
			WeightsStore0[8] <= WeightsStore0[764];
			WeightsStore0[9] <= WeightsStore0[765];
			WeightsStore0[10] <= WeightsStore0[766];
			WeightsStore0[11] <= WeightsStore0[767];
			WeightsStore0[12] <= WeightsStore0[768];
			WeightsStore0[13] <= WeightsStore0[769];
			WeightsStore0[14] <= WeightsStore0[770];
			WeightsStore0[15] <= WeightsStore0[771];
			WeightsStore0[16] <= WeightsStore0[772];
			WeightsStore0[17] <= WeightsStore0[773];
			WeightsStore0[18] <= WeightsStore0[774];
			WeightsStore0[19] <= WeightsStore0[775];
			WeightsStore0[20] <= WeightsStore0[776];
			WeightsStore0[21] <= WeightsStore0[777];
			WeightsStore0[22] <= WeightsStore0[778];
			WeightsStore0[23] <= WeightsStore0[779];
			WeightsStore0[24] <= WeightsStore0[780];
			WeightsStore0[25] <= WeightsStore0[781];
			WeightsStore0[26] <= WeightsStore0[782];
			WeightsStore0[27] <= WeightsStore0[783];
			WeightsStore1[0] <= WeightsStore1[756];
			WeightsStore1[1] <= WeightsStore1[757];
			WeightsStore1[2] <= WeightsStore1[758];
			WeightsStore1[3] <= WeightsStore1[759];
			WeightsStore1[4] <= WeightsStore1[760];
			WeightsStore1[5] <= WeightsStore1[761];
			WeightsStore1[6] <= WeightsStore1[762];
			WeightsStore1[7] <= WeightsStore1[763];
			WeightsStore1[8] <= WeightsStore1[764];
			WeightsStore1[9] <= WeightsStore1[765];
			WeightsStore1[10] <= WeightsStore1[766];
			WeightsStore1[11] <= WeightsStore1[767];
			WeightsStore1[12] <= WeightsStore1[768];
			WeightsStore1[13] <= WeightsStore1[769];
			WeightsStore1[14] <= WeightsStore1[770];
			WeightsStore1[15] <= WeightsStore1[771];
			WeightsStore1[16] <= WeightsStore1[772];
			WeightsStore1[17] <= WeightsStore1[773];
			WeightsStore1[18] <= WeightsStore1[774];
			WeightsStore1[19] <= WeightsStore1[775];
			WeightsStore1[20] <= WeightsStore1[776];
			WeightsStore1[21] <= WeightsStore1[777];
			WeightsStore1[22] <= WeightsStore1[778];
			WeightsStore1[23] <= WeightsStore1[779];
			WeightsStore1[24] <= WeightsStore1[780];
			WeightsStore1[25] <= WeightsStore1[781];
			WeightsStore1[26] <= WeightsStore1[782];
			WeightsStore1[27] <= WeightsStore1[783];
			WeightsStore2[0] <= WeightsStore2[756];
			WeightsStore2[1] <= WeightsStore2[757];
			WeightsStore2[2] <= WeightsStore2[758];
			WeightsStore2[3] <= WeightsStore2[759];
			WeightsStore2[4] <= WeightsStore2[760];
			WeightsStore2[5] <= WeightsStore2[761];
			WeightsStore2[6] <= WeightsStore2[762];
			WeightsStore2[7] <= WeightsStore2[763];
			WeightsStore2[8] <= WeightsStore2[764];
			WeightsStore2[9] <= WeightsStore2[765];
			WeightsStore2[10] <= WeightsStore2[766];
			WeightsStore2[11] <= WeightsStore2[767];
			WeightsStore2[12] <= WeightsStore2[768];
			WeightsStore2[13] <= WeightsStore2[769];
			WeightsStore2[14] <= WeightsStore2[770];
			WeightsStore2[15] <= WeightsStore2[771];
			WeightsStore2[16] <= WeightsStore2[772];
			WeightsStore2[17] <= WeightsStore2[773];
			WeightsStore2[18] <= WeightsStore2[774];
			WeightsStore2[19] <= WeightsStore2[775];
			WeightsStore2[20] <= WeightsStore2[776];
			WeightsStore2[21] <= WeightsStore2[777];
			WeightsStore2[22] <= WeightsStore2[778];
			WeightsStore2[23] <= WeightsStore2[779];
			WeightsStore2[24] <= WeightsStore2[780];
			WeightsStore2[25] <= WeightsStore2[781];
			WeightsStore2[26] <= WeightsStore2[782];
			WeightsStore2[27] <= WeightsStore2[783];
			WeightsStore3[0] <= WeightsStore3[756];
			WeightsStore3[1] <= WeightsStore3[757];
			WeightsStore3[2] <= WeightsStore3[758];
			WeightsStore3[3] <= WeightsStore3[759];
			WeightsStore3[4] <= WeightsStore3[760];
			WeightsStore3[5] <= WeightsStore3[761];
			WeightsStore3[6] <= WeightsStore3[762];
			WeightsStore3[7] <= WeightsStore3[763];
			WeightsStore3[8] <= WeightsStore3[764];
			WeightsStore3[9] <= WeightsStore3[765];
			WeightsStore3[10] <= WeightsStore3[766];
			WeightsStore3[11] <= WeightsStore3[767];
			WeightsStore3[12] <= WeightsStore3[768];
			WeightsStore3[13] <= WeightsStore3[769];
			WeightsStore3[14] <= WeightsStore3[770];
			WeightsStore3[15] <= WeightsStore3[771];
			WeightsStore3[16] <= WeightsStore3[772];
			WeightsStore3[17] <= WeightsStore3[773];
			WeightsStore3[18] <= WeightsStore3[774];
			WeightsStore3[19] <= WeightsStore3[775];
			WeightsStore3[20] <= WeightsStore3[776];
			WeightsStore3[21] <= WeightsStore3[777];
			WeightsStore3[22] <= WeightsStore3[778];
			WeightsStore3[23] <= WeightsStore3[779];
			WeightsStore3[24] <= WeightsStore3[780];
			WeightsStore3[25] <= WeightsStore3[781];
			WeightsStore3[26] <= WeightsStore3[782];
			WeightsStore3[27] <= WeightsStore3[783];
			WeightsStore4[0] <= WeightsStore4[756];
			WeightsStore4[1] <= WeightsStore4[757];
			WeightsStore4[2] <= WeightsStore4[758];
			WeightsStore4[3] <= WeightsStore4[759];
			WeightsStore4[4] <= WeightsStore4[760];
			WeightsStore4[5] <= WeightsStore4[761];
			WeightsStore4[6] <= WeightsStore4[762];
			WeightsStore4[7] <= WeightsStore4[763];
			WeightsStore4[8] <= WeightsStore4[764];
			WeightsStore4[9] <= WeightsStore4[765];
			WeightsStore4[10] <= WeightsStore4[766];
			WeightsStore4[11] <= WeightsStore4[767];
			WeightsStore4[12] <= WeightsStore4[768];
			WeightsStore4[13] <= WeightsStore4[769];
			WeightsStore4[14] <= WeightsStore4[770];
			WeightsStore4[15] <= WeightsStore4[771];
			WeightsStore4[16] <= WeightsStore4[772];
			WeightsStore4[17] <= WeightsStore4[773];
			WeightsStore4[18] <= WeightsStore4[774];
			WeightsStore4[19] <= WeightsStore4[775];
			WeightsStore4[20] <= WeightsStore4[776];
			WeightsStore4[21] <= WeightsStore4[777];
			WeightsStore4[22] <= WeightsStore4[778];
			WeightsStore4[23] <= WeightsStore4[779];
			WeightsStore4[24] <= WeightsStore4[780];
			WeightsStore4[25] <= WeightsStore4[781];
			WeightsStore4[26] <= WeightsStore4[782];
			WeightsStore4[27] <= WeightsStore4[783];
			WeightsStore5[0] <= WeightsStore5[756];
			WeightsStore5[1] <= WeightsStore5[757];
			WeightsStore5[2] <= WeightsStore5[758];
			WeightsStore5[3] <= WeightsStore5[759];
			WeightsStore5[4] <= WeightsStore5[760];
			WeightsStore5[5] <= WeightsStore5[761];
			WeightsStore5[6] <= WeightsStore5[762];
			WeightsStore5[7] <= WeightsStore5[763];
			WeightsStore5[8] <= WeightsStore5[764];
			WeightsStore5[9] <= WeightsStore5[765];
			WeightsStore5[10] <= WeightsStore5[766];
			WeightsStore5[11] <= WeightsStore5[767];
			WeightsStore5[12] <= WeightsStore5[768];
			WeightsStore5[13] <= WeightsStore5[769];
			WeightsStore5[14] <= WeightsStore5[770];
			WeightsStore5[15] <= WeightsStore5[771];
			WeightsStore5[16] <= WeightsStore5[772];
			WeightsStore5[17] <= WeightsStore5[773];
			WeightsStore5[18] <= WeightsStore5[774];
			WeightsStore5[19] <= WeightsStore5[775];
			WeightsStore5[20] <= WeightsStore5[776];
			WeightsStore5[21] <= WeightsStore5[777];
			WeightsStore5[22] <= WeightsStore5[778];
			WeightsStore5[23] <= WeightsStore5[779];
			WeightsStore5[24] <= WeightsStore5[780];
			WeightsStore5[25] <= WeightsStore5[781];
			WeightsStore5[26] <= WeightsStore5[782];
			WeightsStore5[27] <= WeightsStore5[783];
			WeightsStore6[0] <= WeightsStore6[756];
			WeightsStore6[1] <= WeightsStore6[757];
			WeightsStore6[2] <= WeightsStore6[758];
			WeightsStore6[3] <= WeightsStore6[759];
			WeightsStore6[4] <= WeightsStore6[760];
			WeightsStore6[5] <= WeightsStore6[761];
			WeightsStore6[6] <= WeightsStore6[762];
			WeightsStore6[7] <= WeightsStore6[763];
			WeightsStore6[8] <= WeightsStore6[764];
			WeightsStore6[9] <= WeightsStore6[765];
			WeightsStore6[10] <= WeightsStore6[766];
			WeightsStore6[11] <= WeightsStore6[767];
			WeightsStore6[12] <= WeightsStore6[768];
			WeightsStore6[13] <= WeightsStore6[769];
			WeightsStore6[14] <= WeightsStore6[770];
			WeightsStore6[15] <= WeightsStore6[771];
			WeightsStore6[16] <= WeightsStore6[772];
			WeightsStore6[17] <= WeightsStore6[773];
			WeightsStore6[18] <= WeightsStore6[774];
			WeightsStore6[19] <= WeightsStore6[775];
			WeightsStore6[20] <= WeightsStore6[776];
			WeightsStore6[21] <= WeightsStore6[777];
			WeightsStore6[22] <= WeightsStore6[778];
			WeightsStore6[23] <= WeightsStore6[779];
			WeightsStore6[24] <= WeightsStore6[780];
			WeightsStore6[25] <= WeightsStore6[781];
			WeightsStore6[26] <= WeightsStore6[782];
			WeightsStore6[27] <= WeightsStore6[783];
			WeightsStore7[0] <= WeightsStore7[756];
			WeightsStore7[1] <= WeightsStore7[757];
			WeightsStore7[2] <= WeightsStore7[758];
			WeightsStore7[3] <= WeightsStore7[759];
			WeightsStore7[4] <= WeightsStore7[760];
			WeightsStore7[5] <= WeightsStore7[761];
			WeightsStore7[6] <= WeightsStore7[762];
			WeightsStore7[7] <= WeightsStore7[763];
			WeightsStore7[8] <= WeightsStore7[764];
			WeightsStore7[9] <= WeightsStore7[765];
			WeightsStore7[10] <= WeightsStore7[766];
			WeightsStore7[11] <= WeightsStore7[767];
			WeightsStore7[12] <= WeightsStore7[768];
			WeightsStore7[13] <= WeightsStore7[769];
			WeightsStore7[14] <= WeightsStore7[770];
			WeightsStore7[15] <= WeightsStore7[771];
			WeightsStore7[16] <= WeightsStore7[772];
			WeightsStore7[17] <= WeightsStore7[773];
			WeightsStore7[18] <= WeightsStore7[774];
			WeightsStore7[19] <= WeightsStore7[775];
			WeightsStore7[20] <= WeightsStore7[776];
			WeightsStore7[21] <= WeightsStore7[777];
			WeightsStore7[22] <= WeightsStore7[778];
			WeightsStore7[23] <= WeightsStore7[779];
			WeightsStore7[24] <= WeightsStore7[780];
			WeightsStore7[25] <= WeightsStore7[781];
			WeightsStore7[26] <= WeightsStore7[782];
			WeightsStore7[27] <= WeightsStore7[783];
			WeightsStore8[0] <= WeightsStore8[756];
			WeightsStore8[1] <= WeightsStore8[757];
			WeightsStore8[2] <= WeightsStore8[758];
			WeightsStore8[3] <= WeightsStore8[759];
			WeightsStore8[4] <= WeightsStore8[760];
			WeightsStore8[5] <= WeightsStore8[761];
			WeightsStore8[6] <= WeightsStore8[762];
			WeightsStore8[7] <= WeightsStore8[763];
			WeightsStore8[8] <= WeightsStore8[764];
			WeightsStore8[9] <= WeightsStore8[765];
			WeightsStore8[10] <= WeightsStore8[766];
			WeightsStore8[11] <= WeightsStore8[767];
			WeightsStore8[12] <= WeightsStore8[768];
			WeightsStore8[13] <= WeightsStore8[769];
			WeightsStore8[14] <= WeightsStore8[770];
			WeightsStore8[15] <= WeightsStore8[771];
			WeightsStore8[16] <= WeightsStore8[772];
			WeightsStore8[17] <= WeightsStore8[773];
			WeightsStore8[18] <= WeightsStore8[774];
			WeightsStore8[19] <= WeightsStore8[775];
			WeightsStore8[20] <= WeightsStore8[776];
			WeightsStore8[21] <= WeightsStore8[777];
			WeightsStore8[22] <= WeightsStore8[778];
			WeightsStore8[23] <= WeightsStore8[779];
			WeightsStore8[24] <= WeightsStore8[780];
			WeightsStore8[25] <= WeightsStore8[781];
			WeightsStore8[26] <= WeightsStore8[782];
			WeightsStore8[27] <= WeightsStore8[783];
			WeightsStore9[0] <= WeightsStore9[756];
			WeightsStore9[1] <= WeightsStore9[757];
			WeightsStore9[2] <= WeightsStore9[758];
			WeightsStore9[3] <= WeightsStore9[759];
			WeightsStore9[4] <= WeightsStore9[760];
			WeightsStore9[5] <= WeightsStore9[761];
			WeightsStore9[6] <= WeightsStore9[762];
			WeightsStore9[7] <= WeightsStore9[763];
			WeightsStore9[8] <= WeightsStore9[764];
			WeightsStore9[9] <= WeightsStore9[765];
			WeightsStore9[10] <= WeightsStore9[766];
			WeightsStore9[11] <= WeightsStore9[767];
			WeightsStore9[12] <= WeightsStore9[768];
			WeightsStore9[13] <= WeightsStore9[769];
			WeightsStore9[14] <= WeightsStore9[770];
			WeightsStore9[15] <= WeightsStore9[771];
			WeightsStore9[16] <= WeightsStore9[772];
			WeightsStore9[17] <= WeightsStore9[773];
			WeightsStore9[18] <= WeightsStore9[774];
			WeightsStore9[19] <= WeightsStore9[775];
			WeightsStore9[20] <= WeightsStore9[776];
			WeightsStore9[21] <= WeightsStore9[777];
			WeightsStore9[22] <= WeightsStore9[778];
			WeightsStore9[23] <= WeightsStore9[779];
			WeightsStore9[24] <= WeightsStore9[780];
			WeightsStore9[25] <= WeightsStore9[781];
			WeightsStore9[26] <= WeightsStore9[782];
			WeightsStore9[27] <= WeightsStore9[783];
		end else if(switchCounter == 32'd299) begin
			ready <= 1'b1;
			$display("%d %b.%b", switchCounter, value[259:252],value[251:234]);
			$display("%d %b.%b", switchCounter, value[233:226],value[225:208]);
			$display("%d %b.%b", switchCounter, value[207:200],value[199:182]);
			$display("%d %b.%b", switchCounter, value[181:174],value[173:156]);
			$display("%d %b.%b", switchCounter, value[155:148],value[147:130]);
			$display("%d %b.%b", switchCounter, value[129:122],value[121:104]);
			$display("%d %b.%b", switchCounter, value[103:96],value[95:78]);
			$display("%d %b.%b", switchCounter, value[77:70],value[69:52]);
			$display("%d %b.%b", switchCounter, value[51:44],value[43:26]);
			$display("%d %b.%b", switchCounter, value[25:18],value[17:0]);
		end
	end
end
endmodule
