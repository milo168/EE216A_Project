module test
#(parameter PIXEL_N = 784,
parameter WEIGHT_SIZE = 19,
parameter PIXEL_SIZE = 10)
(
input clk,
input GlobalReset,
input [PIXEL_N*PIXEL_SIZE-1:0] Pixels,
input [PIXEL_N*WEIGHT_SIZE-1:0] Weights,
output [25:0] value
);

wire[18:0] A [0:783];
wire[9:0] B [0:783];
reg[18:0] A1;
reg[18:0] A2;
reg[9:0] B1;
reg[9:0] B2;
wire[25:0] FPMAns1;
wire[25:0] FPMAns2;
wire[25:0] FPAAns;
reg[25:0] addAns [0:391];
reg[25:0] addInput [0:1];
reg[31:0] switchCounter = 32'd0;
assign value = addAns[0];

assign A[0] = Weights[18:0];
assign A[1] = Weights[37:19];
assign A[2] = Weights[56:38];
assign A[3] = Weights[75:57];
assign A[4] = Weights[94:76];
assign A[5] = Weights[113:95];
assign A[6] = Weights[132:114];
assign A[7] = Weights[151:133];
assign A[8] = Weights[170:152];
assign A[9] = Weights[189:171];
assign A[10] = Weights[208:190];
assign A[11] = Weights[227:209];
assign A[12] = Weights[246:228];
assign A[13] = Weights[265:247];
assign A[14] = Weights[284:266];
assign A[15] = Weights[303:285];
assign A[16] = Weights[322:304];
assign A[17] = Weights[341:323];
assign A[18] = Weights[360:342];
assign A[19] = Weights[379:361];
assign A[20] = Weights[398:380];
assign A[21] = Weights[417:399];
assign A[22] = Weights[436:418];
assign A[23] = Weights[455:437];
assign A[24] = Weights[474:456];
assign A[25] = Weights[493:475];
assign A[26] = Weights[512:494];
assign A[27] = Weights[531:513];
assign A[28] = Weights[550:532];
assign A[29] = Weights[569:551];
assign A[30] = Weights[588:570];
assign A[31] = Weights[607:589];
assign A[32] = Weights[626:608];
assign A[33] = Weights[645:627];
assign A[34] = Weights[664:646];
assign A[35] = Weights[683:665];
assign A[36] = Weights[702:684];
assign A[37] = Weights[721:703];
assign A[38] = Weights[740:722];
assign A[39] = Weights[759:741];
assign A[40] = Weights[778:760];
assign A[41] = Weights[797:779];
assign A[42] = Weights[816:798];
assign A[43] = Weights[835:817];
assign A[44] = Weights[854:836];
assign A[45] = Weights[873:855];
assign A[46] = Weights[892:874];
assign A[47] = Weights[911:893];
assign A[48] = Weights[930:912];
assign A[49] = Weights[949:931];
assign A[50] = Weights[968:950];
assign A[51] = Weights[987:969];
assign A[52] = Weights[1006:988];
assign A[53] = Weights[1025:1007];
assign A[54] = Weights[1044:1026];
assign A[55] = Weights[1063:1045];
assign A[56] = Weights[1082:1064];
assign A[57] = Weights[1101:1083];
assign A[58] = Weights[1120:1102];
assign A[59] = Weights[1139:1121];
assign A[60] = Weights[1158:1140];
assign A[61] = Weights[1177:1159];
assign A[62] = Weights[1196:1178];
assign A[63] = Weights[1215:1197];
assign A[64] = Weights[1234:1216];
assign A[65] = Weights[1253:1235];
assign A[66] = Weights[1272:1254];
assign A[67] = Weights[1291:1273];
assign A[68] = Weights[1310:1292];
assign A[69] = Weights[1329:1311];
assign A[70] = Weights[1348:1330];
assign A[71] = Weights[1367:1349];
assign A[72] = Weights[1386:1368];
assign A[73] = Weights[1405:1387];
assign A[74] = Weights[1424:1406];
assign A[75] = Weights[1443:1425];
assign A[76] = Weights[1462:1444];
assign A[77] = Weights[1481:1463];
assign A[78] = Weights[1500:1482];
assign A[79] = Weights[1519:1501];
assign A[80] = Weights[1538:1520];
assign A[81] = Weights[1557:1539];
assign A[82] = Weights[1576:1558];
assign A[83] = Weights[1595:1577];
assign A[84] = Weights[1614:1596];
assign A[85] = Weights[1633:1615];
assign A[86] = Weights[1652:1634];
assign A[87] = Weights[1671:1653];
assign A[88] = Weights[1690:1672];
assign A[89] = Weights[1709:1691];
assign A[90] = Weights[1728:1710];
assign A[91] = Weights[1747:1729];
assign A[92] = Weights[1766:1748];
assign A[93] = Weights[1785:1767];
assign A[94] = Weights[1804:1786];
assign A[95] = Weights[1823:1805];
assign A[96] = Weights[1842:1824];
assign A[97] = Weights[1861:1843];
assign A[98] = Weights[1880:1862];
assign A[99] = Weights[1899:1881];
assign A[100] = Weights[1918:1900];
assign A[101] = Weights[1937:1919];
assign A[102] = Weights[1956:1938];
assign A[103] = Weights[1975:1957];
assign A[104] = Weights[1994:1976];
assign A[105] = Weights[2013:1995];
assign A[106] = Weights[2032:2014];
assign A[107] = Weights[2051:2033];
assign A[108] = Weights[2070:2052];
assign A[109] = Weights[2089:2071];
assign A[110] = Weights[2108:2090];
assign A[111] = Weights[2127:2109];
assign A[112] = Weights[2146:2128];
assign A[113] = Weights[2165:2147];
assign A[114] = Weights[2184:2166];
assign A[115] = Weights[2203:2185];
assign A[116] = Weights[2222:2204];
assign A[117] = Weights[2241:2223];
assign A[118] = Weights[2260:2242];
assign A[119] = Weights[2279:2261];
assign A[120] = Weights[2298:2280];
assign A[121] = Weights[2317:2299];
assign A[122] = Weights[2336:2318];
assign A[123] = Weights[2355:2337];
assign A[124] = Weights[2374:2356];
assign A[125] = Weights[2393:2375];
assign A[126] = Weights[2412:2394];
assign A[127] = Weights[2431:2413];
assign A[128] = Weights[2450:2432];
assign A[129] = Weights[2469:2451];
assign A[130] = Weights[2488:2470];
assign A[131] = Weights[2507:2489];
assign A[132] = Weights[2526:2508];
assign A[133] = Weights[2545:2527];
assign A[134] = Weights[2564:2546];
assign A[135] = Weights[2583:2565];
assign A[136] = Weights[2602:2584];
assign A[137] = Weights[2621:2603];
assign A[138] = Weights[2640:2622];
assign A[139] = Weights[2659:2641];
assign A[140] = Weights[2678:2660];
assign A[141] = Weights[2697:2679];
assign A[142] = Weights[2716:2698];
assign A[143] = Weights[2735:2717];
assign A[144] = Weights[2754:2736];
assign A[145] = Weights[2773:2755];
assign A[146] = Weights[2792:2774];
assign A[147] = Weights[2811:2793];
assign A[148] = Weights[2830:2812];
assign A[149] = Weights[2849:2831];
assign A[150] = Weights[2868:2850];
assign A[151] = Weights[2887:2869];
assign A[152] = Weights[2906:2888];
assign A[153] = Weights[2925:2907];
assign A[154] = Weights[2944:2926];
assign A[155] = Weights[2963:2945];
assign A[156] = Weights[2982:2964];
assign A[157] = Weights[3001:2983];
assign A[158] = Weights[3020:3002];
assign A[159] = Weights[3039:3021];
assign A[160] = Weights[3058:3040];
assign A[161] = Weights[3077:3059];
assign A[162] = Weights[3096:3078];
assign A[163] = Weights[3115:3097];
assign A[164] = Weights[3134:3116];
assign A[165] = Weights[3153:3135];
assign A[166] = Weights[3172:3154];
assign A[167] = Weights[3191:3173];
assign A[168] = Weights[3210:3192];
assign A[169] = Weights[3229:3211];
assign A[170] = Weights[3248:3230];
assign A[171] = Weights[3267:3249];
assign A[172] = Weights[3286:3268];
assign A[173] = Weights[3305:3287];
assign A[174] = Weights[3324:3306];
assign A[175] = Weights[3343:3325];
assign A[176] = Weights[3362:3344];
assign A[177] = Weights[3381:3363];
assign A[178] = Weights[3400:3382];
assign A[179] = Weights[3419:3401];
assign A[180] = Weights[3438:3420];
assign A[181] = Weights[3457:3439];
assign A[182] = Weights[3476:3458];
assign A[183] = Weights[3495:3477];
assign A[184] = Weights[3514:3496];
assign A[185] = Weights[3533:3515];
assign A[186] = Weights[3552:3534];
assign A[187] = Weights[3571:3553];
assign A[188] = Weights[3590:3572];
assign A[189] = Weights[3609:3591];
assign A[190] = Weights[3628:3610];
assign A[191] = Weights[3647:3629];
assign A[192] = Weights[3666:3648];
assign A[193] = Weights[3685:3667];
assign A[194] = Weights[3704:3686];
assign A[195] = Weights[3723:3705];
assign A[196] = Weights[3742:3724];
assign A[197] = Weights[3761:3743];
assign A[198] = Weights[3780:3762];
assign A[199] = Weights[3799:3781];
assign A[200] = Weights[3818:3800];
assign A[201] = Weights[3837:3819];
assign A[202] = Weights[3856:3838];
assign A[203] = Weights[3875:3857];
assign A[204] = Weights[3894:3876];
assign A[205] = Weights[3913:3895];
assign A[206] = Weights[3932:3914];
assign A[207] = Weights[3951:3933];
assign A[208] = Weights[3970:3952];
assign A[209] = Weights[3989:3971];
assign A[210] = Weights[4008:3990];
assign A[211] = Weights[4027:4009];
assign A[212] = Weights[4046:4028];
assign A[213] = Weights[4065:4047];
assign A[214] = Weights[4084:4066];
assign A[215] = Weights[4103:4085];
assign A[216] = Weights[4122:4104];
assign A[217] = Weights[4141:4123];
assign A[218] = Weights[4160:4142];
assign A[219] = Weights[4179:4161];
assign A[220] = Weights[4198:4180];
assign A[221] = Weights[4217:4199];
assign A[222] = Weights[4236:4218];
assign A[223] = Weights[4255:4237];
assign A[224] = Weights[4274:4256];
assign A[225] = Weights[4293:4275];
assign A[226] = Weights[4312:4294];
assign A[227] = Weights[4331:4313];
assign A[228] = Weights[4350:4332];
assign A[229] = Weights[4369:4351];
assign A[230] = Weights[4388:4370];
assign A[231] = Weights[4407:4389];
assign A[232] = Weights[4426:4408];
assign A[233] = Weights[4445:4427];
assign A[234] = Weights[4464:4446];
assign A[235] = Weights[4483:4465];
assign A[236] = Weights[4502:4484];
assign A[237] = Weights[4521:4503];
assign A[238] = Weights[4540:4522];
assign A[239] = Weights[4559:4541];
assign A[240] = Weights[4578:4560];
assign A[241] = Weights[4597:4579];
assign A[242] = Weights[4616:4598];
assign A[243] = Weights[4635:4617];
assign A[244] = Weights[4654:4636];
assign A[245] = Weights[4673:4655];
assign A[246] = Weights[4692:4674];
assign A[247] = Weights[4711:4693];
assign A[248] = Weights[4730:4712];
assign A[249] = Weights[4749:4731];
assign A[250] = Weights[4768:4750];
assign A[251] = Weights[4787:4769];
assign A[252] = Weights[4806:4788];
assign A[253] = Weights[4825:4807];
assign A[254] = Weights[4844:4826];
assign A[255] = Weights[4863:4845];
assign A[256] = Weights[4882:4864];
assign A[257] = Weights[4901:4883];
assign A[258] = Weights[4920:4902];
assign A[259] = Weights[4939:4921];
assign A[260] = Weights[4958:4940];
assign A[261] = Weights[4977:4959];
assign A[262] = Weights[4996:4978];
assign A[263] = Weights[5015:4997];
assign A[264] = Weights[5034:5016];
assign A[265] = Weights[5053:5035];
assign A[266] = Weights[5072:5054];
assign A[267] = Weights[5091:5073];
assign A[268] = Weights[5110:5092];
assign A[269] = Weights[5129:5111];
assign A[270] = Weights[5148:5130];
assign A[271] = Weights[5167:5149];
assign A[272] = Weights[5186:5168];
assign A[273] = Weights[5205:5187];
assign A[274] = Weights[5224:5206];
assign A[275] = Weights[5243:5225];
assign A[276] = Weights[5262:5244];
assign A[277] = Weights[5281:5263];
assign A[278] = Weights[5300:5282];
assign A[279] = Weights[5319:5301];
assign A[280] = Weights[5338:5320];
assign A[281] = Weights[5357:5339];
assign A[282] = Weights[5376:5358];
assign A[283] = Weights[5395:5377];
assign A[284] = Weights[5414:5396];
assign A[285] = Weights[5433:5415];
assign A[286] = Weights[5452:5434];
assign A[287] = Weights[5471:5453];
assign A[288] = Weights[5490:5472];
assign A[289] = Weights[5509:5491];
assign A[290] = Weights[5528:5510];
assign A[291] = Weights[5547:5529];
assign A[292] = Weights[5566:5548];
assign A[293] = Weights[5585:5567];
assign A[294] = Weights[5604:5586];
assign A[295] = Weights[5623:5605];
assign A[296] = Weights[5642:5624];
assign A[297] = Weights[5661:5643];
assign A[298] = Weights[5680:5662];
assign A[299] = Weights[5699:5681];
assign A[300] = Weights[5718:5700];
assign A[301] = Weights[5737:5719];
assign A[302] = Weights[5756:5738];
assign A[303] = Weights[5775:5757];
assign A[304] = Weights[5794:5776];
assign A[305] = Weights[5813:5795];
assign A[306] = Weights[5832:5814];
assign A[307] = Weights[5851:5833];
assign A[308] = Weights[5870:5852];
assign A[309] = Weights[5889:5871];
assign A[310] = Weights[5908:5890];
assign A[311] = Weights[5927:5909];
assign A[312] = Weights[5946:5928];
assign A[313] = Weights[5965:5947];
assign A[314] = Weights[5984:5966];
assign A[315] = Weights[6003:5985];
assign A[316] = Weights[6022:6004];
assign A[317] = Weights[6041:6023];
assign A[318] = Weights[6060:6042];
assign A[319] = Weights[6079:6061];
assign A[320] = Weights[6098:6080];
assign A[321] = Weights[6117:6099];
assign A[322] = Weights[6136:6118];
assign A[323] = Weights[6155:6137];
assign A[324] = Weights[6174:6156];
assign A[325] = Weights[6193:6175];
assign A[326] = Weights[6212:6194];
assign A[327] = Weights[6231:6213];
assign A[328] = Weights[6250:6232];
assign A[329] = Weights[6269:6251];
assign A[330] = Weights[6288:6270];
assign A[331] = Weights[6307:6289];
assign A[332] = Weights[6326:6308];
assign A[333] = Weights[6345:6327];
assign A[334] = Weights[6364:6346];
assign A[335] = Weights[6383:6365];
assign A[336] = Weights[6402:6384];
assign A[337] = Weights[6421:6403];
assign A[338] = Weights[6440:6422];
assign A[339] = Weights[6459:6441];
assign A[340] = Weights[6478:6460];
assign A[341] = Weights[6497:6479];
assign A[342] = Weights[6516:6498];
assign A[343] = Weights[6535:6517];
assign A[344] = Weights[6554:6536];
assign A[345] = Weights[6573:6555];
assign A[346] = Weights[6592:6574];
assign A[347] = Weights[6611:6593];
assign A[348] = Weights[6630:6612];
assign A[349] = Weights[6649:6631];
assign A[350] = Weights[6668:6650];
assign A[351] = Weights[6687:6669];
assign A[352] = Weights[6706:6688];
assign A[353] = Weights[6725:6707];
assign A[354] = Weights[6744:6726];
assign A[355] = Weights[6763:6745];
assign A[356] = Weights[6782:6764];
assign A[357] = Weights[6801:6783];
assign A[358] = Weights[6820:6802];
assign A[359] = Weights[6839:6821];
assign A[360] = Weights[6858:6840];
assign A[361] = Weights[6877:6859];
assign A[362] = Weights[6896:6878];
assign A[363] = Weights[6915:6897];
assign A[364] = Weights[6934:6916];
assign A[365] = Weights[6953:6935];
assign A[366] = Weights[6972:6954];
assign A[367] = Weights[6991:6973];
assign A[368] = Weights[7010:6992];
assign A[369] = Weights[7029:7011];
assign A[370] = Weights[7048:7030];
assign A[371] = Weights[7067:7049];
assign A[372] = Weights[7086:7068];
assign A[373] = Weights[7105:7087];
assign A[374] = Weights[7124:7106];
assign A[375] = Weights[7143:7125];
assign A[376] = Weights[7162:7144];
assign A[377] = Weights[7181:7163];
assign A[378] = Weights[7200:7182];
assign A[379] = Weights[7219:7201];
assign A[380] = Weights[7238:7220];
assign A[381] = Weights[7257:7239];
assign A[382] = Weights[7276:7258];
assign A[383] = Weights[7295:7277];
assign A[384] = Weights[7314:7296];
assign A[385] = Weights[7333:7315];
assign A[386] = Weights[7352:7334];
assign A[387] = Weights[7371:7353];
assign A[388] = Weights[7390:7372];
assign A[389] = Weights[7409:7391];
assign A[390] = Weights[7428:7410];
assign A[391] = Weights[7447:7429];
assign A[392] = Weights[7466:7448];
assign A[393] = Weights[7485:7467];
assign A[394] = Weights[7504:7486];
assign A[395] = Weights[7523:7505];
assign A[396] = Weights[7542:7524];
assign A[397] = Weights[7561:7543];
assign A[398] = Weights[7580:7562];
assign A[399] = Weights[7599:7581];
assign A[400] = Weights[7618:7600];
assign A[401] = Weights[7637:7619];
assign A[402] = Weights[7656:7638];
assign A[403] = Weights[7675:7657];
assign A[404] = Weights[7694:7676];
assign A[405] = Weights[7713:7695];
assign A[406] = Weights[7732:7714];
assign A[407] = Weights[7751:7733];
assign A[408] = Weights[7770:7752];
assign A[409] = Weights[7789:7771];
assign A[410] = Weights[7808:7790];
assign A[411] = Weights[7827:7809];
assign A[412] = Weights[7846:7828];
assign A[413] = Weights[7865:7847];
assign A[414] = Weights[7884:7866];
assign A[415] = Weights[7903:7885];
assign A[416] = Weights[7922:7904];
assign A[417] = Weights[7941:7923];
assign A[418] = Weights[7960:7942];
assign A[419] = Weights[7979:7961];
assign A[420] = Weights[7998:7980];
assign A[421] = Weights[8017:7999];
assign A[422] = Weights[8036:8018];
assign A[423] = Weights[8055:8037];
assign A[424] = Weights[8074:8056];
assign A[425] = Weights[8093:8075];
assign A[426] = Weights[8112:8094];
assign A[427] = Weights[8131:8113];
assign A[428] = Weights[8150:8132];
assign A[429] = Weights[8169:8151];
assign A[430] = Weights[8188:8170];
assign A[431] = Weights[8207:8189];
assign A[432] = Weights[8226:8208];
assign A[433] = Weights[8245:8227];
assign A[434] = Weights[8264:8246];
assign A[435] = Weights[8283:8265];
assign A[436] = Weights[8302:8284];
assign A[437] = Weights[8321:8303];
assign A[438] = Weights[8340:8322];
assign A[439] = Weights[8359:8341];
assign A[440] = Weights[8378:8360];
assign A[441] = Weights[8397:8379];
assign A[442] = Weights[8416:8398];
assign A[443] = Weights[8435:8417];
assign A[444] = Weights[8454:8436];
assign A[445] = Weights[8473:8455];
assign A[446] = Weights[8492:8474];
assign A[447] = Weights[8511:8493];
assign A[448] = Weights[8530:8512];
assign A[449] = Weights[8549:8531];
assign A[450] = Weights[8568:8550];
assign A[451] = Weights[8587:8569];
assign A[452] = Weights[8606:8588];
assign A[453] = Weights[8625:8607];
assign A[454] = Weights[8644:8626];
assign A[455] = Weights[8663:8645];
assign A[456] = Weights[8682:8664];
assign A[457] = Weights[8701:8683];
assign A[458] = Weights[8720:8702];
assign A[459] = Weights[8739:8721];
assign A[460] = Weights[8758:8740];
assign A[461] = Weights[8777:8759];
assign A[462] = Weights[8796:8778];
assign A[463] = Weights[8815:8797];
assign A[464] = Weights[8834:8816];
assign A[465] = Weights[8853:8835];
assign A[466] = Weights[8872:8854];
assign A[467] = Weights[8891:8873];
assign A[468] = Weights[8910:8892];
assign A[469] = Weights[8929:8911];
assign A[470] = Weights[8948:8930];
assign A[471] = Weights[8967:8949];
assign A[472] = Weights[8986:8968];
assign A[473] = Weights[9005:8987];
assign A[474] = Weights[9024:9006];
assign A[475] = Weights[9043:9025];
assign A[476] = Weights[9062:9044];
assign A[477] = Weights[9081:9063];
assign A[478] = Weights[9100:9082];
assign A[479] = Weights[9119:9101];
assign A[480] = Weights[9138:9120];
assign A[481] = Weights[9157:9139];
assign A[482] = Weights[9176:9158];
assign A[483] = Weights[9195:9177];
assign A[484] = Weights[9214:9196];
assign A[485] = Weights[9233:9215];
assign A[486] = Weights[9252:9234];
assign A[487] = Weights[9271:9253];
assign A[488] = Weights[9290:9272];
assign A[489] = Weights[9309:9291];
assign A[490] = Weights[9328:9310];
assign A[491] = Weights[9347:9329];
assign A[492] = Weights[9366:9348];
assign A[493] = Weights[9385:9367];
assign A[494] = Weights[9404:9386];
assign A[495] = Weights[9423:9405];
assign A[496] = Weights[9442:9424];
assign A[497] = Weights[9461:9443];
assign A[498] = Weights[9480:9462];
assign A[499] = Weights[9499:9481];
assign A[500] = Weights[9518:9500];
assign A[501] = Weights[9537:9519];
assign A[502] = Weights[9556:9538];
assign A[503] = Weights[9575:9557];
assign A[504] = Weights[9594:9576];
assign A[505] = Weights[9613:9595];
assign A[506] = Weights[9632:9614];
assign A[507] = Weights[9651:9633];
assign A[508] = Weights[9670:9652];
assign A[509] = Weights[9689:9671];
assign A[510] = Weights[9708:9690];
assign A[511] = Weights[9727:9709];
assign A[512] = Weights[9746:9728];
assign A[513] = Weights[9765:9747];
assign A[514] = Weights[9784:9766];
assign A[515] = Weights[9803:9785];
assign A[516] = Weights[9822:9804];
assign A[517] = Weights[9841:9823];
assign A[518] = Weights[9860:9842];
assign A[519] = Weights[9879:9861];
assign A[520] = Weights[9898:9880];
assign A[521] = Weights[9917:9899];
assign A[522] = Weights[9936:9918];
assign A[523] = Weights[9955:9937];
assign A[524] = Weights[9974:9956];
assign A[525] = Weights[9993:9975];
assign A[526] = Weights[10012:9994];
assign A[527] = Weights[10031:10013];
assign A[528] = Weights[10050:10032];
assign A[529] = Weights[10069:10051];
assign A[530] = Weights[10088:10070];
assign A[531] = Weights[10107:10089];
assign A[532] = Weights[10126:10108];
assign A[533] = Weights[10145:10127];
assign A[534] = Weights[10164:10146];
assign A[535] = Weights[10183:10165];
assign A[536] = Weights[10202:10184];
assign A[537] = Weights[10221:10203];
assign A[538] = Weights[10240:10222];
assign A[539] = Weights[10259:10241];
assign A[540] = Weights[10278:10260];
assign A[541] = Weights[10297:10279];
assign A[542] = Weights[10316:10298];
assign A[543] = Weights[10335:10317];
assign A[544] = Weights[10354:10336];
assign A[545] = Weights[10373:10355];
assign A[546] = Weights[10392:10374];
assign A[547] = Weights[10411:10393];
assign A[548] = Weights[10430:10412];
assign A[549] = Weights[10449:10431];
assign A[550] = Weights[10468:10450];
assign A[551] = Weights[10487:10469];
assign A[552] = Weights[10506:10488];
assign A[553] = Weights[10525:10507];
assign A[554] = Weights[10544:10526];
assign A[555] = Weights[10563:10545];
assign A[556] = Weights[10582:10564];
assign A[557] = Weights[10601:10583];
assign A[558] = Weights[10620:10602];
assign A[559] = Weights[10639:10621];
assign A[560] = Weights[10658:10640];
assign A[561] = Weights[10677:10659];
assign A[562] = Weights[10696:10678];
assign A[563] = Weights[10715:10697];
assign A[564] = Weights[10734:10716];
assign A[565] = Weights[10753:10735];
assign A[566] = Weights[10772:10754];
assign A[567] = Weights[10791:10773];
assign A[568] = Weights[10810:10792];
assign A[569] = Weights[10829:10811];
assign A[570] = Weights[10848:10830];
assign A[571] = Weights[10867:10849];
assign A[572] = Weights[10886:10868];
assign A[573] = Weights[10905:10887];
assign A[574] = Weights[10924:10906];
assign A[575] = Weights[10943:10925];
assign A[576] = Weights[10962:10944];
assign A[577] = Weights[10981:10963];
assign A[578] = Weights[11000:10982];
assign A[579] = Weights[11019:11001];
assign A[580] = Weights[11038:11020];
assign A[581] = Weights[11057:11039];
assign A[582] = Weights[11076:11058];
assign A[583] = Weights[11095:11077];
assign A[584] = Weights[11114:11096];
assign A[585] = Weights[11133:11115];
assign A[586] = Weights[11152:11134];
assign A[587] = Weights[11171:11153];
assign A[588] = Weights[11190:11172];
assign A[589] = Weights[11209:11191];
assign A[590] = Weights[11228:11210];
assign A[591] = Weights[11247:11229];
assign A[592] = Weights[11266:11248];
assign A[593] = Weights[11285:11267];
assign A[594] = Weights[11304:11286];
assign A[595] = Weights[11323:11305];
assign A[596] = Weights[11342:11324];
assign A[597] = Weights[11361:11343];
assign A[598] = Weights[11380:11362];
assign A[599] = Weights[11399:11381];
assign A[600] = Weights[11418:11400];
assign A[601] = Weights[11437:11419];
assign A[602] = Weights[11456:11438];
assign A[603] = Weights[11475:11457];
assign A[604] = Weights[11494:11476];
assign A[605] = Weights[11513:11495];
assign A[606] = Weights[11532:11514];
assign A[607] = Weights[11551:11533];
assign A[608] = Weights[11570:11552];
assign A[609] = Weights[11589:11571];
assign A[610] = Weights[11608:11590];
assign A[611] = Weights[11627:11609];
assign A[612] = Weights[11646:11628];
assign A[613] = Weights[11665:11647];
assign A[614] = Weights[11684:11666];
assign A[615] = Weights[11703:11685];
assign A[616] = Weights[11722:11704];
assign A[617] = Weights[11741:11723];
assign A[618] = Weights[11760:11742];
assign A[619] = Weights[11779:11761];
assign A[620] = Weights[11798:11780];
assign A[621] = Weights[11817:11799];
assign A[622] = Weights[11836:11818];
assign A[623] = Weights[11855:11837];
assign A[624] = Weights[11874:11856];
assign A[625] = Weights[11893:11875];
assign A[626] = Weights[11912:11894];
assign A[627] = Weights[11931:11913];
assign A[628] = Weights[11950:11932];
assign A[629] = Weights[11969:11951];
assign A[630] = Weights[11988:11970];
assign A[631] = Weights[12007:11989];
assign A[632] = Weights[12026:12008];
assign A[633] = Weights[12045:12027];
assign A[634] = Weights[12064:12046];
assign A[635] = Weights[12083:12065];
assign A[636] = Weights[12102:12084];
assign A[637] = Weights[12121:12103];
assign A[638] = Weights[12140:12122];
assign A[639] = Weights[12159:12141];
assign A[640] = Weights[12178:12160];
assign A[641] = Weights[12197:12179];
assign A[642] = Weights[12216:12198];
assign A[643] = Weights[12235:12217];
assign A[644] = Weights[12254:12236];
assign A[645] = Weights[12273:12255];
assign A[646] = Weights[12292:12274];
assign A[647] = Weights[12311:12293];
assign A[648] = Weights[12330:12312];
assign A[649] = Weights[12349:12331];
assign A[650] = Weights[12368:12350];
assign A[651] = Weights[12387:12369];
assign A[652] = Weights[12406:12388];
assign A[653] = Weights[12425:12407];
assign A[654] = Weights[12444:12426];
assign A[655] = Weights[12463:12445];
assign A[656] = Weights[12482:12464];
assign A[657] = Weights[12501:12483];
assign A[658] = Weights[12520:12502];
assign A[659] = Weights[12539:12521];
assign A[660] = Weights[12558:12540];
assign A[661] = Weights[12577:12559];
assign A[662] = Weights[12596:12578];
assign A[663] = Weights[12615:12597];
assign A[664] = Weights[12634:12616];
assign A[665] = Weights[12653:12635];
assign A[666] = Weights[12672:12654];
assign A[667] = Weights[12691:12673];
assign A[668] = Weights[12710:12692];
assign A[669] = Weights[12729:12711];
assign A[670] = Weights[12748:12730];
assign A[671] = Weights[12767:12749];
assign A[672] = Weights[12786:12768];
assign A[673] = Weights[12805:12787];
assign A[674] = Weights[12824:12806];
assign A[675] = Weights[12843:12825];
assign A[676] = Weights[12862:12844];
assign A[677] = Weights[12881:12863];
assign A[678] = Weights[12900:12882];
assign A[679] = Weights[12919:12901];
assign A[680] = Weights[12938:12920];
assign A[681] = Weights[12957:12939];
assign A[682] = Weights[12976:12958];
assign A[683] = Weights[12995:12977];
assign A[684] = Weights[13014:12996];
assign A[685] = Weights[13033:13015];
assign A[686] = Weights[13052:13034];
assign A[687] = Weights[13071:13053];
assign A[688] = Weights[13090:13072];
assign A[689] = Weights[13109:13091];
assign A[690] = Weights[13128:13110];
assign A[691] = Weights[13147:13129];
assign A[692] = Weights[13166:13148];
assign A[693] = Weights[13185:13167];
assign A[694] = Weights[13204:13186];
assign A[695] = Weights[13223:13205];
assign A[696] = Weights[13242:13224];
assign A[697] = Weights[13261:13243];
assign A[698] = Weights[13280:13262];
assign A[699] = Weights[13299:13281];
assign A[700] = Weights[13318:13300];
assign A[701] = Weights[13337:13319];
assign A[702] = Weights[13356:13338];
assign A[703] = Weights[13375:13357];
assign A[704] = Weights[13394:13376];
assign A[705] = Weights[13413:13395];
assign A[706] = Weights[13432:13414];
assign A[707] = Weights[13451:13433];
assign A[708] = Weights[13470:13452];
assign A[709] = Weights[13489:13471];
assign A[710] = Weights[13508:13490];
assign A[711] = Weights[13527:13509];
assign A[712] = Weights[13546:13528];
assign A[713] = Weights[13565:13547];
assign A[714] = Weights[13584:13566];
assign A[715] = Weights[13603:13585];
assign A[716] = Weights[13622:13604];
assign A[717] = Weights[13641:13623];
assign A[718] = Weights[13660:13642];
assign A[719] = Weights[13679:13661];
assign A[720] = Weights[13698:13680];
assign A[721] = Weights[13717:13699];
assign A[722] = Weights[13736:13718];
assign A[723] = Weights[13755:13737];
assign A[724] = Weights[13774:13756];
assign A[725] = Weights[13793:13775];
assign A[726] = Weights[13812:13794];
assign A[727] = Weights[13831:13813];
assign A[728] = Weights[13850:13832];
assign A[729] = Weights[13869:13851];
assign A[730] = Weights[13888:13870];
assign A[731] = Weights[13907:13889];
assign A[732] = Weights[13926:13908];
assign A[733] = Weights[13945:13927];
assign A[734] = Weights[13964:13946];
assign A[735] = Weights[13983:13965];
assign A[736] = Weights[14002:13984];
assign A[737] = Weights[14021:14003];
assign A[738] = Weights[14040:14022];
assign A[739] = Weights[14059:14041];
assign A[740] = Weights[14078:14060];
assign A[741] = Weights[14097:14079];
assign A[742] = Weights[14116:14098];
assign A[743] = Weights[14135:14117];
assign A[744] = Weights[14154:14136];
assign A[745] = Weights[14173:14155];
assign A[746] = Weights[14192:14174];
assign A[747] = Weights[14211:14193];
assign A[748] = Weights[14230:14212];
assign A[749] = Weights[14249:14231];
assign A[750] = Weights[14268:14250];
assign A[751] = Weights[14287:14269];
assign A[752] = Weights[14306:14288];
assign A[753] = Weights[14325:14307];
assign A[754] = Weights[14344:14326];
assign A[755] = Weights[14363:14345];
assign A[756] = Weights[14382:14364];
assign A[757] = Weights[14401:14383];
assign A[758] = Weights[14420:14402];
assign A[759] = Weights[14439:14421];
assign A[760] = Weights[14458:14440];
assign A[761] = Weights[14477:14459];
assign A[762] = Weights[14496:14478];
assign A[763] = Weights[14515:14497];
assign A[764] = Weights[14534:14516];
assign A[765] = Weights[14553:14535];
assign A[766] = Weights[14572:14554];
assign A[767] = Weights[14591:14573];
assign A[768] = Weights[14610:14592];
assign A[769] = Weights[14629:14611];
assign A[770] = Weights[14648:14630];
assign A[771] = Weights[14667:14649];
assign A[772] = Weights[14686:14668];
assign A[773] = Weights[14705:14687];
assign A[774] = Weights[14724:14706];
assign A[775] = Weights[14743:14725];
assign A[776] = Weights[14762:14744];
assign A[777] = Weights[14781:14763];
assign A[778] = Weights[14800:14782];
assign A[779] = Weights[14819:14801];
assign A[780] = Weights[14838:14820];
assign A[781] = Weights[14857:14839];
assign A[782] = Weights[14876:14858];
assign A[783] = Weights[14895:14877];
assign B[0] = Pixels[9:0];
assign B[1] = Pixels[19:10];
assign B[2] = Pixels[29:20];
assign B[3] = Pixels[39:30];
assign B[4] = Pixels[49:40];
assign B[5] = Pixels[59:50];
assign B[6] = Pixels[69:60];
assign B[7] = Pixels[79:70];
assign B[8] = Pixels[89:80];
assign B[9] = Pixels[99:90];
assign B[10] = Pixels[109:100];
assign B[11] = Pixels[119:110];
assign B[12] = Pixels[129:120];
assign B[13] = Pixels[139:130];
assign B[14] = Pixels[149:140];
assign B[15] = Pixels[159:150];
assign B[16] = Pixels[169:160];
assign B[17] = Pixels[179:170];
assign B[18] = Pixels[189:180];
assign B[19] = Pixels[199:190];
assign B[20] = Pixels[209:200];
assign B[21] = Pixels[219:210];
assign B[22] = Pixels[229:220];
assign B[23] = Pixels[239:230];
assign B[24] = Pixels[249:240];
assign B[25] = Pixels[259:250];
assign B[26] = Pixels[269:260];
assign B[27] = Pixels[279:270];
assign B[28] = Pixels[289:280];
assign B[29] = Pixels[299:290];
assign B[30] = Pixels[309:300];
assign B[31] = Pixels[319:310];
assign B[32] = Pixels[329:320];
assign B[33] = Pixels[339:330];
assign B[34] = Pixels[349:340];
assign B[35] = Pixels[359:350];
assign B[36] = Pixels[369:360];
assign B[37] = Pixels[379:370];
assign B[38] = Pixels[389:380];
assign B[39] = Pixels[399:390];
assign B[40] = Pixels[409:400];
assign B[41] = Pixels[419:410];
assign B[42] = Pixels[429:420];
assign B[43] = Pixels[439:430];
assign B[44] = Pixels[449:440];
assign B[45] = Pixels[459:450];
assign B[46] = Pixels[469:460];
assign B[47] = Pixels[479:470];
assign B[48] = Pixels[489:480];
assign B[49] = Pixels[499:490];
assign B[50] = Pixels[509:500];
assign B[51] = Pixels[519:510];
assign B[52] = Pixels[529:520];
assign B[53] = Pixels[539:530];
assign B[54] = Pixels[549:540];
assign B[55] = Pixels[559:550];
assign B[56] = Pixels[569:560];
assign B[57] = Pixels[579:570];
assign B[58] = Pixels[589:580];
assign B[59] = Pixels[599:590];
assign B[60] = Pixels[609:600];
assign B[61] = Pixels[619:610];
assign B[62] = Pixels[629:620];
assign B[63] = Pixels[639:630];
assign B[64] = Pixels[649:640];
assign B[65] = Pixels[659:650];
assign B[66] = Pixels[669:660];
assign B[67] = Pixels[679:670];
assign B[68] = Pixels[689:680];
assign B[69] = Pixels[699:690];
assign B[70] = Pixels[709:700];
assign B[71] = Pixels[719:710];
assign B[72] = Pixels[729:720];
assign B[73] = Pixels[739:730];
assign B[74] = Pixels[749:740];
assign B[75] = Pixels[759:750];
assign B[76] = Pixels[769:760];
assign B[77] = Pixels[779:770];
assign B[78] = Pixels[789:780];
assign B[79] = Pixels[799:790];
assign B[80] = Pixels[809:800];
assign B[81] = Pixels[819:810];
assign B[82] = Pixels[829:820];
assign B[83] = Pixels[839:830];
assign B[84] = Pixels[849:840];
assign B[85] = Pixels[859:850];
assign B[86] = Pixels[869:860];
assign B[87] = Pixels[879:870];
assign B[88] = Pixels[889:880];
assign B[89] = Pixels[899:890];
assign B[90] = Pixels[909:900];
assign B[91] = Pixels[919:910];
assign B[92] = Pixels[929:920];
assign B[93] = Pixels[939:930];
assign B[94] = Pixels[949:940];
assign B[95] = Pixels[959:950];
assign B[96] = Pixels[969:960];
assign B[97] = Pixels[979:970];
assign B[98] = Pixels[989:980];
assign B[99] = Pixels[999:990];
assign B[100] = Pixels[1009:1000];
assign B[101] = Pixels[1019:1010];
assign B[102] = Pixels[1029:1020];
assign B[103] = Pixels[1039:1030];
assign B[104] = Pixels[1049:1040];
assign B[105] = Pixels[1059:1050];
assign B[106] = Pixels[1069:1060];
assign B[107] = Pixels[1079:1070];
assign B[108] = Pixels[1089:1080];
assign B[109] = Pixels[1099:1090];
assign B[110] = Pixels[1109:1100];
assign B[111] = Pixels[1119:1110];
assign B[112] = Pixels[1129:1120];
assign B[113] = Pixels[1139:1130];
assign B[114] = Pixels[1149:1140];
assign B[115] = Pixels[1159:1150];
assign B[116] = Pixels[1169:1160];
assign B[117] = Pixels[1179:1170];
assign B[118] = Pixels[1189:1180];
assign B[119] = Pixels[1199:1190];
assign B[120] = Pixels[1209:1200];
assign B[121] = Pixels[1219:1210];
assign B[122] = Pixels[1229:1220];
assign B[123] = Pixels[1239:1230];
assign B[124] = Pixels[1249:1240];
assign B[125] = Pixels[1259:1250];
assign B[126] = Pixels[1269:1260];
assign B[127] = Pixels[1279:1270];
assign B[128] = Pixels[1289:1280];
assign B[129] = Pixels[1299:1290];
assign B[130] = Pixels[1309:1300];
assign B[131] = Pixels[1319:1310];
assign B[132] = Pixels[1329:1320];
assign B[133] = Pixels[1339:1330];
assign B[134] = Pixels[1349:1340];
assign B[135] = Pixels[1359:1350];
assign B[136] = Pixels[1369:1360];
assign B[137] = Pixels[1379:1370];
assign B[138] = Pixels[1389:1380];
assign B[139] = Pixels[1399:1390];
assign B[140] = Pixels[1409:1400];
assign B[141] = Pixels[1419:1410];
assign B[142] = Pixels[1429:1420];
assign B[143] = Pixels[1439:1430];
assign B[144] = Pixels[1449:1440];
assign B[145] = Pixels[1459:1450];
assign B[146] = Pixels[1469:1460];
assign B[147] = Pixels[1479:1470];
assign B[148] = Pixels[1489:1480];
assign B[149] = Pixels[1499:1490];
assign B[150] = Pixels[1509:1500];
assign B[151] = Pixels[1519:1510];
assign B[152] = Pixels[1529:1520];
assign B[153] = Pixels[1539:1530];
assign B[154] = Pixels[1549:1540];
assign B[155] = Pixels[1559:1550];
assign B[156] = Pixels[1569:1560];
assign B[157] = Pixels[1579:1570];
assign B[158] = Pixels[1589:1580];
assign B[159] = Pixels[1599:1590];
assign B[160] = Pixels[1609:1600];
assign B[161] = Pixels[1619:1610];
assign B[162] = Pixels[1629:1620];
assign B[163] = Pixels[1639:1630];
assign B[164] = Pixels[1649:1640];
assign B[165] = Pixels[1659:1650];
assign B[166] = Pixels[1669:1660];
assign B[167] = Pixels[1679:1670];
assign B[168] = Pixels[1689:1680];
assign B[169] = Pixels[1699:1690];
assign B[170] = Pixels[1709:1700];
assign B[171] = Pixels[1719:1710];
assign B[172] = Pixels[1729:1720];
assign B[173] = Pixels[1739:1730];
assign B[174] = Pixels[1749:1740];
assign B[175] = Pixels[1759:1750];
assign B[176] = Pixels[1769:1760];
assign B[177] = Pixels[1779:1770];
assign B[178] = Pixels[1789:1780];
assign B[179] = Pixels[1799:1790];
assign B[180] = Pixels[1809:1800];
assign B[181] = Pixels[1819:1810];
assign B[182] = Pixels[1829:1820];
assign B[183] = Pixels[1839:1830];
assign B[184] = Pixels[1849:1840];
assign B[185] = Pixels[1859:1850];
assign B[186] = Pixels[1869:1860];
assign B[187] = Pixels[1879:1870];
assign B[188] = Pixels[1889:1880];
assign B[189] = Pixels[1899:1890];
assign B[190] = Pixels[1909:1900];
assign B[191] = Pixels[1919:1910];
assign B[192] = Pixels[1929:1920];
assign B[193] = Pixels[1939:1930];
assign B[194] = Pixels[1949:1940];
assign B[195] = Pixels[1959:1950];
assign B[196] = Pixels[1969:1960];
assign B[197] = Pixels[1979:1970];
assign B[198] = Pixels[1989:1980];
assign B[199] = Pixels[1999:1990];
assign B[200] = Pixels[2009:2000];
assign B[201] = Pixels[2019:2010];
assign B[202] = Pixels[2029:2020];
assign B[203] = Pixels[2039:2030];
assign B[204] = Pixels[2049:2040];
assign B[205] = Pixels[2059:2050];
assign B[206] = Pixels[2069:2060];
assign B[207] = Pixels[2079:2070];
assign B[208] = Pixels[2089:2080];
assign B[209] = Pixels[2099:2090];
assign B[210] = Pixels[2109:2100];
assign B[211] = Pixels[2119:2110];
assign B[212] = Pixels[2129:2120];
assign B[213] = Pixels[2139:2130];
assign B[214] = Pixels[2149:2140];
assign B[215] = Pixels[2159:2150];
assign B[216] = Pixels[2169:2160];
assign B[217] = Pixels[2179:2170];
assign B[218] = Pixels[2189:2180];
assign B[219] = Pixels[2199:2190];
assign B[220] = Pixels[2209:2200];
assign B[221] = Pixels[2219:2210];
assign B[222] = Pixels[2229:2220];
assign B[223] = Pixels[2239:2230];
assign B[224] = Pixels[2249:2240];
assign B[225] = Pixels[2259:2250];
assign B[226] = Pixels[2269:2260];
assign B[227] = Pixels[2279:2270];
assign B[228] = Pixels[2289:2280];
assign B[229] = Pixels[2299:2290];
assign B[230] = Pixels[2309:2300];
assign B[231] = Pixels[2319:2310];
assign B[232] = Pixels[2329:2320];
assign B[233] = Pixels[2339:2330];
assign B[234] = Pixels[2349:2340];
assign B[235] = Pixels[2359:2350];
assign B[236] = Pixels[2369:2360];
assign B[237] = Pixels[2379:2370];
assign B[238] = Pixels[2389:2380];
assign B[239] = Pixels[2399:2390];
assign B[240] = Pixels[2409:2400];
assign B[241] = Pixels[2419:2410];
assign B[242] = Pixels[2429:2420];
assign B[243] = Pixels[2439:2430];
assign B[244] = Pixels[2449:2440];
assign B[245] = Pixels[2459:2450];
assign B[246] = Pixels[2469:2460];
assign B[247] = Pixels[2479:2470];
assign B[248] = Pixels[2489:2480];
assign B[249] = Pixels[2499:2490];
assign B[250] = Pixels[2509:2500];
assign B[251] = Pixels[2519:2510];
assign B[252] = Pixels[2529:2520];
assign B[253] = Pixels[2539:2530];
assign B[254] = Pixels[2549:2540];
assign B[255] = Pixels[2559:2550];
assign B[256] = Pixels[2569:2560];
assign B[257] = Pixels[2579:2570];
assign B[258] = Pixels[2589:2580];
assign B[259] = Pixels[2599:2590];
assign B[260] = Pixels[2609:2600];
assign B[261] = Pixels[2619:2610];
assign B[262] = Pixels[2629:2620];
assign B[263] = Pixels[2639:2630];
assign B[264] = Pixels[2649:2640];
assign B[265] = Pixels[2659:2650];
assign B[266] = Pixels[2669:2660];
assign B[267] = Pixels[2679:2670];
assign B[268] = Pixels[2689:2680];
assign B[269] = Pixels[2699:2690];
assign B[270] = Pixels[2709:2700];
assign B[271] = Pixels[2719:2710];
assign B[272] = Pixels[2729:2720];
assign B[273] = Pixels[2739:2730];
assign B[274] = Pixels[2749:2740];
assign B[275] = Pixels[2759:2750];
assign B[276] = Pixels[2769:2760];
assign B[277] = Pixels[2779:2770];
assign B[278] = Pixels[2789:2780];
assign B[279] = Pixels[2799:2790];
assign B[280] = Pixels[2809:2800];
assign B[281] = Pixels[2819:2810];
assign B[282] = Pixels[2829:2820];
assign B[283] = Pixels[2839:2830];
assign B[284] = Pixels[2849:2840];
assign B[285] = Pixels[2859:2850];
assign B[286] = Pixels[2869:2860];
assign B[287] = Pixels[2879:2870];
assign B[288] = Pixels[2889:2880];
assign B[289] = Pixels[2899:2890];
assign B[290] = Pixels[2909:2900];
assign B[291] = Pixels[2919:2910];
assign B[292] = Pixels[2929:2920];
assign B[293] = Pixels[2939:2930];
assign B[294] = Pixels[2949:2940];
assign B[295] = Pixels[2959:2950];
assign B[296] = Pixels[2969:2960];
assign B[297] = Pixels[2979:2970];
assign B[298] = Pixels[2989:2980];
assign B[299] = Pixels[2999:2990];
assign B[300] = Pixels[3009:3000];
assign B[301] = Pixels[3019:3010];
assign B[302] = Pixels[3029:3020];
assign B[303] = Pixels[3039:3030];
assign B[304] = Pixels[3049:3040];
assign B[305] = Pixels[3059:3050];
assign B[306] = Pixels[3069:3060];
assign B[307] = Pixels[3079:3070];
assign B[308] = Pixels[3089:3080];
assign B[309] = Pixels[3099:3090];
assign B[310] = Pixels[3109:3100];
assign B[311] = Pixels[3119:3110];
assign B[312] = Pixels[3129:3120];
assign B[313] = Pixels[3139:3130];
assign B[314] = Pixels[3149:3140];
assign B[315] = Pixels[3159:3150];
assign B[316] = Pixels[3169:3160];
assign B[317] = Pixels[3179:3170];
assign B[318] = Pixels[3189:3180];
assign B[319] = Pixels[3199:3190];
assign B[320] = Pixels[3209:3200];
assign B[321] = Pixels[3219:3210];
assign B[322] = Pixels[3229:3220];
assign B[323] = Pixels[3239:3230];
assign B[324] = Pixels[3249:3240];
assign B[325] = Pixels[3259:3250];
assign B[326] = Pixels[3269:3260];
assign B[327] = Pixels[3279:3270];
assign B[328] = Pixels[3289:3280];
assign B[329] = Pixels[3299:3290];
assign B[330] = Pixels[3309:3300];
assign B[331] = Pixels[3319:3310];
assign B[332] = Pixels[3329:3320];
assign B[333] = Pixels[3339:3330];
assign B[334] = Pixels[3349:3340];
assign B[335] = Pixels[3359:3350];
assign B[336] = Pixels[3369:3360];
assign B[337] = Pixels[3379:3370];
assign B[338] = Pixels[3389:3380];
assign B[339] = Pixels[3399:3390];
assign B[340] = Pixels[3409:3400];
assign B[341] = Pixels[3419:3410];
assign B[342] = Pixels[3429:3420];
assign B[343] = Pixels[3439:3430];
assign B[344] = Pixels[3449:3440];
assign B[345] = Pixels[3459:3450];
assign B[346] = Pixels[3469:3460];
assign B[347] = Pixels[3479:3470];
assign B[348] = Pixels[3489:3480];
assign B[349] = Pixels[3499:3490];
assign B[350] = Pixels[3509:3500];
assign B[351] = Pixels[3519:3510];
assign B[352] = Pixels[3529:3520];
assign B[353] = Pixels[3539:3530];
assign B[354] = Pixels[3549:3540];
assign B[355] = Pixels[3559:3550];
assign B[356] = Pixels[3569:3560];
assign B[357] = Pixels[3579:3570];
assign B[358] = Pixels[3589:3580];
assign B[359] = Pixels[3599:3590];
assign B[360] = Pixels[3609:3600];
assign B[361] = Pixels[3619:3610];
assign B[362] = Pixels[3629:3620];
assign B[363] = Pixels[3639:3630];
assign B[364] = Pixels[3649:3640];
assign B[365] = Pixels[3659:3650];
assign B[366] = Pixels[3669:3660];
assign B[367] = Pixels[3679:3670];
assign B[368] = Pixels[3689:3680];
assign B[369] = Pixels[3699:3690];
assign B[370] = Pixels[3709:3700];
assign B[371] = Pixels[3719:3710];
assign B[372] = Pixels[3729:3720];
assign B[373] = Pixels[3739:3730];
assign B[374] = Pixels[3749:3740];
assign B[375] = Pixels[3759:3750];
assign B[376] = Pixels[3769:3760];
assign B[377] = Pixels[3779:3770];
assign B[378] = Pixels[3789:3780];
assign B[379] = Pixels[3799:3790];
assign B[380] = Pixels[3809:3800];
assign B[381] = Pixels[3819:3810];
assign B[382] = Pixels[3829:3820];
assign B[383] = Pixels[3839:3830];
assign B[384] = Pixels[3849:3840];
assign B[385] = Pixels[3859:3850];
assign B[386] = Pixels[3869:3860];
assign B[387] = Pixels[3879:3870];
assign B[388] = Pixels[3889:3880];
assign B[389] = Pixels[3899:3890];
assign B[390] = Pixels[3909:3900];
assign B[391] = Pixels[3919:3910];
assign B[392] = Pixels[3929:3920];
assign B[393] = Pixels[3939:3930];
assign B[394] = Pixels[3949:3940];
assign B[395] = Pixels[3959:3950];
assign B[396] = Pixels[3969:3960];
assign B[397] = Pixels[3979:3970];
assign B[398] = Pixels[3989:3980];
assign B[399] = Pixels[3999:3990];
assign B[400] = Pixels[4009:4000];
assign B[401] = Pixels[4019:4010];
assign B[402] = Pixels[4029:4020];
assign B[403] = Pixels[4039:4030];
assign B[404] = Pixels[4049:4040];
assign B[405] = Pixels[4059:4050];
assign B[406] = Pixels[4069:4060];
assign B[407] = Pixels[4079:4070];
assign B[408] = Pixels[4089:4080];
assign B[409] = Pixels[4099:4090];
assign B[410] = Pixels[4109:4100];
assign B[411] = Pixels[4119:4110];
assign B[412] = Pixels[4129:4120];
assign B[413] = Pixels[4139:4130];
assign B[414] = Pixels[4149:4140];
assign B[415] = Pixels[4159:4150];
assign B[416] = Pixels[4169:4160];
assign B[417] = Pixels[4179:4170];
assign B[418] = Pixels[4189:4180];
assign B[419] = Pixels[4199:4190];
assign B[420] = Pixels[4209:4200];
assign B[421] = Pixels[4219:4210];
assign B[422] = Pixels[4229:4220];
assign B[423] = Pixels[4239:4230];
assign B[424] = Pixels[4249:4240];
assign B[425] = Pixels[4259:4250];
assign B[426] = Pixels[4269:4260];
assign B[427] = Pixels[4279:4270];
assign B[428] = Pixels[4289:4280];
assign B[429] = Pixels[4299:4290];
assign B[430] = Pixels[4309:4300];
assign B[431] = Pixels[4319:4310];
assign B[432] = Pixels[4329:4320];
assign B[433] = Pixels[4339:4330];
assign B[434] = Pixels[4349:4340];
assign B[435] = Pixels[4359:4350];
assign B[436] = Pixels[4369:4360];
assign B[437] = Pixels[4379:4370];
assign B[438] = Pixels[4389:4380];
assign B[439] = Pixels[4399:4390];
assign B[440] = Pixels[4409:4400];
assign B[441] = Pixels[4419:4410];
assign B[442] = Pixels[4429:4420];
assign B[443] = Pixels[4439:4430];
assign B[444] = Pixels[4449:4440];
assign B[445] = Pixels[4459:4450];
assign B[446] = Pixels[4469:4460];
assign B[447] = Pixels[4479:4470];
assign B[448] = Pixels[4489:4480];
assign B[449] = Pixels[4499:4490];
assign B[450] = Pixels[4509:4500];
assign B[451] = Pixels[4519:4510];
assign B[452] = Pixels[4529:4520];
assign B[453] = Pixels[4539:4530];
assign B[454] = Pixels[4549:4540];
assign B[455] = Pixels[4559:4550];
assign B[456] = Pixels[4569:4560];
assign B[457] = Pixels[4579:4570];
assign B[458] = Pixels[4589:4580];
assign B[459] = Pixels[4599:4590];
assign B[460] = Pixels[4609:4600];
assign B[461] = Pixels[4619:4610];
assign B[462] = Pixels[4629:4620];
assign B[463] = Pixels[4639:4630];
assign B[464] = Pixels[4649:4640];
assign B[465] = Pixels[4659:4650];
assign B[466] = Pixels[4669:4660];
assign B[467] = Pixels[4679:4670];
assign B[468] = Pixels[4689:4680];
assign B[469] = Pixels[4699:4690];
assign B[470] = Pixels[4709:4700];
assign B[471] = Pixels[4719:4710];
assign B[472] = Pixels[4729:4720];
assign B[473] = Pixels[4739:4730];
assign B[474] = Pixels[4749:4740];
assign B[475] = Pixels[4759:4750];
assign B[476] = Pixels[4769:4760];
assign B[477] = Pixels[4779:4770];
assign B[478] = Pixels[4789:4780];
assign B[479] = Pixels[4799:4790];
assign B[480] = Pixels[4809:4800];
assign B[481] = Pixels[4819:4810];
assign B[482] = Pixels[4829:4820];
assign B[483] = Pixels[4839:4830];
assign B[484] = Pixels[4849:4840];
assign B[485] = Pixels[4859:4850];
assign B[486] = Pixels[4869:4860];
assign B[487] = Pixels[4879:4870];
assign B[488] = Pixels[4889:4880];
assign B[489] = Pixels[4899:4890];
assign B[490] = Pixels[4909:4900];
assign B[491] = Pixels[4919:4910];
assign B[492] = Pixels[4929:4920];
assign B[493] = Pixels[4939:4930];
assign B[494] = Pixels[4949:4940];
assign B[495] = Pixels[4959:4950];
assign B[496] = Pixels[4969:4960];
assign B[497] = Pixels[4979:4970];
assign B[498] = Pixels[4989:4980];
assign B[499] = Pixels[4999:4990];
assign B[500] = Pixels[5009:5000];
assign B[501] = Pixels[5019:5010];
assign B[502] = Pixels[5029:5020];
assign B[503] = Pixels[5039:5030];
assign B[504] = Pixels[5049:5040];
assign B[505] = Pixels[5059:5050];
assign B[506] = Pixels[5069:5060];
assign B[507] = Pixels[5079:5070];
assign B[508] = Pixels[5089:5080];
assign B[509] = Pixels[5099:5090];
assign B[510] = Pixels[5109:5100];
assign B[511] = Pixels[5119:5110];
assign B[512] = Pixels[5129:5120];
assign B[513] = Pixels[5139:5130];
assign B[514] = Pixels[5149:5140];
assign B[515] = Pixels[5159:5150];
assign B[516] = Pixels[5169:5160];
assign B[517] = Pixels[5179:5170];
assign B[518] = Pixels[5189:5180];
assign B[519] = Pixels[5199:5190];
assign B[520] = Pixels[5209:5200];
assign B[521] = Pixels[5219:5210];
assign B[522] = Pixels[5229:5220];
assign B[523] = Pixels[5239:5230];
assign B[524] = Pixels[5249:5240];
assign B[525] = Pixels[5259:5250];
assign B[526] = Pixels[5269:5260];
assign B[527] = Pixels[5279:5270];
assign B[528] = Pixels[5289:5280];
assign B[529] = Pixels[5299:5290];
assign B[530] = Pixels[5309:5300];
assign B[531] = Pixels[5319:5310];
assign B[532] = Pixels[5329:5320];
assign B[533] = Pixels[5339:5330];
assign B[534] = Pixels[5349:5340];
assign B[535] = Pixels[5359:5350];
assign B[536] = Pixels[5369:5360];
assign B[537] = Pixels[5379:5370];
assign B[538] = Pixels[5389:5380];
assign B[539] = Pixels[5399:5390];
assign B[540] = Pixels[5409:5400];
assign B[541] = Pixels[5419:5410];
assign B[542] = Pixels[5429:5420];
assign B[543] = Pixels[5439:5430];
assign B[544] = Pixels[5449:5440];
assign B[545] = Pixels[5459:5450];
assign B[546] = Pixels[5469:5460];
assign B[547] = Pixels[5479:5470];
assign B[548] = Pixels[5489:5480];
assign B[549] = Pixels[5499:5490];
assign B[550] = Pixels[5509:5500];
assign B[551] = Pixels[5519:5510];
assign B[552] = Pixels[5529:5520];
assign B[553] = Pixels[5539:5530];
assign B[554] = Pixels[5549:5540];
assign B[555] = Pixels[5559:5550];
assign B[556] = Pixels[5569:5560];
assign B[557] = Pixels[5579:5570];
assign B[558] = Pixels[5589:5580];
assign B[559] = Pixels[5599:5590];
assign B[560] = Pixels[5609:5600];
assign B[561] = Pixels[5619:5610];
assign B[562] = Pixels[5629:5620];
assign B[563] = Pixels[5639:5630];
assign B[564] = Pixels[5649:5640];
assign B[565] = Pixels[5659:5650];
assign B[566] = Pixels[5669:5660];
assign B[567] = Pixels[5679:5670];
assign B[568] = Pixels[5689:5680];
assign B[569] = Pixels[5699:5690];
assign B[570] = Pixels[5709:5700];
assign B[571] = Pixels[5719:5710];
assign B[572] = Pixels[5729:5720];
assign B[573] = Pixels[5739:5730];
assign B[574] = Pixels[5749:5740];
assign B[575] = Pixels[5759:5750];
assign B[576] = Pixels[5769:5760];
assign B[577] = Pixels[5779:5770];
assign B[578] = Pixels[5789:5780];
assign B[579] = Pixels[5799:5790];
assign B[580] = Pixels[5809:5800];
assign B[581] = Pixels[5819:5810];
assign B[582] = Pixels[5829:5820];
assign B[583] = Pixels[5839:5830];
assign B[584] = Pixels[5849:5840];
assign B[585] = Pixels[5859:5850];
assign B[586] = Pixels[5869:5860];
assign B[587] = Pixels[5879:5870];
assign B[588] = Pixels[5889:5880];
assign B[589] = Pixels[5899:5890];
assign B[590] = Pixels[5909:5900];
assign B[591] = Pixels[5919:5910];
assign B[592] = Pixels[5929:5920];
assign B[593] = Pixels[5939:5930];
assign B[594] = Pixels[5949:5940];
assign B[595] = Pixels[5959:5950];
assign B[596] = Pixels[5969:5960];
assign B[597] = Pixels[5979:5970];
assign B[598] = Pixels[5989:5980];
assign B[599] = Pixels[5999:5990];
assign B[600] = Pixels[6009:6000];
assign B[601] = Pixels[6019:6010];
assign B[602] = Pixels[6029:6020];
assign B[603] = Pixels[6039:6030];
assign B[604] = Pixels[6049:6040];
assign B[605] = Pixels[6059:6050];
assign B[606] = Pixels[6069:6060];
assign B[607] = Pixels[6079:6070];
assign B[608] = Pixels[6089:6080];
assign B[609] = Pixels[6099:6090];
assign B[610] = Pixels[6109:6100];
assign B[611] = Pixels[6119:6110];
assign B[612] = Pixels[6129:6120];
assign B[613] = Pixels[6139:6130];
assign B[614] = Pixels[6149:6140];
assign B[615] = Pixels[6159:6150];
assign B[616] = Pixels[6169:6160];
assign B[617] = Pixels[6179:6170];
assign B[618] = Pixels[6189:6180];
assign B[619] = Pixels[6199:6190];
assign B[620] = Pixels[6209:6200];
assign B[621] = Pixels[6219:6210];
assign B[622] = Pixels[6229:6220];
assign B[623] = Pixels[6239:6230];
assign B[624] = Pixels[6249:6240];
assign B[625] = Pixels[6259:6250];
assign B[626] = Pixels[6269:6260];
assign B[627] = Pixels[6279:6270];
assign B[628] = Pixels[6289:6280];
assign B[629] = Pixels[6299:6290];
assign B[630] = Pixels[6309:6300];
assign B[631] = Pixels[6319:6310];
assign B[632] = Pixels[6329:6320];
assign B[633] = Pixels[6339:6330];
assign B[634] = Pixels[6349:6340];
assign B[635] = Pixels[6359:6350];
assign B[636] = Pixels[6369:6360];
assign B[637] = Pixels[6379:6370];
assign B[638] = Pixels[6389:6380];
assign B[639] = Pixels[6399:6390];
assign B[640] = Pixels[6409:6400];
assign B[641] = Pixels[6419:6410];
assign B[642] = Pixels[6429:6420];
assign B[643] = Pixels[6439:6430];
assign B[644] = Pixels[6449:6440];
assign B[645] = Pixels[6459:6450];
assign B[646] = Pixels[6469:6460];
assign B[647] = Pixels[6479:6470];
assign B[648] = Pixels[6489:6480];
assign B[649] = Pixels[6499:6490];
assign B[650] = Pixels[6509:6500];
assign B[651] = Pixels[6519:6510];
assign B[652] = Pixels[6529:6520];
assign B[653] = Pixels[6539:6530];
assign B[654] = Pixels[6549:6540];
assign B[655] = Pixels[6559:6550];
assign B[656] = Pixels[6569:6560];
assign B[657] = Pixels[6579:6570];
assign B[658] = Pixels[6589:6580];
assign B[659] = Pixels[6599:6590];
assign B[660] = Pixels[6609:6600];
assign B[661] = Pixels[6619:6610];
assign B[662] = Pixels[6629:6620];
assign B[663] = Pixels[6639:6630];
assign B[664] = Pixels[6649:6640];
assign B[665] = Pixels[6659:6650];
assign B[666] = Pixels[6669:6660];
assign B[667] = Pixels[6679:6670];
assign B[668] = Pixels[6689:6680];
assign B[669] = Pixels[6699:6690];
assign B[670] = Pixels[6709:6700];
assign B[671] = Pixels[6719:6710];
assign B[672] = Pixels[6729:6720];
assign B[673] = Pixels[6739:6730];
assign B[674] = Pixels[6749:6740];
assign B[675] = Pixels[6759:6750];
assign B[676] = Pixels[6769:6760];
assign B[677] = Pixels[6779:6770];
assign B[678] = Pixels[6789:6780];
assign B[679] = Pixels[6799:6790];
assign B[680] = Pixels[6809:6800];
assign B[681] = Pixels[6819:6810];
assign B[682] = Pixels[6829:6820];
assign B[683] = Pixels[6839:6830];
assign B[684] = Pixels[6849:6840];
assign B[685] = Pixels[6859:6850];
assign B[686] = Pixels[6869:6860];
assign B[687] = Pixels[6879:6870];
assign B[688] = Pixels[6889:6880];
assign B[689] = Pixels[6899:6890];
assign B[690] = Pixels[6909:6900];
assign B[691] = Pixels[6919:6910];
assign B[692] = Pixels[6929:6920];
assign B[693] = Pixels[6939:6930];
assign B[694] = Pixels[6949:6940];
assign B[695] = Pixels[6959:6950];
assign B[696] = Pixels[6969:6960];
assign B[697] = Pixels[6979:6970];
assign B[698] = Pixels[6989:6980];
assign B[699] = Pixels[6999:6990];
assign B[700] = Pixels[7009:7000];
assign B[701] = Pixels[7019:7010];
assign B[702] = Pixels[7029:7020];
assign B[703] = Pixels[7039:7030];
assign B[704] = Pixels[7049:7040];
assign B[705] = Pixels[7059:7050];
assign B[706] = Pixels[7069:7060];
assign B[707] = Pixels[7079:7070];
assign B[708] = Pixels[7089:7080];
assign B[709] = Pixels[7099:7090];
assign B[710] = Pixels[7109:7100];
assign B[711] = Pixels[7119:7110];
assign B[712] = Pixels[7129:7120];
assign B[713] = Pixels[7139:7130];
assign B[714] = Pixels[7149:7140];
assign B[715] = Pixels[7159:7150];
assign B[716] = Pixels[7169:7160];
assign B[717] = Pixels[7179:7170];
assign B[718] = Pixels[7189:7180];
assign B[719] = Pixels[7199:7190];
assign B[720] = Pixels[7209:7200];
assign B[721] = Pixels[7219:7210];
assign B[722] = Pixels[7229:7220];
assign B[723] = Pixels[7239:7230];
assign B[724] = Pixels[7249:7240];
assign B[725] = Pixels[7259:7250];
assign B[726] = Pixels[7269:7260];
assign B[727] = Pixels[7279:7270];
assign B[728] = Pixels[7289:7280];
assign B[729] = Pixels[7299:7290];
assign B[730] = Pixels[7309:7300];
assign B[731] = Pixels[7319:7310];
assign B[732] = Pixels[7329:7320];
assign B[733] = Pixels[7339:7330];
assign B[734] = Pixels[7349:7340];
assign B[735] = Pixels[7359:7350];
assign B[736] = Pixels[7369:7360];
assign B[737] = Pixels[7379:7370];
assign B[738] = Pixels[7389:7380];
assign B[739] = Pixels[7399:7390];
assign B[740] = Pixels[7409:7400];
assign B[741] = Pixels[7419:7410];
assign B[742] = Pixels[7429:7420];
assign B[743] = Pixels[7439:7430];
assign B[744] = Pixels[7449:7440];
assign B[745] = Pixels[7459:7450];
assign B[746] = Pixels[7469:7460];
assign B[747] = Pixels[7479:7470];
assign B[748] = Pixels[7489:7480];
assign B[749] = Pixels[7499:7490];
assign B[750] = Pixels[7509:7500];
assign B[751] = Pixels[7519:7510];
assign B[752] = Pixels[7529:7520];
assign B[753] = Pixels[7539:7530];
assign B[754] = Pixels[7549:7540];
assign B[755] = Pixels[7559:7550];
assign B[756] = Pixels[7569:7560];
assign B[757] = Pixels[7579:7570];
assign B[758] = Pixels[7589:7580];
assign B[759] = Pixels[7599:7590];
assign B[760] = Pixels[7609:7600];
assign B[761] = Pixels[7619:7610];
assign B[762] = Pixels[7629:7620];
assign B[763] = Pixels[7639:7630];
assign B[764] = Pixels[7649:7640];
assign B[765] = Pixels[7659:7650];
assign B[766] = Pixels[7669:7660];
assign B[767] = Pixels[7679:7670];
assign B[768] = Pixels[7689:7680];
assign B[769] = Pixels[7699:7690];
assign B[770] = Pixels[7709:7700];
assign B[771] = Pixels[7719:7710];
assign B[772] = Pixels[7729:7720];
assign B[773] = Pixels[7739:7730];
assign B[774] = Pixels[7749:7740];
assign B[775] = Pixels[7759:7750];
assign B[776] = Pixels[7769:7760];
assign B[777] = Pixels[7779:7770];
assign B[778] = Pixels[7789:7780];
assign B[779] = Pixels[7799:7790];
assign B[780] = Pixels[7809:7800];
assign B[781] = Pixels[7819:7810];
assign B[782] = Pixels[7829:7820];
assign B[783] = Pixels[7839:7830];

FixedPointMultiplier FPM1(.clk(clk),.GlobalReset(GlobalReset),.WeightPort(A1),.PixelPort(B1),.Output_syn(FPMAns1));
FixedPointMultiplier FPM2(.clk(clk),.GlobalReset(GlobalReset),.WeightPort(A2),.PixelPort(B2),.Output_syn(FPMAns2));
FixedPointAdder FPA1(.clk(clk),.GlobalReset(GlobalReset),.Port2(addInput[1]),.Port1(addInput[0]),.Output_syn(FPAAns));

always@(posedge clk)begin
	if(GlobalReset == 1'b1)begin
		A1 <= A[0];
		A2 <= A[392];
		B1 <= B[0];
		B2 <= B[392];
		addInput[0] <= 26'd0;
		addInput[1] <= 26'd0;
		switchCounter <= 32'd0;
		addAns[0] <= 26'd0;
		addAns[1] <= 26'd0;
		addAns[2] <= 26'd0;
		addAns[3] <= 26'd0;
		addAns[4] <= 26'd0;
		addAns[5] <= 26'd0;
		addAns[6] <= 26'd0;
		addAns[7] <= 26'd0;
		addAns[8] <= 26'd0;
		addAns[9] <= 26'd0;
		addAns[10] <= 26'd0;
		addAns[11] <= 26'd0;
		addAns[12] <= 26'd0;
		addAns[13] <= 26'd0;
		addAns[14] <= 26'd0;
		addAns[15] <= 26'd0;
		addAns[16] <= 26'd0;
		addAns[17] <= 26'd0;
		addAns[18] <= 26'd0;
		addAns[19] <= 26'd0;
		addAns[20] <= 26'd0;
		addAns[21] <= 26'd0;
		addAns[22] <= 26'd0;
		addAns[23] <= 26'd0;
		addAns[24] <= 26'd0;
		addAns[25] <= 26'd0;
		addAns[26] <= 26'd0;
		addAns[27] <= 26'd0;
		addAns[28] <= 26'd0;
		addAns[29] <= 26'd0;
		addAns[30] <= 26'd0;
		addAns[31] <= 26'd0;
		addAns[32] <= 26'd0;
		addAns[33] <= 26'd0;
		addAns[34] <= 26'd0;
		addAns[35] <= 26'd0;
		addAns[36] <= 26'd0;
		addAns[37] <= 26'd0;
		addAns[38] <= 26'd0;
		addAns[39] <= 26'd0;
		addAns[40] <= 26'd0;
		addAns[41] <= 26'd0;
		addAns[42] <= 26'd0;
		addAns[43] <= 26'd0;
		addAns[44] <= 26'd0;
		addAns[45] <= 26'd0;
		addAns[46] <= 26'd0;
		addAns[47] <= 26'd0;
		addAns[48] <= 26'd0;
		addAns[49] <= 26'd0;
		addAns[50] <= 26'd0;
		addAns[51] <= 26'd0;
		addAns[52] <= 26'd0;
		addAns[53] <= 26'd0;
		addAns[54] <= 26'd0;
		addAns[55] <= 26'd0;
		addAns[56] <= 26'd0;
		addAns[57] <= 26'd0;
		addAns[58] <= 26'd0;
		addAns[59] <= 26'd0;
		addAns[60] <= 26'd0;
		addAns[61] <= 26'd0;
		addAns[62] <= 26'd0;
		addAns[63] <= 26'd0;
		addAns[64] <= 26'd0;
		addAns[65] <= 26'd0;
		addAns[66] <= 26'd0;
		addAns[67] <= 26'd0;
		addAns[68] <= 26'd0;
		addAns[69] <= 26'd0;
		addAns[70] <= 26'd0;
		addAns[71] <= 26'd0;
		addAns[72] <= 26'd0;
		addAns[73] <= 26'd0;
		addAns[74] <= 26'd0;
		addAns[75] <= 26'd0;
		addAns[76] <= 26'd0;
		addAns[77] <= 26'd0;
		addAns[78] <= 26'd0;
		addAns[79] <= 26'd0;
		addAns[80] <= 26'd0;
		addAns[81] <= 26'd0;
		addAns[82] <= 26'd0;
		addAns[83] <= 26'd0;
		addAns[84] <= 26'd0;
		addAns[85] <= 26'd0;
		addAns[86] <= 26'd0;
		addAns[87] <= 26'd0;
		addAns[88] <= 26'd0;
		addAns[89] <= 26'd0;
		addAns[90] <= 26'd0;
		addAns[91] <= 26'd0;
		addAns[92] <= 26'd0;
		addAns[93] <= 26'd0;
		addAns[94] <= 26'd0;
		addAns[95] <= 26'd0;
		addAns[96] <= 26'd0;
		addAns[97] <= 26'd0;
		addAns[98] <= 26'd0;
		addAns[99] <= 26'd0;
		addAns[100] <= 26'd0;
		addAns[101] <= 26'd0;
		addAns[102] <= 26'd0;
		addAns[103] <= 26'd0;
		addAns[104] <= 26'd0;
		addAns[105] <= 26'd0;
		addAns[106] <= 26'd0;
		addAns[107] <= 26'd0;
		addAns[108] <= 26'd0;
		addAns[109] <= 26'd0;
		addAns[110] <= 26'd0;
		addAns[111] <= 26'd0;
		addAns[112] <= 26'd0;
		addAns[113] <= 26'd0;
		addAns[114] <= 26'd0;
		addAns[115] <= 26'd0;
		addAns[116] <= 26'd0;
		addAns[117] <= 26'd0;
		addAns[118] <= 26'd0;
		addAns[119] <= 26'd0;
		addAns[120] <= 26'd0;
		addAns[121] <= 26'd0;
		addAns[122] <= 26'd0;
		addAns[123] <= 26'd0;
		addAns[124] <= 26'd0;
		addAns[125] <= 26'd0;
		addAns[126] <= 26'd0;
		addAns[127] <= 26'd0;
		addAns[128] <= 26'd0;
		addAns[129] <= 26'd0;
		addAns[130] <= 26'd0;
		addAns[131] <= 26'd0;
		addAns[132] <= 26'd0;
		addAns[133] <= 26'd0;
		addAns[134] <= 26'd0;
		addAns[135] <= 26'd0;
		addAns[136] <= 26'd0;
		addAns[137] <= 26'd0;
		addAns[138] <= 26'd0;
		addAns[139] <= 26'd0;
		addAns[140] <= 26'd0;
		addAns[141] <= 26'd0;
		addAns[142] <= 26'd0;
		addAns[143] <= 26'd0;
		addAns[144] <= 26'd0;
		addAns[145] <= 26'd0;
		addAns[146] <= 26'd0;
		addAns[147] <= 26'd0;
		addAns[148] <= 26'd0;
		addAns[149] <= 26'd0;
		addAns[150] <= 26'd0;
		addAns[151] <= 26'd0;
		addAns[152] <= 26'd0;
		addAns[153] <= 26'd0;
		addAns[154] <= 26'd0;
		addAns[155] <= 26'd0;
		addAns[156] <= 26'd0;
		addAns[157] <= 26'd0;
		addAns[158] <= 26'd0;
		addAns[159] <= 26'd0;
		addAns[160] <= 26'd0;
		addAns[161] <= 26'd0;
		addAns[162] <= 26'd0;
		addAns[163] <= 26'd0;
		addAns[164] <= 26'd0;
		addAns[165] <= 26'd0;
		addAns[166] <= 26'd0;
		addAns[167] <= 26'd0;
		addAns[168] <= 26'd0;
		addAns[169] <= 26'd0;
		addAns[170] <= 26'd0;
		addAns[171] <= 26'd0;
		addAns[172] <= 26'd0;
		addAns[173] <= 26'd0;
		addAns[174] <= 26'd0;
		addAns[175] <= 26'd0;
		addAns[176] <= 26'd0;
		addAns[177] <= 26'd0;
		addAns[178] <= 26'd0;
		addAns[179] <= 26'd0;
		addAns[180] <= 26'd0;
		addAns[181] <= 26'd0;
		addAns[182] <= 26'd0;
		addAns[183] <= 26'd0;
		addAns[184] <= 26'd0;
		addAns[185] <= 26'd0;
		addAns[186] <= 26'd0;
		addAns[187] <= 26'd0;
		addAns[188] <= 26'd0;
		addAns[189] <= 26'd0;
		addAns[190] <= 26'd0;
		addAns[191] <= 26'd0;
		addAns[192] <= 26'd0;
		addAns[193] <= 26'd0;
		addAns[194] <= 26'd0;
		addAns[195] <= 26'd0;
		addAns[196] <= 26'd0;
		addAns[197] <= 26'd0;
		addAns[198] <= 26'd0;
		addAns[199] <= 26'd0;
		addAns[200] <= 26'd0;
		addAns[201] <= 26'd0;
		addAns[202] <= 26'd0;
		addAns[203] <= 26'd0;
		addAns[204] <= 26'd0;
		addAns[205] <= 26'd0;
		addAns[206] <= 26'd0;
		addAns[207] <= 26'd0;
		addAns[208] <= 26'd0;
		addAns[209] <= 26'd0;
		addAns[210] <= 26'd0;
		addAns[211] <= 26'd0;
		addAns[212] <= 26'd0;
		addAns[213] <= 26'd0;
		addAns[214] <= 26'd0;
		addAns[215] <= 26'd0;
		addAns[216] <= 26'd0;
		addAns[217] <= 26'd0;
		addAns[218] <= 26'd0;
		addAns[219] <= 26'd0;
		addAns[220] <= 26'd0;
		addAns[221] <= 26'd0;
		addAns[222] <= 26'd0;
		addAns[223] <= 26'd0;
		addAns[224] <= 26'd0;
		addAns[225] <= 26'd0;
		addAns[226] <= 26'd0;
		addAns[227] <= 26'd0;
		addAns[228] <= 26'd0;
		addAns[229] <= 26'd0;
		addAns[230] <= 26'd0;
		addAns[231] <= 26'd0;
		addAns[232] <= 26'd0;
		addAns[233] <= 26'd0;
		addAns[234] <= 26'd0;
		addAns[235] <= 26'd0;
		addAns[236] <= 26'd0;
		addAns[237] <= 26'd0;
		addAns[238] <= 26'd0;
		addAns[239] <= 26'd0;
		addAns[240] <= 26'd0;
		addAns[241] <= 26'd0;
		addAns[242] <= 26'd0;
		addAns[243] <= 26'd0;
		addAns[244] <= 26'd0;
		addAns[245] <= 26'd0;
		addAns[246] <= 26'd0;
		addAns[247] <= 26'd0;
		addAns[248] <= 26'd0;
		addAns[249] <= 26'd0;
		addAns[250] <= 26'd0;
		addAns[251] <= 26'd0;
		addAns[252] <= 26'd0;
		addAns[253] <= 26'd0;
		addAns[254] <= 26'd0;
		addAns[255] <= 26'd0;
		addAns[256] <= 26'd0;
		addAns[257] <= 26'd0;
		addAns[258] <= 26'd0;
		addAns[259] <= 26'd0;
		addAns[260] <= 26'd0;
		addAns[261] <= 26'd0;
		addAns[262] <= 26'd0;
		addAns[263] <= 26'd0;
		addAns[264] <= 26'd0;
		addAns[265] <= 26'd0;
		addAns[266] <= 26'd0;
		addAns[267] <= 26'd0;
		addAns[268] <= 26'd0;
		addAns[269] <= 26'd0;
		addAns[270] <= 26'd0;
		addAns[271] <= 26'd0;
		addAns[272] <= 26'd0;
		addAns[273] <= 26'd0;
		addAns[274] <= 26'd0;
		addAns[275] <= 26'd0;
		addAns[276] <= 26'd0;
		addAns[277] <= 26'd0;
		addAns[278] <= 26'd0;
		addAns[279] <= 26'd0;
		addAns[280] <= 26'd0;
		addAns[281] <= 26'd0;
		addAns[282] <= 26'd0;
		addAns[283] <= 26'd0;
		addAns[284] <= 26'd0;
		addAns[285] <= 26'd0;
		addAns[286] <= 26'd0;
		addAns[287] <= 26'd0;
		addAns[288] <= 26'd0;
		addAns[289] <= 26'd0;
		addAns[290] <= 26'd0;
		addAns[291] <= 26'd0;
		addAns[292] <= 26'd0;
		addAns[293] <= 26'd0;
		addAns[294] <= 26'd0;
		addAns[295] <= 26'd0;
		addAns[296] <= 26'd0;
		addAns[297] <= 26'd0;
		addAns[298] <= 26'd0;
		addAns[299] <= 26'd0;
		addAns[300] <= 26'd0;
		addAns[301] <= 26'd0;
		addAns[302] <= 26'd0;
		addAns[303] <= 26'd0;
		addAns[304] <= 26'd0;
		addAns[305] <= 26'd0;
		addAns[306] <= 26'd0;
		addAns[307] <= 26'd0;
		addAns[308] <= 26'd0;
		addAns[309] <= 26'd0;
		addAns[310] <= 26'd0;
		addAns[311] <= 26'd0;
		addAns[312] <= 26'd0;
		addAns[313] <= 26'd0;
		addAns[314] <= 26'd0;
		addAns[315] <= 26'd0;
		addAns[316] <= 26'd0;
		addAns[317] <= 26'd0;
		addAns[318] <= 26'd0;
		addAns[319] <= 26'd0;
		addAns[320] <= 26'd0;
		addAns[321] <= 26'd0;
		addAns[322] <= 26'd0;
		addAns[323] <= 26'd0;
		addAns[324] <= 26'd0;
		addAns[325] <= 26'd0;
		addAns[326] <= 26'd0;
		addAns[327] <= 26'd0;
		addAns[328] <= 26'd0;
		addAns[329] <= 26'd0;
		addAns[330] <= 26'd0;
		addAns[331] <= 26'd0;
		addAns[332] <= 26'd0;
		addAns[333] <= 26'd0;
		addAns[334] <= 26'd0;
		addAns[335] <= 26'd0;
		addAns[336] <= 26'd0;
		addAns[337] <= 26'd0;
		addAns[338] <= 26'd0;
		addAns[339] <= 26'd0;
		addAns[340] <= 26'd0;
		addAns[341] <= 26'd0;
		addAns[342] <= 26'd0;
		addAns[343] <= 26'd0;
		addAns[344] <= 26'd0;
		addAns[345] <= 26'd0;
		addAns[346] <= 26'd0;
		addAns[347] <= 26'd0;
		addAns[348] <= 26'd0;
		addAns[349] <= 26'd0;
		addAns[350] <= 26'd0;
		addAns[351] <= 26'd0;
		addAns[352] <= 26'd0;
		addAns[353] <= 26'd0;
		addAns[354] <= 26'd0;
		addAns[355] <= 26'd0;
		addAns[356] <= 26'd0;
		addAns[357] <= 26'd0;
		addAns[358] <= 26'd0;
		addAns[359] <= 26'd0;
		addAns[360] <= 26'd0;
		addAns[361] <= 26'd0;
		addAns[362] <= 26'd0;
		addAns[363] <= 26'd0;
		addAns[364] <= 26'd0;
		addAns[365] <= 26'd0;
		addAns[366] <= 26'd0;
		addAns[367] <= 26'd0;
		addAns[368] <= 26'd0;
		addAns[369] <= 26'd0;
		addAns[370] <= 26'd0;
		addAns[371] <= 26'd0;
		addAns[372] <= 26'd0;
		addAns[373] <= 26'd0;
		addAns[374] <= 26'd0;
		addAns[375] <= 26'd0;
		addAns[376] <= 26'd0;
		addAns[377] <= 26'd0;
		addAns[378] <= 26'd0;
		addAns[379] <= 26'd0;
		addAns[380] <= 26'd0;
		addAns[381] <= 26'd0;
		addAns[382] <= 26'd0;
		addAns[383] <= 26'd0;
		addAns[384] <= 26'd0;
		addAns[385] <= 26'd0;
		addAns[386] <= 26'd0;
		addAns[387] <= 26'd0;
		addAns[388] <= 26'd0;
		addAns[389] <= 26'd0;
		addAns[390] <= 26'd0;
		addAns[391] <= 26'd0;
	end else begin
		case(switchCounter)
			0: begin
				A1 <= A[0];
				A2 <= A[392];
				B1 <= B[0];
				B2 <= B[392];
			end
			1: begin
				A1 <= A[1];
				A2 <= A[393];
				B1 <= B[1];
				B2 <= B[393];
			end
			2: begin
				A1 <= A[2];
				A2 <= A[394];
				B1 <= B[2];
				B2 <= B[394];
			end
			3: begin
				A1 <= A[3];
				A2 <= A[395];
				B1 <= B[3];
				B2 <= B[395];
			end
			4: begin
				A1 <= A[4];
				A2 <= A[396];
				B1 <= B[4];
				B2 <= B[396];
			end
			5: begin
				A1 <= A[5];
				A2 <= A[397];
				B1 <= B[5];
				B2 <= B[397];
			end
			6: begin
				A1 <= A[6];
				A2 <= A[398];
				B1 <= B[6];
				B2 <= B[398];
			end
			7: begin
				A1 <= A[7];
				A2 <= A[399];
				B1 <= B[7];
				B2 <= B[399];
			end
			8: begin
				A1 <= A[8];
				A2 <= A[400];
				B1 <= B[8];
				B2 <= B[400];
			end
			9: begin
				A1 <= A[9];
				A2 <= A[401];
				B1 <= B[9];
				B2 <= B[401];
			end
			10: begin
				A1 <= A[10];
				A2 <= A[402];
				B1 <= B[10];
				B2 <= B[402];
			end
			11: begin
				A1 <= A[11];
				A2 <= A[403];
				B1 <= B[11];
				B2 <= B[403];
			end
			12: begin
				A1 <= A[12];
				A2 <= A[404];
				B1 <= B[12];
				B2 <= B[404];
			end
			13: begin
				A1 <= A[13];
				A2 <= A[405];
				B1 <= B[13];
				B2 <= B[405];
			end
			14: begin
				A1 <= A[14];
				A2 <= A[406];
				B1 <= B[14];
				B2 <= B[406];
			end
			15: begin
				A1 <= A[15];
				A2 <= A[407];
				B1 <= B[15];
				B2 <= B[407];
			end
			16: begin
				A1 <= A[16];
				A2 <= A[408];
				B1 <= B[16];
				B2 <= B[408];
			end
			17: begin
				A1 <= A[17];
				A2 <= A[409];
				B1 <= B[17];
				B2 <= B[409];
			end
			18: begin
				A1 <= A[18];
				A2 <= A[410];
				B1 <= B[18];
				B2 <= B[410];
			end
			19: begin
				A1 <= A[19];
				A2 <= A[411];
				B1 <= B[19];
				B2 <= B[411];
			end
			20: begin
				A1 <= A[20];
				A2 <= A[412];
				B1 <= B[20];
				B2 <= B[412];
			end
			21: begin
				A1 <= A[21];
				A2 <= A[413];
				B1 <= B[21];
				B2 <= B[413];
			end
			22: begin
				A1 <= A[22];
				A2 <= A[414];
				B1 <= B[22];
				B2 <= B[414];
			end
			23: begin
				A1 <= A[23];
				A2 <= A[415];
				B1 <= B[23];
				B2 <= B[415];
			end
			24: begin
				A1 <= A[24];
				A2 <= A[416];
				B1 <= B[24];
				B2 <= B[416];
			end
			25: begin
				A1 <= A[25];
				A2 <= A[417];
				B1 <= B[25];
				B2 <= B[417];
			end
			26: begin
				A1 <= A[26];
				A2 <= A[418];
				B1 <= B[26];
				B2 <= B[418];
			end
			27: begin
				A1 <= A[27];
				A2 <= A[419];
				B1 <= B[27];
				B2 <= B[419];
			end
			28: begin
				A1 <= A[28];
				A2 <= A[420];
				B1 <= B[28];
				B2 <= B[420];
			end
			29: begin
				A1 <= A[29];
				A2 <= A[421];
				B1 <= B[29];
				B2 <= B[421];
			end
			30: begin
				A1 <= A[30];
				A2 <= A[422];
				B1 <= B[30];
				B2 <= B[422];
			end
			31: begin
				A1 <= A[31];
				A2 <= A[423];
				B1 <= B[31];
				B2 <= B[423];
			end
			32: begin
				A1 <= A[32];
				A2 <= A[424];
				B1 <= B[32];
				B2 <= B[424];
			end
			33: begin
				A1 <= A[33];
				A2 <= A[425];
				B1 <= B[33];
				B2 <= B[425];
			end
			34: begin
				A1 <= A[34];
				A2 <= A[426];
				B1 <= B[34];
				B2 <= B[426];
			end
			35: begin
				A1 <= A[35];
				A2 <= A[427];
				B1 <= B[35];
				B2 <= B[427];
			end
			36: begin
				A1 <= A[36];
				A2 <= A[428];
				B1 <= B[36];
				B2 <= B[428];
			end
			37: begin
				A1 <= A[37];
				A2 <= A[429];
				B1 <= B[37];
				B2 <= B[429];
			end
			38: begin
				A1 <= A[38];
				A2 <= A[430];
				B1 <= B[38];
				B2 <= B[430];
			end
			39: begin
				A1 <= A[39];
				A2 <= A[431];
				B1 <= B[39];
				B2 <= B[431];
			end
			40: begin
				A1 <= A[40];
				A2 <= A[432];
				B1 <= B[40];
				B2 <= B[432];
			end
			41: begin
				A1 <= A[41];
				A2 <= A[433];
				B1 <= B[41];
				B2 <= B[433];
			end
			42: begin
				A1 <= A[42];
				A2 <= A[434];
				B1 <= B[42];
				B2 <= B[434];
			end
			43: begin
				A1 <= A[43];
				A2 <= A[435];
				B1 <= B[43];
				B2 <= B[435];
			end
			44: begin
				A1 <= A[44];
				A2 <= A[436];
				B1 <= B[44];
				B2 <= B[436];
			end
			45: begin
				A1 <= A[45];
				A2 <= A[437];
				B1 <= B[45];
				B2 <= B[437];
			end
			46: begin
				A1 <= A[46];
				A2 <= A[438];
				B1 <= B[46];
				B2 <= B[438];
			end
			47: begin
				A1 <= A[47];
				A2 <= A[439];
				B1 <= B[47];
				B2 <= B[439];
			end
			48: begin
				A1 <= A[48];
				A2 <= A[440];
				B1 <= B[48];
				B2 <= B[440];
			end
			49: begin
				A1 <= A[49];
				A2 <= A[441];
				B1 <= B[49];
				B2 <= B[441];
			end
			50: begin
				A1 <= A[50];
				A2 <= A[442];
				B1 <= B[50];
				B2 <= B[442];
			end
			51: begin
				A1 <= A[51];
				A2 <= A[443];
				B1 <= B[51];
				B2 <= B[443];
			end
			52: begin
				A1 <= A[52];
				A2 <= A[444];
				B1 <= B[52];
				B2 <= B[444];
			end
			53: begin
				A1 <= A[53];
				A2 <= A[445];
				B1 <= B[53];
				B2 <= B[445];
			end
			54: begin
				A1 <= A[54];
				A2 <= A[446];
				B1 <= B[54];
				B2 <= B[446];
			end
			55: begin
				A1 <= A[55];
				A2 <= A[447];
				B1 <= B[55];
				B2 <= B[447];
			end
			56: begin
				A1 <= A[56];
				A2 <= A[448];
				B1 <= B[56];
				B2 <= B[448];
			end
			57: begin
				A1 <= A[57];
				A2 <= A[449];
				B1 <= B[57];
				B2 <= B[449];
			end
			58: begin
				A1 <= A[58];
				A2 <= A[450];
				B1 <= B[58];
				B2 <= B[450];
			end
			59: begin
				A1 <= A[59];
				A2 <= A[451];
				B1 <= B[59];
				B2 <= B[451];
			end
			60: begin
				A1 <= A[60];
				A2 <= A[452];
				B1 <= B[60];
				B2 <= B[452];
			end
			61: begin
				A1 <= A[61];
				A2 <= A[453];
				B1 <= B[61];
				B2 <= B[453];
			end
			62: begin
				A1 <= A[62];
				A2 <= A[454];
				B1 <= B[62];
				B2 <= B[454];
			end
			63: begin
				A1 <= A[63];
				A2 <= A[455];
				B1 <= B[63];
				B2 <= B[455];
			end
			64: begin
				A1 <= A[64];
				A2 <= A[456];
				B1 <= B[64];
				B2 <= B[456];
			end
			65: begin
				A1 <= A[65];
				A2 <= A[457];
				B1 <= B[65];
				B2 <= B[457];
			end
			66: begin
				A1 <= A[66];
				A2 <= A[458];
				B1 <= B[66];
				B2 <= B[458];
			end
			67: begin
				A1 <= A[67];
				A2 <= A[459];
				B1 <= B[67];
				B2 <= B[459];
			end
			68: begin
				A1 <= A[68];
				A2 <= A[460];
				B1 <= B[68];
				B2 <= B[460];
			end
			69: begin
				A1 <= A[69];
				A2 <= A[461];
				B1 <= B[69];
				B2 <= B[461];
			end
			70: begin
				A1 <= A[70];
				A2 <= A[462];
				B1 <= B[70];
				B2 <= B[462];
			end
			71: begin
				A1 <= A[71];
				A2 <= A[463];
				B1 <= B[71];
				B2 <= B[463];
			end
			72: begin
				A1 <= A[72];
				A2 <= A[464];
				B1 <= B[72];
				B2 <= B[464];
			end
			73: begin
				A1 <= A[73];
				A2 <= A[465];
				B1 <= B[73];
				B2 <= B[465];
			end
			74: begin
				A1 <= A[74];
				A2 <= A[466];
				B1 <= B[74];
				B2 <= B[466];
			end
			75: begin
				A1 <= A[75];
				A2 <= A[467];
				B1 <= B[75];
				B2 <= B[467];
			end
			76: begin
				A1 <= A[76];
				A2 <= A[468];
				B1 <= B[76];
				B2 <= B[468];
			end
			77: begin
				A1 <= A[77];
				A2 <= A[469];
				B1 <= B[77];
				B2 <= B[469];
			end
			78: begin
				A1 <= A[78];
				A2 <= A[470];
				B1 <= B[78];
				B2 <= B[470];
			end
			79: begin
				A1 <= A[79];
				A2 <= A[471];
				B1 <= B[79];
				B2 <= B[471];
			end
			80: begin
				A1 <= A[80];
				A2 <= A[472];
				B1 <= B[80];
				B2 <= B[472];
			end
			81: begin
				A1 <= A[81];
				A2 <= A[473];
				B1 <= B[81];
				B2 <= B[473];
			end
			82: begin
				A1 <= A[82];
				A2 <= A[474];
				B1 <= B[82];
				B2 <= B[474];
			end
			83: begin
				A1 <= A[83];
				A2 <= A[475];
				B1 <= B[83];
				B2 <= B[475];
			end
			84: begin
				A1 <= A[84];
				A2 <= A[476];
				B1 <= B[84];
				B2 <= B[476];
			end
			85: begin
				A1 <= A[85];
				A2 <= A[477];
				B1 <= B[85];
				B2 <= B[477];
			end
			86: begin
				A1 <= A[86];
				A2 <= A[478];
				B1 <= B[86];
				B2 <= B[478];
			end
			87: begin
				A1 <= A[87];
				A2 <= A[479];
				B1 <= B[87];
				B2 <= B[479];
			end
			88: begin
				A1 <= A[88];
				A2 <= A[480];
				B1 <= B[88];
				B2 <= B[480];
			end
			89: begin
				A1 <= A[89];
				A2 <= A[481];
				B1 <= B[89];
				B2 <= B[481];
			end
			90: begin
				A1 <= A[90];
				A2 <= A[482];
				B1 <= B[90];
				B2 <= B[482];
			end
			91: begin
				A1 <= A[91];
				A2 <= A[483];
				B1 <= B[91];
				B2 <= B[483];
			end
			92: begin
				A1 <= A[92];
				A2 <= A[484];
				B1 <= B[92];
				B2 <= B[484];
			end
			93: begin
				A1 <= A[93];
				A2 <= A[485];
				B1 <= B[93];
				B2 <= B[485];
			end
			94: begin
				A1 <= A[94];
				A2 <= A[486];
				B1 <= B[94];
				B2 <= B[486];
			end
			95: begin
				A1 <= A[95];
				A2 <= A[487];
				B1 <= B[95];
				B2 <= B[487];
			end
			96: begin
				A1 <= A[96];
				A2 <= A[488];
				B1 <= B[96];
				B2 <= B[488];
			end
			97: begin
				A1 <= A[97];
				A2 <= A[489];
				B1 <= B[97];
				B2 <= B[489];
			end
			98: begin
				A1 <= A[98];
				A2 <= A[490];
				B1 <= B[98];
				B2 <= B[490];
			end
			99: begin
				A1 <= A[99];
				A2 <= A[491];
				B1 <= B[99];
				B2 <= B[491];
			end
			100: begin
				A1 <= A[100];
				A2 <= A[492];
				B1 <= B[100];
				B2 <= B[492];
			end
			101: begin
				A1 <= A[101];
				A2 <= A[493];
				B1 <= B[101];
				B2 <= B[493];
			end
			102: begin
				A1 <= A[102];
				A2 <= A[494];
				B1 <= B[102];
				B2 <= B[494];
			end
			103: begin
				A1 <= A[103];
				A2 <= A[495];
				B1 <= B[103];
				B2 <= B[495];
			end
			104: begin
				A1 <= A[104];
				A2 <= A[496];
				B1 <= B[104];
				B2 <= B[496];
			end
			105: begin
				A1 <= A[105];
				A2 <= A[497];
				B1 <= B[105];
				B2 <= B[497];
			end
			106: begin
				A1 <= A[106];
				A2 <= A[498];
				B1 <= B[106];
				B2 <= B[498];
			end
			107: begin
				A1 <= A[107];
				A2 <= A[499];
				B1 <= B[107];
				B2 <= B[499];
			end
			108: begin
				A1 <= A[108];
				A2 <= A[500];
				B1 <= B[108];
				B2 <= B[500];
			end
			109: begin
				A1 <= A[109];
				A2 <= A[501];
				B1 <= B[109];
				B2 <= B[501];
			end
			110: begin
				A1 <= A[110];
				A2 <= A[502];
				B1 <= B[110];
				B2 <= B[502];
			end
			111: begin
				A1 <= A[111];
				A2 <= A[503];
				B1 <= B[111];
				B2 <= B[503];
			end
			112: begin
				A1 <= A[112];
				A2 <= A[504];
				B1 <= B[112];
				B2 <= B[504];
			end
			113: begin
				A1 <= A[113];
				A2 <= A[505];
				B1 <= B[113];
				B2 <= B[505];
			end
			114: begin
				A1 <= A[114];
				A2 <= A[506];
				B1 <= B[114];
				B2 <= B[506];
			end
			115: begin
				A1 <= A[115];
				A2 <= A[507];
				B1 <= B[115];
				B2 <= B[507];
			end
			116: begin
				A1 <= A[116];
				A2 <= A[508];
				B1 <= B[116];
				B2 <= B[508];
			end
			117: begin
				A1 <= A[117];
				A2 <= A[509];
				B1 <= B[117];
				B2 <= B[509];
			end
			118: begin
				A1 <= A[118];
				A2 <= A[510];
				B1 <= B[118];
				B2 <= B[510];
			end
			119: begin
				A1 <= A[119];
				A2 <= A[511];
				B1 <= B[119];
				B2 <= B[511];
			end
			120: begin
				A1 <= A[120];
				A2 <= A[512];
				B1 <= B[120];
				B2 <= B[512];
			end
			121: begin
				A1 <= A[121];
				A2 <= A[513];
				B1 <= B[121];
				B2 <= B[513];
			end
			122: begin
				A1 <= A[122];
				A2 <= A[514];
				B1 <= B[122];
				B2 <= B[514];
			end
			123: begin
				A1 <= A[123];
				A2 <= A[515];
				B1 <= B[123];
				B2 <= B[515];
			end
			124: begin
				A1 <= A[124];
				A2 <= A[516];
				B1 <= B[124];
				B2 <= B[516];
			end
			125: begin
				A1 <= A[125];
				A2 <= A[517];
				B1 <= B[125];
				B2 <= B[517];
			end
			126: begin
				A1 <= A[126];
				A2 <= A[518];
				B1 <= B[126];
				B2 <= B[518];
			end
			127: begin
				A1 <= A[127];
				A2 <= A[519];
				B1 <= B[127];
				B2 <= B[519];
			end
			128: begin
				A1 <= A[128];
				A2 <= A[520];
				B1 <= B[128];
				B2 <= B[520];
			end
			129: begin
				A1 <= A[129];
				A2 <= A[521];
				B1 <= B[129];
				B2 <= B[521];
			end
			130: begin
				A1 <= A[130];
				A2 <= A[522];
				B1 <= B[130];
				B2 <= B[522];
			end
			131: begin
				A1 <= A[131];
				A2 <= A[523];
				B1 <= B[131];
				B2 <= B[523];
			end
			132: begin
				A1 <= A[132];
				A2 <= A[524];
				B1 <= B[132];
				B2 <= B[524];
			end
			133: begin
				A1 <= A[133];
				A2 <= A[525];
				B1 <= B[133];
				B2 <= B[525];
			end
			134: begin
				A1 <= A[134];
				A2 <= A[526];
				B1 <= B[134];
				B2 <= B[526];
			end
			135: begin
				A1 <= A[135];
				A2 <= A[527];
				B1 <= B[135];
				B2 <= B[527];
			end
			136: begin
				A1 <= A[136];
				A2 <= A[528];
				B1 <= B[136];
				B2 <= B[528];
			end
			137: begin
				A1 <= A[137];
				A2 <= A[529];
				B1 <= B[137];
				B2 <= B[529];
			end
			138: begin
				A1 <= A[138];
				A2 <= A[530];
				B1 <= B[138];
				B2 <= B[530];
			end
			139: begin
				A1 <= A[139];
				A2 <= A[531];
				B1 <= B[139];
				B2 <= B[531];
			end
			140: begin
				A1 <= A[140];
				A2 <= A[532];
				B1 <= B[140];
				B2 <= B[532];
			end
			141: begin
				A1 <= A[141];
				A2 <= A[533];
				B1 <= B[141];
				B2 <= B[533];
			end
			142: begin
				A1 <= A[142];
				A2 <= A[534];
				B1 <= B[142];
				B2 <= B[534];
			end
			143: begin
				A1 <= A[143];
				A2 <= A[535];
				B1 <= B[143];
				B2 <= B[535];
			end
			144: begin
				A1 <= A[144];
				A2 <= A[536];
				B1 <= B[144];
				B2 <= B[536];
			end
			145: begin
				A1 <= A[145];
				A2 <= A[537];
				B1 <= B[145];
				B2 <= B[537];
			end
			146: begin
				A1 <= A[146];
				A2 <= A[538];
				B1 <= B[146];
				B2 <= B[538];
			end
			147: begin
				A1 <= A[147];
				A2 <= A[539];
				B1 <= B[147];
				B2 <= B[539];
			end
			148: begin
				A1 <= A[148];
				A2 <= A[540];
				B1 <= B[148];
				B2 <= B[540];
			end
			149: begin
				A1 <= A[149];
				A2 <= A[541];
				B1 <= B[149];
				B2 <= B[541];
			end
			150: begin
				A1 <= A[150];
				A2 <= A[542];
				B1 <= B[150];
				B2 <= B[542];
			end
			151: begin
				A1 <= A[151];
				A2 <= A[543];
				B1 <= B[151];
				B2 <= B[543];
			end
			152: begin
				A1 <= A[152];
				A2 <= A[544];
				B1 <= B[152];
				B2 <= B[544];
			end
			153: begin
				A1 <= A[153];
				A2 <= A[545];
				B1 <= B[153];
				B2 <= B[545];
			end
			154: begin
				A1 <= A[154];
				A2 <= A[546];
				B1 <= B[154];
				B2 <= B[546];
			end
			155: begin
				A1 <= A[155];
				A2 <= A[547];
				B1 <= B[155];
				B2 <= B[547];
			end
			156: begin
				A1 <= A[156];
				A2 <= A[548];
				B1 <= B[156];
				B2 <= B[548];
			end
			157: begin
				A1 <= A[157];
				A2 <= A[549];
				B1 <= B[157];
				B2 <= B[549];
			end
			158: begin
				A1 <= A[158];
				A2 <= A[550];
				B1 <= B[158];
				B2 <= B[550];
			end
			159: begin
				A1 <= A[159];
				A2 <= A[551];
				B1 <= B[159];
				B2 <= B[551];
			end
			160: begin
				A1 <= A[160];
				A2 <= A[552];
				B1 <= B[160];
				B2 <= B[552];
			end
			161: begin
				A1 <= A[161];
				A2 <= A[553];
				B1 <= B[161];
				B2 <= B[553];
			end
			162: begin
				A1 <= A[162];
				A2 <= A[554];
				B1 <= B[162];
				B2 <= B[554];
			end
			163: begin
				A1 <= A[163];
				A2 <= A[555];
				B1 <= B[163];
				B2 <= B[555];
			end
			164: begin
				A1 <= A[164];
				A2 <= A[556];
				B1 <= B[164];
				B2 <= B[556];
			end
			165: begin
				A1 <= A[165];
				A2 <= A[557];
				B1 <= B[165];
				B2 <= B[557];
			end
			166: begin
				A1 <= A[166];
				A2 <= A[558];
				B1 <= B[166];
				B2 <= B[558];
			end
			167: begin
				A1 <= A[167];
				A2 <= A[559];
				B1 <= B[167];
				B2 <= B[559];
			end
			168: begin
				A1 <= A[168];
				A2 <= A[560];
				B1 <= B[168];
				B2 <= B[560];
			end
			169: begin
				A1 <= A[169];
				A2 <= A[561];
				B1 <= B[169];
				B2 <= B[561];
			end
			170: begin
				A1 <= A[170];
				A2 <= A[562];
				B1 <= B[170];
				B2 <= B[562];
			end
			171: begin
				A1 <= A[171];
				A2 <= A[563];
				B1 <= B[171];
				B2 <= B[563];
			end
			172: begin
				A1 <= A[172];
				A2 <= A[564];
				B1 <= B[172];
				B2 <= B[564];
			end
			173: begin
				A1 <= A[173];
				A2 <= A[565];
				B1 <= B[173];
				B2 <= B[565];
			end
			174: begin
				A1 <= A[174];
				A2 <= A[566];
				B1 <= B[174];
				B2 <= B[566];
			end
			175: begin
				A1 <= A[175];
				A2 <= A[567];
				B1 <= B[175];
				B2 <= B[567];
			end
			176: begin
				A1 <= A[176];
				A2 <= A[568];
				B1 <= B[176];
				B2 <= B[568];
			end
			177: begin
				A1 <= A[177];
				A2 <= A[569];
				B1 <= B[177];
				B2 <= B[569];
			end
			178: begin
				A1 <= A[178];
				A2 <= A[570];
				B1 <= B[178];
				B2 <= B[570];
			end
			179: begin
				A1 <= A[179];
				A2 <= A[571];
				B1 <= B[179];
				B2 <= B[571];
			end
			180: begin
				A1 <= A[180];
				A2 <= A[572];
				B1 <= B[180];
				B2 <= B[572];
			end
			181: begin
				A1 <= A[181];
				A2 <= A[573];
				B1 <= B[181];
				B2 <= B[573];
			end
			182: begin
				A1 <= A[182];
				A2 <= A[574];
				B1 <= B[182];
				B2 <= B[574];
			end
			183: begin
				A1 <= A[183];
				A2 <= A[575];
				B1 <= B[183];
				B2 <= B[575];
			end
			184: begin
				A1 <= A[184];
				A2 <= A[576];
				B1 <= B[184];
				B2 <= B[576];
			end
			185: begin
				A1 <= A[185];
				A2 <= A[577];
				B1 <= B[185];
				B2 <= B[577];
			end
			186: begin
				A1 <= A[186];
				A2 <= A[578];
				B1 <= B[186];
				B2 <= B[578];
			end
			187: begin
				A1 <= A[187];
				A2 <= A[579];
				B1 <= B[187];
				B2 <= B[579];
			end
			188: begin
				A1 <= A[188];
				A2 <= A[580];
				B1 <= B[188];
				B2 <= B[580];
			end
			189: begin
				A1 <= A[189];
				A2 <= A[581];
				B1 <= B[189];
				B2 <= B[581];
			end
			190: begin
				A1 <= A[190];
				A2 <= A[582];
				B1 <= B[190];
				B2 <= B[582];
			end
			191: begin
				A1 <= A[191];
				A2 <= A[583];
				B1 <= B[191];
				B2 <= B[583];
			end
			192: begin
				A1 <= A[192];
				A2 <= A[584];
				B1 <= B[192];
				B2 <= B[584];
			end
			193: begin
				A1 <= A[193];
				A2 <= A[585];
				B1 <= B[193];
				B2 <= B[585];
			end
			194: begin
				A1 <= A[194];
				A2 <= A[586];
				B1 <= B[194];
				B2 <= B[586];
			end
			195: begin
				A1 <= A[195];
				A2 <= A[587];
				B1 <= B[195];
				B2 <= B[587];
			end
			196: begin
				A1 <= A[196];
				A2 <= A[588];
				B1 <= B[196];
				B2 <= B[588];
			end
			197: begin
				A1 <= A[197];
				A2 <= A[589];
				B1 <= B[197];
				B2 <= B[589];
			end
			198: begin
				A1 <= A[198];
				A2 <= A[590];
				B1 <= B[198];
				B2 <= B[590];
			end
			199: begin
				A1 <= A[199];
				A2 <= A[591];
				B1 <= B[199];
				B2 <= B[591];
			end
			200: begin
				A1 <= A[200];
				A2 <= A[592];
				B1 <= B[200];
				B2 <= B[592];
			end
			201: begin
				A1 <= A[201];
				A2 <= A[593];
				B1 <= B[201];
				B2 <= B[593];
			end
			202: begin
				A1 <= A[202];
				A2 <= A[594];
				B1 <= B[202];
				B2 <= B[594];
			end
			203: begin
				A1 <= A[203];
				A2 <= A[595];
				B1 <= B[203];
				B2 <= B[595];
			end
			204: begin
				A1 <= A[204];
				A2 <= A[596];
				B1 <= B[204];
				B2 <= B[596];
			end
			205: begin
				A1 <= A[205];
				A2 <= A[597];
				B1 <= B[205];
				B2 <= B[597];
			end
			206: begin
				A1 <= A[206];
				A2 <= A[598];
				B1 <= B[206];
				B2 <= B[598];
			end
			207: begin
				A1 <= A[207];
				A2 <= A[599];
				B1 <= B[207];
				B2 <= B[599];
			end
			208: begin
				A1 <= A[208];
				A2 <= A[600];
				B1 <= B[208];
				B2 <= B[600];
			end
			209: begin
				A1 <= A[209];
				A2 <= A[601];
				B1 <= B[209];
				B2 <= B[601];
			end
			210: begin
				A1 <= A[210];
				A2 <= A[602];
				B1 <= B[210];
				B2 <= B[602];
			end
			211: begin
				A1 <= A[211];
				A2 <= A[603];
				B1 <= B[211];
				B2 <= B[603];
			end
			212: begin
				A1 <= A[212];
				A2 <= A[604];
				B1 <= B[212];
				B2 <= B[604];
			end
			213: begin
				A1 <= A[213];
				A2 <= A[605];
				B1 <= B[213];
				B2 <= B[605];
			end
			214: begin
				A1 <= A[214];
				A2 <= A[606];
				B1 <= B[214];
				B2 <= B[606];
			end
			215: begin
				A1 <= A[215];
				A2 <= A[607];
				B1 <= B[215];
				B2 <= B[607];
			end
			216: begin
				A1 <= A[216];
				A2 <= A[608];
				B1 <= B[216];
				B2 <= B[608];
			end
			217: begin
				A1 <= A[217];
				A2 <= A[609];
				B1 <= B[217];
				B2 <= B[609];
			end
			218: begin
				A1 <= A[218];
				A2 <= A[610];
				B1 <= B[218];
				B2 <= B[610];
			end
			219: begin
				A1 <= A[219];
				A2 <= A[611];
				B1 <= B[219];
				B2 <= B[611];
			end
			220: begin
				A1 <= A[220];
				A2 <= A[612];
				B1 <= B[220];
				B2 <= B[612];
			end
			221: begin
				A1 <= A[221];
				A2 <= A[613];
				B1 <= B[221];
				B2 <= B[613];
			end
			222: begin
				A1 <= A[222];
				A2 <= A[614];
				B1 <= B[222];
				B2 <= B[614];
			end
			223: begin
				A1 <= A[223];
				A2 <= A[615];
				B1 <= B[223];
				B2 <= B[615];
			end
			224: begin
				A1 <= A[224];
				A2 <= A[616];
				B1 <= B[224];
				B2 <= B[616];
			end
			225: begin
				A1 <= A[225];
				A2 <= A[617];
				B1 <= B[225];
				B2 <= B[617];
			end
			226: begin
				A1 <= A[226];
				A2 <= A[618];
				B1 <= B[226];
				B2 <= B[618];
			end
			227: begin
				A1 <= A[227];
				A2 <= A[619];
				B1 <= B[227];
				B2 <= B[619];
			end
			228: begin
				A1 <= A[228];
				A2 <= A[620];
				B1 <= B[228];
				B2 <= B[620];
			end
			229: begin
				A1 <= A[229];
				A2 <= A[621];
				B1 <= B[229];
				B2 <= B[621];
			end
			230: begin
				A1 <= A[230];
				A2 <= A[622];
				B1 <= B[230];
				B2 <= B[622];
			end
			231: begin
				A1 <= A[231];
				A2 <= A[623];
				B1 <= B[231];
				B2 <= B[623];
			end
			232: begin
				A1 <= A[232];
				A2 <= A[624];
				B1 <= B[232];
				B2 <= B[624];
			end
			233: begin
				A1 <= A[233];
				A2 <= A[625];
				B1 <= B[233];
				B2 <= B[625];
			end
			234: begin
				A1 <= A[234];
				A2 <= A[626];
				B1 <= B[234];
				B2 <= B[626];
			end
			235: begin
				A1 <= A[235];
				A2 <= A[627];
				B1 <= B[235];
				B2 <= B[627];
			end
			236: begin
				A1 <= A[236];
				A2 <= A[628];
				B1 <= B[236];
				B2 <= B[628];
			end
			237: begin
				A1 <= A[237];
				A2 <= A[629];
				B1 <= B[237];
				B2 <= B[629];
			end
			238: begin
				A1 <= A[238];
				A2 <= A[630];
				B1 <= B[238];
				B2 <= B[630];
			end
			239: begin
				A1 <= A[239];
				A2 <= A[631];
				B1 <= B[239];
				B2 <= B[631];
			end
			240: begin
				A1 <= A[240];
				A2 <= A[632];
				B1 <= B[240];
				B2 <= B[632];
			end
			241: begin
				A1 <= A[241];
				A2 <= A[633];
				B1 <= B[241];
				B2 <= B[633];
			end
			242: begin
				A1 <= A[242];
				A2 <= A[634];
				B1 <= B[242];
				B2 <= B[634];
			end
			243: begin
				A1 <= A[243];
				A2 <= A[635];
				B1 <= B[243];
				B2 <= B[635];
			end
			244: begin
				A1 <= A[244];
				A2 <= A[636];
				B1 <= B[244];
				B2 <= B[636];
			end
			245: begin
				A1 <= A[245];
				A2 <= A[637];
				B1 <= B[245];
				B2 <= B[637];
			end
			246: begin
				A1 <= A[246];
				A2 <= A[638];
				B1 <= B[246];
				B2 <= B[638];
			end
			247: begin
				A1 <= A[247];
				A2 <= A[639];
				B1 <= B[247];
				B2 <= B[639];
			end
			248: begin
				A1 <= A[248];
				A2 <= A[640];
				B1 <= B[248];
				B2 <= B[640];
			end
			249: begin
				A1 <= A[249];
				A2 <= A[641];
				B1 <= B[249];
				B2 <= B[641];
			end
			250: begin
				A1 <= A[250];
				A2 <= A[642];
				B1 <= B[250];
				B2 <= B[642];
			end
			251: begin
				A1 <= A[251];
				A2 <= A[643];
				B1 <= B[251];
				B2 <= B[643];
			end
			252: begin
				A1 <= A[252];
				A2 <= A[644];
				B1 <= B[252];
				B2 <= B[644];
			end
			253: begin
				A1 <= A[253];
				A2 <= A[645];
				B1 <= B[253];
				B2 <= B[645];
			end
			254: begin
				A1 <= A[254];
				A2 <= A[646];
				B1 <= B[254];
				B2 <= B[646];
			end
			255: begin
				A1 <= A[255];
				A2 <= A[647];
				B1 <= B[255];
				B2 <= B[647];
			end
			256: begin
				A1 <= A[256];
				A2 <= A[648];
				B1 <= B[256];
				B2 <= B[648];
			end
			257: begin
				A1 <= A[257];
				A2 <= A[649];
				B1 <= B[257];
				B2 <= B[649];
			end
			258: begin
				A1 <= A[258];
				A2 <= A[650];
				B1 <= B[258];
				B2 <= B[650];
			end
			259: begin
				A1 <= A[259];
				A2 <= A[651];
				B1 <= B[259];
				B2 <= B[651];
			end
			260: begin
				A1 <= A[260];
				A2 <= A[652];
				B1 <= B[260];
				B2 <= B[652];
			end
			261: begin
				A1 <= A[261];
				A2 <= A[653];
				B1 <= B[261];
				B2 <= B[653];
			end
			262: begin
				A1 <= A[262];
				A2 <= A[654];
				B1 <= B[262];
				B2 <= B[654];
			end
			263: begin
				A1 <= A[263];
				A2 <= A[655];
				B1 <= B[263];
				B2 <= B[655];
			end
			264: begin
				A1 <= A[264];
				A2 <= A[656];
				B1 <= B[264];
				B2 <= B[656];
			end
			265: begin
				A1 <= A[265];
				A2 <= A[657];
				B1 <= B[265];
				B2 <= B[657];
			end
			266: begin
				A1 <= A[266];
				A2 <= A[658];
				B1 <= B[266];
				B2 <= B[658];
			end
			267: begin
				A1 <= A[267];
				A2 <= A[659];
				B1 <= B[267];
				B2 <= B[659];
			end
			268: begin
				A1 <= A[268];
				A2 <= A[660];
				B1 <= B[268];
				B2 <= B[660];
			end
			269: begin
				A1 <= A[269];
				A2 <= A[661];
				B1 <= B[269];
				B2 <= B[661];
			end
			270: begin
				A1 <= A[270];
				A2 <= A[662];
				B1 <= B[270];
				B2 <= B[662];
			end
			271: begin
				A1 <= A[271];
				A2 <= A[663];
				B1 <= B[271];
				B2 <= B[663];
			end
			272: begin
				A1 <= A[272];
				A2 <= A[664];
				B1 <= B[272];
				B2 <= B[664];
			end
			273: begin
				A1 <= A[273];
				A2 <= A[665];
				B1 <= B[273];
				B2 <= B[665];
			end
			274: begin
				A1 <= A[274];
				A2 <= A[666];
				B1 <= B[274];
				B2 <= B[666];
			end
			275: begin
				A1 <= A[275];
				A2 <= A[667];
				B1 <= B[275];
				B2 <= B[667];
			end
			276: begin
				A1 <= A[276];
				A2 <= A[668];
				B1 <= B[276];
				B2 <= B[668];
			end
			277: begin
				A1 <= A[277];
				A2 <= A[669];
				B1 <= B[277];
				B2 <= B[669];
			end
			278: begin
				A1 <= A[278];
				A2 <= A[670];
				B1 <= B[278];
				B2 <= B[670];
			end
			279: begin
				A1 <= A[279];
				A2 <= A[671];
				B1 <= B[279];
				B2 <= B[671];
			end
			280: begin
				A1 <= A[280];
				A2 <= A[672];
				B1 <= B[280];
				B2 <= B[672];
			end
			281: begin
				A1 <= A[281];
				A2 <= A[673];
				B1 <= B[281];
				B2 <= B[673];
			end
			282: begin
				A1 <= A[282];
				A2 <= A[674];
				B1 <= B[282];
				B2 <= B[674];
			end
			283: begin
				A1 <= A[283];
				A2 <= A[675];
				B1 <= B[283];
				B2 <= B[675];
			end
			284: begin
				A1 <= A[284];
				A2 <= A[676];
				B1 <= B[284];
				B2 <= B[676];
			end
			285: begin
				A1 <= A[285];
				A2 <= A[677];
				B1 <= B[285];
				B2 <= B[677];
			end
			286: begin
				A1 <= A[286];
				A2 <= A[678];
				B1 <= B[286];
				B2 <= B[678];
			end
			287: begin
				A1 <= A[287];
				A2 <= A[679];
				B1 <= B[287];
				B2 <= B[679];
			end
			288: begin
				A1 <= A[288];
				A2 <= A[680];
				B1 <= B[288];
				B2 <= B[680];
			end
			289: begin
				A1 <= A[289];
				A2 <= A[681];
				B1 <= B[289];
				B2 <= B[681];
			end
			290: begin
				A1 <= A[290];
				A2 <= A[682];
				B1 <= B[290];
				B2 <= B[682];
			end
			291: begin
				A1 <= A[291];
				A2 <= A[683];
				B1 <= B[291];
				B2 <= B[683];
			end
			292: begin
				A1 <= A[292];
				A2 <= A[684];
				B1 <= B[292];
				B2 <= B[684];
			end
			293: begin
				A1 <= A[293];
				A2 <= A[685];
				B1 <= B[293];
				B2 <= B[685];
			end
			294: begin
				A1 <= A[294];
				A2 <= A[686];
				B1 <= B[294];
				B2 <= B[686];
			end
			295: begin
				A1 <= A[295];
				A2 <= A[687];
				B1 <= B[295];
				B2 <= B[687];
			end
			296: begin
				A1 <= A[296];
				A2 <= A[688];
				B1 <= B[296];
				B2 <= B[688];
			end
			297: begin
				A1 <= A[297];
				A2 <= A[689];
				B1 <= B[297];
				B2 <= B[689];
			end
			298: begin
				A1 <= A[298];
				A2 <= A[690];
				B1 <= B[298];
				B2 <= B[690];
			end
			299: begin
				A1 <= A[299];
				A2 <= A[691];
				B1 <= B[299];
				B2 <= B[691];
			end
			300: begin
				A1 <= A[300];
				A2 <= A[692];
				B1 <= B[300];
				B2 <= B[692];
			end
			301: begin
				A1 <= A[301];
				A2 <= A[693];
				B1 <= B[301];
				B2 <= B[693];
			end
			302: begin
				A1 <= A[302];
				A2 <= A[694];
				B1 <= B[302];
				B2 <= B[694];
			end
			303: begin
				A1 <= A[303];
				A2 <= A[695];
				B1 <= B[303];
				B2 <= B[695];
			end
			304: begin
				A1 <= A[304];
				A2 <= A[696];
				B1 <= B[304];
				B2 <= B[696];
			end
			305: begin
				A1 <= A[305];
				A2 <= A[697];
				B1 <= B[305];
				B2 <= B[697];
			end
			306: begin
				A1 <= A[306];
				A2 <= A[698];
				B1 <= B[306];
				B2 <= B[698];
			end
			307: begin
				A1 <= A[307];
				A2 <= A[699];
				B1 <= B[307];
				B2 <= B[699];
			end
			308: begin
				A1 <= A[308];
				A2 <= A[700];
				B1 <= B[308];
				B2 <= B[700];
			end
			309: begin
				A1 <= A[309];
				A2 <= A[701];
				B1 <= B[309];
				B2 <= B[701];
			end
			310: begin
				A1 <= A[310];
				A2 <= A[702];
				B1 <= B[310];
				B2 <= B[702];
			end
			311: begin
				A1 <= A[311];
				A2 <= A[703];
				B1 <= B[311];
				B2 <= B[703];
			end
			312: begin
				A1 <= A[312];
				A2 <= A[704];
				B1 <= B[312];
				B2 <= B[704];
			end
			313: begin
				A1 <= A[313];
				A2 <= A[705];
				B1 <= B[313];
				B2 <= B[705];
			end
			314: begin
				A1 <= A[314];
				A2 <= A[706];
				B1 <= B[314];
				B2 <= B[706];
			end
			315: begin
				A1 <= A[315];
				A2 <= A[707];
				B1 <= B[315];
				B2 <= B[707];
			end
			316: begin
				A1 <= A[316];
				A2 <= A[708];
				B1 <= B[316];
				B2 <= B[708];
			end
			317: begin
				A1 <= A[317];
				A2 <= A[709];
				B1 <= B[317];
				B2 <= B[709];
			end
			318: begin
				A1 <= A[318];
				A2 <= A[710];
				B1 <= B[318];
				B2 <= B[710];
			end
			319: begin
				A1 <= A[319];
				A2 <= A[711];
				B1 <= B[319];
				B2 <= B[711];
			end
			320: begin
				A1 <= A[320];
				A2 <= A[712];
				B1 <= B[320];
				B2 <= B[712];
			end
			321: begin
				A1 <= A[321];
				A2 <= A[713];
				B1 <= B[321];
				B2 <= B[713];
			end
			322: begin
				A1 <= A[322];
				A2 <= A[714];
				B1 <= B[322];
				B2 <= B[714];
			end
			323: begin
				A1 <= A[323];
				A2 <= A[715];
				B1 <= B[323];
				B2 <= B[715];
			end
			324: begin
				A1 <= A[324];
				A2 <= A[716];
				B1 <= B[324];
				B2 <= B[716];
			end
			325: begin
				A1 <= A[325];
				A2 <= A[717];
				B1 <= B[325];
				B2 <= B[717];
			end
			326: begin
				A1 <= A[326];
				A2 <= A[718];
				B1 <= B[326];
				B2 <= B[718];
			end
			327: begin
				A1 <= A[327];
				A2 <= A[719];
				B1 <= B[327];
				B2 <= B[719];
			end
			328: begin
				A1 <= A[328];
				A2 <= A[720];
				B1 <= B[328];
				B2 <= B[720];
			end
			329: begin
				A1 <= A[329];
				A2 <= A[721];
				B1 <= B[329];
				B2 <= B[721];
			end
			330: begin
				A1 <= A[330];
				A2 <= A[722];
				B1 <= B[330];
				B2 <= B[722];
			end
			331: begin
				A1 <= A[331];
				A2 <= A[723];
				B1 <= B[331];
				B2 <= B[723];
			end
			332: begin
				A1 <= A[332];
				A2 <= A[724];
				B1 <= B[332];
				B2 <= B[724];
			end
			333: begin
				A1 <= A[333];
				A2 <= A[725];
				B1 <= B[333];
				B2 <= B[725];
			end
			334: begin
				A1 <= A[334];
				A2 <= A[726];
				B1 <= B[334];
				B2 <= B[726];
			end
			335: begin
				A1 <= A[335];
				A2 <= A[727];
				B1 <= B[335];
				B2 <= B[727];
			end
			336: begin
				A1 <= A[336];
				A2 <= A[728];
				B1 <= B[336];
				B2 <= B[728];
			end
			337: begin
				A1 <= A[337];
				A2 <= A[729];
				B1 <= B[337];
				B2 <= B[729];
			end
			338: begin
				A1 <= A[338];
				A2 <= A[730];
				B1 <= B[338];
				B2 <= B[730];
			end
			339: begin
				A1 <= A[339];
				A2 <= A[731];
				B1 <= B[339];
				B2 <= B[731];
			end
			340: begin
				A1 <= A[340];
				A2 <= A[732];
				B1 <= B[340];
				B2 <= B[732];
			end
			341: begin
				A1 <= A[341];
				A2 <= A[733];
				B1 <= B[341];
				B2 <= B[733];
			end
			342: begin
				A1 <= A[342];
				A2 <= A[734];
				B1 <= B[342];
				B2 <= B[734];
			end
			343: begin
				A1 <= A[343];
				A2 <= A[735];
				B1 <= B[343];
				B2 <= B[735];
			end
			344: begin
				A1 <= A[344];
				A2 <= A[736];
				B1 <= B[344];
				B2 <= B[736];
			end
			345: begin
				A1 <= A[345];
				A2 <= A[737];
				B1 <= B[345];
				B2 <= B[737];
			end
			346: begin
				A1 <= A[346];
				A2 <= A[738];
				B1 <= B[346];
				B2 <= B[738];
			end
			347: begin
				A1 <= A[347];
				A2 <= A[739];
				B1 <= B[347];
				B2 <= B[739];
			end
			348: begin
				A1 <= A[348];
				A2 <= A[740];
				B1 <= B[348];
				B2 <= B[740];
			end
			349: begin
				A1 <= A[349];
				A2 <= A[741];
				B1 <= B[349];
				B2 <= B[741];
			end
			350: begin
				A1 <= A[350];
				A2 <= A[742];
				B1 <= B[350];
				B2 <= B[742];
			end
			351: begin
				A1 <= A[351];
				A2 <= A[743];
				B1 <= B[351];
				B2 <= B[743];
			end
			352: begin
				A1 <= A[352];
				A2 <= A[744];
				B1 <= B[352];
				B2 <= B[744];
			end
			353: begin
				A1 <= A[353];
				A2 <= A[745];
				B1 <= B[353];
				B2 <= B[745];
			end
			354: begin
				A1 <= A[354];
				A2 <= A[746];
				B1 <= B[354];
				B2 <= B[746];
			end
			355: begin
				A1 <= A[355];
				A2 <= A[747];
				B1 <= B[355];
				B2 <= B[747];
			end
			356: begin
				A1 <= A[356];
				A2 <= A[748];
				B1 <= B[356];
				B2 <= B[748];
			end
			357: begin
				A1 <= A[357];
				A2 <= A[749];
				B1 <= B[357];
				B2 <= B[749];
			end
			358: begin
				A1 <= A[358];
				A2 <= A[750];
				B1 <= B[358];
				B2 <= B[750];
			end
			359: begin
				A1 <= A[359];
				A2 <= A[751];
				B1 <= B[359];
				B2 <= B[751];
			end
			360: begin
				A1 <= A[360];
				A2 <= A[752];
				B1 <= B[360];
				B2 <= B[752];
			end
			361: begin
				A1 <= A[361];
				A2 <= A[753];
				B1 <= B[361];
				B2 <= B[753];
			end
			362: begin
				A1 <= A[362];
				A2 <= A[754];
				B1 <= B[362];
				B2 <= B[754];
			end
			363: begin
				A1 <= A[363];
				A2 <= A[755];
				B1 <= B[363];
				B2 <= B[755];
			end
			364: begin
				A1 <= A[364];
				A2 <= A[756];
				B1 <= B[364];
				B2 <= B[756];
			end
			365: begin
				A1 <= A[365];
				A2 <= A[757];
				B1 <= B[365];
				B2 <= B[757];
			end
			366: begin
				A1 <= A[366];
				A2 <= A[758];
				B1 <= B[366];
				B2 <= B[758];
			end
			367: begin
				A1 <= A[367];
				A2 <= A[759];
				B1 <= B[367];
				B2 <= B[759];
			end
			368: begin
				A1 <= A[368];
				A2 <= A[760];
				B1 <= B[368];
				B2 <= B[760];
			end
			369: begin
				A1 <= A[369];
				A2 <= A[761];
				B1 <= B[369];
				B2 <= B[761];
			end
			370: begin
				A1 <= A[370];
				A2 <= A[762];
				B1 <= B[370];
				B2 <= B[762];
			end
			371: begin
				A1 <= A[371];
				A2 <= A[763];
				B1 <= B[371];
				B2 <= B[763];
			end
			372: begin
				A1 <= A[372];
				A2 <= A[764];
				B1 <= B[372];
				B2 <= B[764];
			end
			373: begin
				A1 <= A[373];
				A2 <= A[765];
				B1 <= B[373];
				B2 <= B[765];
			end
			374: begin
				A1 <= A[374];
				A2 <= A[766];
				B1 <= B[374];
				B2 <= B[766];
			end
			375: begin
				A1 <= A[375];
				A2 <= A[767];
				B1 <= B[375];
				B2 <= B[767];
			end
			376: begin
				A1 <= A[376];
				A2 <= A[768];
				B1 <= B[376];
				B2 <= B[768];
			end
			377: begin
				A1 <= A[377];
				A2 <= A[769];
				B1 <= B[377];
				B2 <= B[769];
			end
			378: begin
				A1 <= A[378];
				A2 <= A[770];
				B1 <= B[378];
				B2 <= B[770];
			end
			379: begin
				A1 <= A[379];
				A2 <= A[771];
				B1 <= B[379];
				B2 <= B[771];
			end
			380: begin
				A1 <= A[380];
				A2 <= A[772];
				B1 <= B[380];
				B2 <= B[772];
			end
			381: begin
				A1 <= A[381];
				A2 <= A[773];
				B1 <= B[381];
				B2 <= B[773];
			end
			382: begin
				A1 <= A[382];
				A2 <= A[774];
				B1 <= B[382];
				B2 <= B[774];
			end
			383: begin
				A1 <= A[383];
				A2 <= A[775];
				B1 <= B[383];
				B2 <= B[775];
			end
			384: begin
				A1 <= A[384];
				A2 <= A[776];
				B1 <= B[384];
				B2 <= B[776];
			end
			385: begin
				A1 <= A[385];
				A2 <= A[777];
				B1 <= B[385];
				B2 <= B[777];
			end
			386: begin
				A1 <= A[386];
				A2 <= A[778];
				B1 <= B[386];
				B2 <= B[778];
			end
			387: begin
				A1 <= A[387];
				A2 <= A[779];
				B1 <= B[387];
				B2 <= B[779];
			end
			388: begin
				A1 <= A[388];
				A2 <= A[780];
				B1 <= B[388];
				B2 <= B[780];
			end
			389: begin
				A1 <= A[389];
				A2 <= A[781];
				B1 <= B[389];
				B2 <= B[781];
			end
			390: begin
				A1 <= A[390];
				A2 <= A[782];
				B1 <= B[390];
				B2 <= B[782];
			end
			391: begin
				A1 <= A[391];
				A2 <= A[783];
				B1 <= B[391];
				B2 <= B[783];
			end
			default: begin
				A1 <= A1;
				A2 <= A2;
				B1 <= B1;
				B2 <= B2;
			end
		endcase

		if(switchCounter >= 32'd7 && switchCounter <= 32'd398) begin
			addInput[0] <= FPMAns1;
			addInput[1] <= FPMAns2;
		end
		if(switchCounter >= 32'd10 && switchCounter <= 32'd401) begin
			addAns[switchCounter - 32'd10] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd399 && switchCounter <= 32'd594) begin
			addInput[0] <= addAns[(switchCounter - 32'd399) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd399) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd402 && switchCounter <= 32'd597) begin
			addAns[switchCounter - 32'd402] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd595 && switchCounter <= 32'd692) begin
			addInput[0] <= addAns[(switchCounter - 32'd595) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd595) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd598 && switchCounter <= 32'd695) begin
			addAns[switchCounter - 32'd598] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd693 && switchCounter <= 32'd741) begin
			addInput[0] <= addAns[(switchCounter - 32'd693) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd693) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd696 && switchCounter <= 32'd744) begin
			addAns[switchCounter - 32'd696] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd742 && switchCounter <= 32'd765) begin
			addInput[0] <= addAns[(switchCounter - 32'd742) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd742) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd745 && switchCounter <= 32'd768) begin
			addAns[switchCounter - 32'd745] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd766 && switchCounter <= 32'd777) begin
			addInput[0] <= addAns[(switchCounter - 32'd766) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd766) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd769 && switchCounter <= 32'd780) begin
			addAns[switchCounter - 32'd769] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd778 && switchCounter <= 32'd783) begin
			addInput[0] <= addAns[(switchCounter - 32'd778) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd778) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd781 && switchCounter <= 32'd786) begin
			addAns[switchCounter - 32'd781] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter >= 32'd786 && switchCounter <= 32'd788) begin
			addInput[0] <= addAns[(switchCounter - 32'd786) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd786) << 1'd1) + 32'd1];
		end
		if(switchCounter >= 32'd789 && switchCounter <= 32'd791) begin
			addAns[switchCounter - 32'd789] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter == 32'd792) begin
			addInput[0] <= addAns[(switchCounter - 32'd792) << 1'd1];
 			addInput[1] <= addAns[((switchCounter - 32'd792) << 1'd1) + 32'd1];
		end
		if(switchCounter == 32'd795) begin
			addAns[switchCounter - 32'd795] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter == 32'd796) begin
			addInput[0] <= addAns[2];
 			addInput[1] <= addAns[48];
		end
		if(switchCounter == 32'd799) begin
			addAns[1] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		if(switchCounter == 32'd802) begin
			addInput[0] <= addAns[0];
 			addInput[1] <= addAns[1];
		end
		if(switchCounter == 32'd805) begin
			addAns[0] <= FPAAns;
			$display("%d %b.%b", switchCounter, FPAAns[25:18],FPAAns[17:0]);
		end
		switchCounter <= switchCounter + 32'd1;
	end
end
endmodule
