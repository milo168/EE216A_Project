module Image_Classifier(
input clk,
input GlobalReset,
input Input_Valid,
input [18:0] Wgt_0_0,
input [18:0] Wgt_0_1,
input [18:0] Wgt_0_2,
input [18:0] Wgt_0_3,
input [18:0] Wgt_0_4,
input [18:0] Wgt_0_5,
input [18:0] Wgt_0_6,
input [18:0] Wgt_0_7,
input [18:0] Wgt_0_8,
input [18:0] Wgt_0_9,
input [18:0] Wgt_0_10,
input [18:0] Wgt_0_11,
input [18:0] Wgt_0_12,
input [18:0] Wgt_0_13,
input [18:0] Wgt_0_14,
input [18:0] Wgt_0_15,
input [18:0] Wgt_0_16,
input [18:0] Wgt_0_17,
input [18:0] Wgt_0_18,
input [18:0] Wgt_0_19,
input [18:0] Wgt_0_20,
input [18:0] Wgt_0_21,
input [18:0] Wgt_0_22,
input [18:0] Wgt_0_23,
input [18:0] Wgt_0_24,
input [18:0] Wgt_0_25,
input [18:0] Wgt_0_26,
input [18:0] Wgt_0_27,
input [18:0] Wgt_0_28,
input [18:0] Wgt_0_29,
input [18:0] Wgt_0_30,
input [18:0] Wgt_0_31,
input [18:0] Wgt_0_32,
input [18:0] Wgt_0_33,
input [18:0] Wgt_0_34,
input [18:0] Wgt_0_35,
input [18:0] Wgt_0_36,
input [18:0] Wgt_0_37,
input [18:0] Wgt_0_38,
input [18:0] Wgt_0_39,
input [18:0] Wgt_0_40,
input [18:0] Wgt_0_41,
input [18:0] Wgt_0_42,
input [18:0] Wgt_0_43,
input [18:0] Wgt_0_44,
input [18:0] Wgt_0_45,
input [18:0] Wgt_0_46,
input [18:0] Wgt_0_47,
input [18:0] Wgt_0_48,
input [18:0] Wgt_0_49,
input [18:0] Wgt_0_50,
input [18:0] Wgt_0_51,
input [18:0] Wgt_0_52,
input [18:0] Wgt_0_53,
input [18:0] Wgt_0_54,
input [18:0] Wgt_0_55,
input [18:0] Wgt_0_56,
input [18:0] Wgt_0_57,
input [18:0] Wgt_0_58,
input [18:0] Wgt_0_59,
input [18:0] Wgt_0_60,
input [18:0] Wgt_0_61,
input [18:0] Wgt_0_62,
input [18:0] Wgt_0_63,
input [18:0] Wgt_0_64,
input [18:0] Wgt_0_65,
input [18:0] Wgt_0_66,
input [18:0] Wgt_0_67,
input [18:0] Wgt_0_68,
input [18:0] Wgt_0_69,
input [18:0] Wgt_0_70,
input [18:0] Wgt_0_71,
input [18:0] Wgt_0_72,
input [18:0] Wgt_0_73,
input [18:0] Wgt_0_74,
input [18:0] Wgt_0_75,
input [18:0] Wgt_0_76,
input [18:0] Wgt_0_77,
input [18:0] Wgt_0_78,
input [18:0] Wgt_0_79,
input [18:0] Wgt_0_80,
input [18:0] Wgt_0_81,
input [18:0] Wgt_0_82,
input [18:0] Wgt_0_83,
input [18:0] Wgt_0_84,
input [18:0] Wgt_0_85,
input [18:0] Wgt_0_86,
input [18:0] Wgt_0_87,
input [18:0] Wgt_0_88,
input [18:0] Wgt_0_89,
input [18:0] Wgt_0_90,
input [18:0] Wgt_0_91,
input [18:0] Wgt_0_92,
input [18:0] Wgt_0_93,
input [18:0] Wgt_0_94,
input [18:0] Wgt_0_95,
input [18:0] Wgt_0_96,
input [18:0] Wgt_0_97,
input [18:0] Wgt_0_98,
input [18:0] Wgt_0_99,
input [18:0] Wgt_0_100,
input [18:0] Wgt_0_101,
input [18:0] Wgt_0_102,
input [18:0] Wgt_0_103,
input [18:0] Wgt_0_104,
input [18:0] Wgt_0_105,
input [18:0] Wgt_0_106,
input [18:0] Wgt_0_107,
input [18:0] Wgt_0_108,
input [18:0] Wgt_0_109,
input [18:0] Wgt_0_110,
input [18:0] Wgt_0_111,
input [18:0] Wgt_0_112,
input [18:0] Wgt_0_113,
input [18:0] Wgt_0_114,
input [18:0] Wgt_0_115,
input [18:0] Wgt_0_116,
input [18:0] Wgt_0_117,
input [18:0] Wgt_0_118,
input [18:0] Wgt_0_119,
input [18:0] Wgt_0_120,
input [18:0] Wgt_0_121,
input [18:0] Wgt_0_122,
input [18:0] Wgt_0_123,
input [18:0] Wgt_0_124,
input [18:0] Wgt_0_125,
input [18:0] Wgt_0_126,
input [18:0] Wgt_0_127,
input [18:0] Wgt_0_128,
input [18:0] Wgt_0_129,
input [18:0] Wgt_0_130,
input [18:0] Wgt_0_131,
input [18:0] Wgt_0_132,
input [18:0] Wgt_0_133,
input [18:0] Wgt_0_134,
input [18:0] Wgt_0_135,
input [18:0] Wgt_0_136,
input [18:0] Wgt_0_137,
input [18:0] Wgt_0_138,
input [18:0] Wgt_0_139,
input [18:0] Wgt_0_140,
input [18:0] Wgt_0_141,
input [18:0] Wgt_0_142,
input [18:0] Wgt_0_143,
input [18:0] Wgt_0_144,
input [18:0] Wgt_0_145,
input [18:0] Wgt_0_146,
input [18:0] Wgt_0_147,
input [18:0] Wgt_0_148,
input [18:0] Wgt_0_149,
input [18:0] Wgt_0_150,
input [18:0] Wgt_0_151,
input [18:0] Wgt_0_152,
input [18:0] Wgt_0_153,
input [18:0] Wgt_0_154,
input [18:0] Wgt_0_155,
input [18:0] Wgt_0_156,
input [18:0] Wgt_0_157,
input [18:0] Wgt_0_158,
input [18:0] Wgt_0_159,
input [18:0] Wgt_0_160,
input [18:0] Wgt_0_161,
input [18:0] Wgt_0_162,
input [18:0] Wgt_0_163,
input [18:0] Wgt_0_164,
input [18:0] Wgt_0_165,
input [18:0] Wgt_0_166,
input [18:0] Wgt_0_167,
input [18:0] Wgt_0_168,
input [18:0] Wgt_0_169,
input [18:0] Wgt_0_170,
input [18:0] Wgt_0_171,
input [18:0] Wgt_0_172,
input [18:0] Wgt_0_173,
input [18:0] Wgt_0_174,
input [18:0] Wgt_0_175,
input [18:0] Wgt_0_176,
input [18:0] Wgt_0_177,
input [18:0] Wgt_0_178,
input [18:0] Wgt_0_179,
input [18:0] Wgt_0_180,
input [18:0] Wgt_0_181,
input [18:0] Wgt_0_182,
input [18:0] Wgt_0_183,
input [18:0] Wgt_0_184,
input [18:0] Wgt_0_185,
input [18:0] Wgt_0_186,
input [18:0] Wgt_0_187,
input [18:0] Wgt_0_188,
input [18:0] Wgt_0_189,
input [18:0] Wgt_0_190,
input [18:0] Wgt_0_191,
input [18:0] Wgt_0_192,
input [18:0] Wgt_0_193,
input [18:0] Wgt_0_194,
input [18:0] Wgt_0_195,
input [18:0] Wgt_0_196,
input [18:0] Wgt_0_197,
input [18:0] Wgt_0_198,
input [18:0] Wgt_0_199,
input [18:0] Wgt_0_200,
input [18:0] Wgt_0_201,
input [18:0] Wgt_0_202,
input [18:0] Wgt_0_203,
input [18:0] Wgt_0_204,
input [18:0] Wgt_0_205,
input [18:0] Wgt_0_206,
input [18:0] Wgt_0_207,
input [18:0] Wgt_0_208,
input [18:0] Wgt_0_209,
input [18:0] Wgt_0_210,
input [18:0] Wgt_0_211,
input [18:0] Wgt_0_212,
input [18:0] Wgt_0_213,
input [18:0] Wgt_0_214,
input [18:0] Wgt_0_215,
input [18:0] Wgt_0_216,
input [18:0] Wgt_0_217,
input [18:0] Wgt_0_218,
input [18:0] Wgt_0_219,
input [18:0] Wgt_0_220,
input [18:0] Wgt_0_221,
input [18:0] Wgt_0_222,
input [18:0] Wgt_0_223,
input [18:0] Wgt_0_224,
input [18:0] Wgt_0_225,
input [18:0] Wgt_0_226,
input [18:0] Wgt_0_227,
input [18:0] Wgt_0_228,
input [18:0] Wgt_0_229,
input [18:0] Wgt_0_230,
input [18:0] Wgt_0_231,
input [18:0] Wgt_0_232,
input [18:0] Wgt_0_233,
input [18:0] Wgt_0_234,
input [18:0] Wgt_0_235,
input [18:0] Wgt_0_236,
input [18:0] Wgt_0_237,
input [18:0] Wgt_0_238,
input [18:0] Wgt_0_239,
input [18:0] Wgt_0_240,
input [18:0] Wgt_0_241,
input [18:0] Wgt_0_242,
input [18:0] Wgt_0_243,
input [18:0] Wgt_0_244,
input [18:0] Wgt_0_245,
input [18:0] Wgt_0_246,
input [18:0] Wgt_0_247,
input [18:0] Wgt_0_248,
input [18:0] Wgt_0_249,
input [18:0] Wgt_0_250,
input [18:0] Wgt_0_251,
input [18:0] Wgt_0_252,
input [18:0] Wgt_0_253,
input [18:0] Wgt_0_254,
input [18:0] Wgt_0_255,
input [18:0] Wgt_0_256,
input [18:0] Wgt_0_257,
input [18:0] Wgt_0_258,
input [18:0] Wgt_0_259,
input [18:0] Wgt_0_260,
input [18:0] Wgt_0_261,
input [18:0] Wgt_0_262,
input [18:0] Wgt_0_263,
input [18:0] Wgt_0_264,
input [18:0] Wgt_0_265,
input [18:0] Wgt_0_266,
input [18:0] Wgt_0_267,
input [18:0] Wgt_0_268,
input [18:0] Wgt_0_269,
input [18:0] Wgt_0_270,
input [18:0] Wgt_0_271,
input [18:0] Wgt_0_272,
input [18:0] Wgt_0_273,
input [18:0] Wgt_0_274,
input [18:0] Wgt_0_275,
input [18:0] Wgt_0_276,
input [18:0] Wgt_0_277,
input [18:0] Wgt_0_278,
input [18:0] Wgt_0_279,
input [18:0] Wgt_0_280,
input [18:0] Wgt_0_281,
input [18:0] Wgt_0_282,
input [18:0] Wgt_0_283,
input [18:0] Wgt_0_284,
input [18:0] Wgt_0_285,
input [18:0] Wgt_0_286,
input [18:0] Wgt_0_287,
input [18:0] Wgt_0_288,
input [18:0] Wgt_0_289,
input [18:0] Wgt_0_290,
input [18:0] Wgt_0_291,
input [18:0] Wgt_0_292,
input [18:0] Wgt_0_293,
input [18:0] Wgt_0_294,
input [18:0] Wgt_0_295,
input [18:0] Wgt_0_296,
input [18:0] Wgt_0_297,
input [18:0] Wgt_0_298,
input [18:0] Wgt_0_299,
input [18:0] Wgt_0_300,
input [18:0] Wgt_0_301,
input [18:0] Wgt_0_302,
input [18:0] Wgt_0_303,
input [18:0] Wgt_0_304,
input [18:0] Wgt_0_305,
input [18:0] Wgt_0_306,
input [18:0] Wgt_0_307,
input [18:0] Wgt_0_308,
input [18:0] Wgt_0_309,
input [18:0] Wgt_0_310,
input [18:0] Wgt_0_311,
input [18:0] Wgt_0_312,
input [18:0] Wgt_0_313,
input [18:0] Wgt_0_314,
input [18:0] Wgt_0_315,
input [18:0] Wgt_0_316,
input [18:0] Wgt_0_317,
input [18:0] Wgt_0_318,
input [18:0] Wgt_0_319,
input [18:0] Wgt_0_320,
input [18:0] Wgt_0_321,
input [18:0] Wgt_0_322,
input [18:0] Wgt_0_323,
input [18:0] Wgt_0_324,
input [18:0] Wgt_0_325,
input [18:0] Wgt_0_326,
input [18:0] Wgt_0_327,
input [18:0] Wgt_0_328,
input [18:0] Wgt_0_329,
input [18:0] Wgt_0_330,
input [18:0] Wgt_0_331,
input [18:0] Wgt_0_332,
input [18:0] Wgt_0_333,
input [18:0] Wgt_0_334,
input [18:0] Wgt_0_335,
input [18:0] Wgt_0_336,
input [18:0] Wgt_0_337,
input [18:0] Wgt_0_338,
input [18:0] Wgt_0_339,
input [18:0] Wgt_0_340,
input [18:0] Wgt_0_341,
input [18:0] Wgt_0_342,
input [18:0] Wgt_0_343,
input [18:0] Wgt_0_344,
input [18:0] Wgt_0_345,
input [18:0] Wgt_0_346,
input [18:0] Wgt_0_347,
input [18:0] Wgt_0_348,
input [18:0] Wgt_0_349,
input [18:0] Wgt_0_350,
input [18:0] Wgt_0_351,
input [18:0] Wgt_0_352,
input [18:0] Wgt_0_353,
input [18:0] Wgt_0_354,
input [18:0] Wgt_0_355,
input [18:0] Wgt_0_356,
input [18:0] Wgt_0_357,
input [18:0] Wgt_0_358,
input [18:0] Wgt_0_359,
input [18:0] Wgt_0_360,
input [18:0] Wgt_0_361,
input [18:0] Wgt_0_362,
input [18:0] Wgt_0_363,
input [18:0] Wgt_0_364,
input [18:0] Wgt_0_365,
input [18:0] Wgt_0_366,
input [18:0] Wgt_0_367,
input [18:0] Wgt_0_368,
input [18:0] Wgt_0_369,
input [18:0] Wgt_0_370,
input [18:0] Wgt_0_371,
input [18:0] Wgt_0_372,
input [18:0] Wgt_0_373,
input [18:0] Wgt_0_374,
input [18:0] Wgt_0_375,
input [18:0] Wgt_0_376,
input [18:0] Wgt_0_377,
input [18:0] Wgt_0_378,
input [18:0] Wgt_0_379,
input [18:0] Wgt_0_380,
input [18:0] Wgt_0_381,
input [18:0] Wgt_0_382,
input [18:0] Wgt_0_383,
input [18:0] Wgt_0_384,
input [18:0] Wgt_0_385,
input [18:0] Wgt_0_386,
input [18:0] Wgt_0_387,
input [18:0] Wgt_0_388,
input [18:0] Wgt_0_389,
input [18:0] Wgt_0_390,
input [18:0] Wgt_0_391,
input [18:0] Wgt_0_392,
input [18:0] Wgt_0_393,
input [18:0] Wgt_0_394,
input [18:0] Wgt_0_395,
input [18:0] Wgt_0_396,
input [18:0] Wgt_0_397,
input [18:0] Wgt_0_398,
input [18:0] Wgt_0_399,
input [18:0] Wgt_0_400,
input [18:0] Wgt_0_401,
input [18:0] Wgt_0_402,
input [18:0] Wgt_0_403,
input [18:0] Wgt_0_404,
input [18:0] Wgt_0_405,
input [18:0] Wgt_0_406,
input [18:0] Wgt_0_407,
input [18:0] Wgt_0_408,
input [18:0] Wgt_0_409,
input [18:0] Wgt_0_410,
input [18:0] Wgt_0_411,
input [18:0] Wgt_0_412,
input [18:0] Wgt_0_413,
input [18:0] Wgt_0_414,
input [18:0] Wgt_0_415,
input [18:0] Wgt_0_416,
input [18:0] Wgt_0_417,
input [18:0] Wgt_0_418,
input [18:0] Wgt_0_419,
input [18:0] Wgt_0_420,
input [18:0] Wgt_0_421,
input [18:0] Wgt_0_422,
input [18:0] Wgt_0_423,
input [18:0] Wgt_0_424,
input [18:0] Wgt_0_425,
input [18:0] Wgt_0_426,
input [18:0] Wgt_0_427,
input [18:0] Wgt_0_428,
input [18:0] Wgt_0_429,
input [18:0] Wgt_0_430,
input [18:0] Wgt_0_431,
input [18:0] Wgt_0_432,
input [18:0] Wgt_0_433,
input [18:0] Wgt_0_434,
input [18:0] Wgt_0_435,
input [18:0] Wgt_0_436,
input [18:0] Wgt_0_437,
input [18:0] Wgt_0_438,
input [18:0] Wgt_0_439,
input [18:0] Wgt_0_440,
input [18:0] Wgt_0_441,
input [18:0] Wgt_0_442,
input [18:0] Wgt_0_443,
input [18:0] Wgt_0_444,
input [18:0] Wgt_0_445,
input [18:0] Wgt_0_446,
input [18:0] Wgt_0_447,
input [18:0] Wgt_0_448,
input [18:0] Wgt_0_449,
input [18:0] Wgt_0_450,
input [18:0] Wgt_0_451,
input [18:0] Wgt_0_452,
input [18:0] Wgt_0_453,
input [18:0] Wgt_0_454,
input [18:0] Wgt_0_455,
input [18:0] Wgt_0_456,
input [18:0] Wgt_0_457,
input [18:0] Wgt_0_458,
input [18:0] Wgt_0_459,
input [18:0] Wgt_0_460,
input [18:0] Wgt_0_461,
input [18:0] Wgt_0_462,
input [18:0] Wgt_0_463,
input [18:0] Wgt_0_464,
input [18:0] Wgt_0_465,
input [18:0] Wgt_0_466,
input [18:0] Wgt_0_467,
input [18:0] Wgt_0_468,
input [18:0] Wgt_0_469,
input [18:0] Wgt_0_470,
input [18:0] Wgt_0_471,
input [18:0] Wgt_0_472,
input [18:0] Wgt_0_473,
input [18:0] Wgt_0_474,
input [18:0] Wgt_0_475,
input [18:0] Wgt_0_476,
input [18:0] Wgt_0_477,
input [18:0] Wgt_0_478,
input [18:0] Wgt_0_479,
input [18:0] Wgt_0_480,
input [18:0] Wgt_0_481,
input [18:0] Wgt_0_482,
input [18:0] Wgt_0_483,
input [18:0] Wgt_0_484,
input [18:0] Wgt_0_485,
input [18:0] Wgt_0_486,
input [18:0] Wgt_0_487,
input [18:0] Wgt_0_488,
input [18:0] Wgt_0_489,
input [18:0] Wgt_0_490,
input [18:0] Wgt_0_491,
input [18:0] Wgt_0_492,
input [18:0] Wgt_0_493,
input [18:0] Wgt_0_494,
input [18:0] Wgt_0_495,
input [18:0] Wgt_0_496,
input [18:0] Wgt_0_497,
input [18:0] Wgt_0_498,
input [18:0] Wgt_0_499,
input [18:0] Wgt_0_500,
input [18:0] Wgt_0_501,
input [18:0] Wgt_0_502,
input [18:0] Wgt_0_503,
input [18:0] Wgt_0_504,
input [18:0] Wgt_0_505,
input [18:0] Wgt_0_506,
input [18:0] Wgt_0_507,
input [18:0] Wgt_0_508,
input [18:0] Wgt_0_509,
input [18:0] Wgt_0_510,
input [18:0] Wgt_0_511,
input [18:0] Wgt_0_512,
input [18:0] Wgt_0_513,
input [18:0] Wgt_0_514,
input [18:0] Wgt_0_515,
input [18:0] Wgt_0_516,
input [18:0] Wgt_0_517,
input [18:0] Wgt_0_518,
input [18:0] Wgt_0_519,
input [18:0] Wgt_0_520,
input [18:0] Wgt_0_521,
input [18:0] Wgt_0_522,
input [18:0] Wgt_0_523,
input [18:0] Wgt_0_524,
input [18:0] Wgt_0_525,
input [18:0] Wgt_0_526,
input [18:0] Wgt_0_527,
input [18:0] Wgt_0_528,
input [18:0] Wgt_0_529,
input [18:0] Wgt_0_530,
input [18:0] Wgt_0_531,
input [18:0] Wgt_0_532,
input [18:0] Wgt_0_533,
input [18:0] Wgt_0_534,
input [18:0] Wgt_0_535,
input [18:0] Wgt_0_536,
input [18:0] Wgt_0_537,
input [18:0] Wgt_0_538,
input [18:0] Wgt_0_539,
input [18:0] Wgt_0_540,
input [18:0] Wgt_0_541,
input [18:0] Wgt_0_542,
input [18:0] Wgt_0_543,
input [18:0] Wgt_0_544,
input [18:0] Wgt_0_545,
input [18:0] Wgt_0_546,
input [18:0] Wgt_0_547,
input [18:0] Wgt_0_548,
input [18:0] Wgt_0_549,
input [18:0] Wgt_0_550,
input [18:0] Wgt_0_551,
input [18:0] Wgt_0_552,
input [18:0] Wgt_0_553,
input [18:0] Wgt_0_554,
input [18:0] Wgt_0_555,
input [18:0] Wgt_0_556,
input [18:0] Wgt_0_557,
input [18:0] Wgt_0_558,
input [18:0] Wgt_0_559,
input [18:0] Wgt_0_560,
input [18:0] Wgt_0_561,
input [18:0] Wgt_0_562,
input [18:0] Wgt_0_563,
input [18:0] Wgt_0_564,
input [18:0] Wgt_0_565,
input [18:0] Wgt_0_566,
input [18:0] Wgt_0_567,
input [18:0] Wgt_0_568,
input [18:0] Wgt_0_569,
input [18:0] Wgt_0_570,
input [18:0] Wgt_0_571,
input [18:0] Wgt_0_572,
input [18:0] Wgt_0_573,
input [18:0] Wgt_0_574,
input [18:0] Wgt_0_575,
input [18:0] Wgt_0_576,
input [18:0] Wgt_0_577,
input [18:0] Wgt_0_578,
input [18:0] Wgt_0_579,
input [18:0] Wgt_0_580,
input [18:0] Wgt_0_581,
input [18:0] Wgt_0_582,
input [18:0] Wgt_0_583,
input [18:0] Wgt_0_584,
input [18:0] Wgt_0_585,
input [18:0] Wgt_0_586,
input [18:0] Wgt_0_587,
input [18:0] Wgt_0_588,
input [18:0] Wgt_0_589,
input [18:0] Wgt_0_590,
input [18:0] Wgt_0_591,
input [18:0] Wgt_0_592,
input [18:0] Wgt_0_593,
input [18:0] Wgt_0_594,
input [18:0] Wgt_0_595,
input [18:0] Wgt_0_596,
input [18:0] Wgt_0_597,
input [18:0] Wgt_0_598,
input [18:0] Wgt_0_599,
input [18:0] Wgt_0_600,
input [18:0] Wgt_0_601,
input [18:0] Wgt_0_602,
input [18:0] Wgt_0_603,
input [18:0] Wgt_0_604,
input [18:0] Wgt_0_605,
input [18:0] Wgt_0_606,
input [18:0] Wgt_0_607,
input [18:0] Wgt_0_608,
input [18:0] Wgt_0_609,
input [18:0] Wgt_0_610,
input [18:0] Wgt_0_611,
input [18:0] Wgt_0_612,
input [18:0] Wgt_0_613,
input [18:0] Wgt_0_614,
input [18:0] Wgt_0_615,
input [18:0] Wgt_0_616,
input [18:0] Wgt_0_617,
input [18:0] Wgt_0_618,
input [18:0] Wgt_0_619,
input [18:0] Wgt_0_620,
input [18:0] Wgt_0_621,
input [18:0] Wgt_0_622,
input [18:0] Wgt_0_623,
input [18:0] Wgt_0_624,
input [18:0] Wgt_0_625,
input [18:0] Wgt_0_626,
input [18:0] Wgt_0_627,
input [18:0] Wgt_0_628,
input [18:0] Wgt_0_629,
input [18:0] Wgt_0_630,
input [18:0] Wgt_0_631,
input [18:0] Wgt_0_632,
input [18:0] Wgt_0_633,
input [18:0] Wgt_0_634,
input [18:0] Wgt_0_635,
input [18:0] Wgt_0_636,
input [18:0] Wgt_0_637,
input [18:0] Wgt_0_638,
input [18:0] Wgt_0_639,
input [18:0] Wgt_0_640,
input [18:0] Wgt_0_641,
input [18:0] Wgt_0_642,
input [18:0] Wgt_0_643,
input [18:0] Wgt_0_644,
input [18:0] Wgt_0_645,
input [18:0] Wgt_0_646,
input [18:0] Wgt_0_647,
input [18:0] Wgt_0_648,
input [18:0] Wgt_0_649,
input [18:0] Wgt_0_650,
input [18:0] Wgt_0_651,
input [18:0] Wgt_0_652,
input [18:0] Wgt_0_653,
input [18:0] Wgt_0_654,
input [18:0] Wgt_0_655,
input [18:0] Wgt_0_656,
input [18:0] Wgt_0_657,
input [18:0] Wgt_0_658,
input [18:0] Wgt_0_659,
input [18:0] Wgt_0_660,
input [18:0] Wgt_0_661,
input [18:0] Wgt_0_662,
input [18:0] Wgt_0_663,
input [18:0] Wgt_0_664,
input [18:0] Wgt_0_665,
input [18:0] Wgt_0_666,
input [18:0] Wgt_0_667,
input [18:0] Wgt_0_668,
input [18:0] Wgt_0_669,
input [18:0] Wgt_0_670,
input [18:0] Wgt_0_671,
input [18:0] Wgt_0_672,
input [18:0] Wgt_0_673,
input [18:0] Wgt_0_674,
input [18:0] Wgt_0_675,
input [18:0] Wgt_0_676,
input [18:0] Wgt_0_677,
input [18:0] Wgt_0_678,
input [18:0] Wgt_0_679,
input [18:0] Wgt_0_680,
input [18:0] Wgt_0_681,
input [18:0] Wgt_0_682,
input [18:0] Wgt_0_683,
input [18:0] Wgt_0_684,
input [18:0] Wgt_0_685,
input [18:0] Wgt_0_686,
input [18:0] Wgt_0_687,
input [18:0] Wgt_0_688,
input [18:0] Wgt_0_689,
input [18:0] Wgt_0_690,
input [18:0] Wgt_0_691,
input [18:0] Wgt_0_692,
input [18:0] Wgt_0_693,
input [18:0] Wgt_0_694,
input [18:0] Wgt_0_695,
input [18:0] Wgt_0_696,
input [18:0] Wgt_0_697,
input [18:0] Wgt_0_698,
input [18:0] Wgt_0_699,
input [18:0] Wgt_0_700,
input [18:0] Wgt_0_701,
input [18:0] Wgt_0_702,
input [18:0] Wgt_0_703,
input [18:0] Wgt_0_704,
input [18:0] Wgt_0_705,
input [18:0] Wgt_0_706,
input [18:0] Wgt_0_707,
input [18:0] Wgt_0_708,
input [18:0] Wgt_0_709,
input [18:0] Wgt_0_710,
input [18:0] Wgt_0_711,
input [18:0] Wgt_0_712,
input [18:0] Wgt_0_713,
input [18:0] Wgt_0_714,
input [18:0] Wgt_0_715,
input [18:0] Wgt_0_716,
input [18:0] Wgt_0_717,
input [18:0] Wgt_0_718,
input [18:0] Wgt_0_719,
input [18:0] Wgt_0_720,
input [18:0] Wgt_0_721,
input [18:0] Wgt_0_722,
input [18:0] Wgt_0_723,
input [18:0] Wgt_0_724,
input [18:0] Wgt_0_725,
input [18:0] Wgt_0_726,
input [18:0] Wgt_0_727,
input [18:0] Wgt_0_728,
input [18:0] Wgt_0_729,
input [18:0] Wgt_0_730,
input [18:0] Wgt_0_731,
input [18:0] Wgt_0_732,
input [18:0] Wgt_0_733,
input [18:0] Wgt_0_734,
input [18:0] Wgt_0_735,
input [18:0] Wgt_0_736,
input [18:0] Wgt_0_737,
input [18:0] Wgt_0_738,
input [18:0] Wgt_0_739,
input [18:0] Wgt_0_740,
input [18:0] Wgt_0_741,
input [18:0] Wgt_0_742,
input [18:0] Wgt_0_743,
input [18:0] Wgt_0_744,
input [18:0] Wgt_0_745,
input [18:0] Wgt_0_746,
input [18:0] Wgt_0_747,
input [18:0] Wgt_0_748,
input [18:0] Wgt_0_749,
input [18:0] Wgt_0_750,
input [18:0] Wgt_0_751,
input [18:0] Wgt_0_752,
input [18:0] Wgt_0_753,
input [18:0] Wgt_0_754,
input [18:0] Wgt_0_755,
input [18:0] Wgt_0_756,
input [18:0] Wgt_0_757,
input [18:0] Wgt_0_758,
input [18:0] Wgt_0_759,
input [18:0] Wgt_0_760,
input [18:0] Wgt_0_761,
input [18:0] Wgt_0_762,
input [18:0] Wgt_0_763,
input [18:0] Wgt_0_764,
input [18:0] Wgt_0_765,
input [18:0] Wgt_0_766,
input [18:0] Wgt_0_767,
input [18:0] Wgt_0_768,
input [18:0] Wgt_0_769,
input [18:0] Wgt_0_770,
input [18:0] Wgt_0_771,
input [18:0] Wgt_0_772,
input [18:0] Wgt_0_773,
input [18:0] Wgt_0_774,
input [18:0] Wgt_0_775,
input [18:0] Wgt_0_776,
input [18:0] Wgt_0_777,
input [18:0] Wgt_0_778,
input [18:0] Wgt_0_779,
input [18:0] Wgt_0_780,
input [18:0] Wgt_0_781,
input [18:0] Wgt_0_782,
input [18:0] Wgt_0_783,
input [18:0] Wgt_0_784,
input [18:0] Wgt_1_0,
input [18:0] Wgt_1_1,
input [18:0] Wgt_1_2,
input [18:0] Wgt_1_3,
input [18:0] Wgt_1_4,
input [18:0] Wgt_1_5,
input [18:0] Wgt_1_6,
input [18:0] Wgt_1_7,
input [18:0] Wgt_1_8,
input [18:0] Wgt_1_9,
input [18:0] Wgt_1_10,
input [18:0] Wgt_1_11,
input [18:0] Wgt_1_12,
input [18:0] Wgt_1_13,
input [18:0] Wgt_1_14,
input [18:0] Wgt_1_15,
input [18:0] Wgt_1_16,
input [18:0] Wgt_1_17,
input [18:0] Wgt_1_18,
input [18:0] Wgt_1_19,
input [18:0] Wgt_1_20,
input [18:0] Wgt_1_21,
input [18:0] Wgt_1_22,
input [18:0] Wgt_1_23,
input [18:0] Wgt_1_24,
input [18:0] Wgt_1_25,
input [18:0] Wgt_1_26,
input [18:0] Wgt_1_27,
input [18:0] Wgt_1_28,
input [18:0] Wgt_1_29,
input [18:0] Wgt_1_30,
input [18:0] Wgt_1_31,
input [18:0] Wgt_1_32,
input [18:0] Wgt_1_33,
input [18:0] Wgt_1_34,
input [18:0] Wgt_1_35,
input [18:0] Wgt_1_36,
input [18:0] Wgt_1_37,
input [18:0] Wgt_1_38,
input [18:0] Wgt_1_39,
input [18:0] Wgt_1_40,
input [18:0] Wgt_1_41,
input [18:0] Wgt_1_42,
input [18:0] Wgt_1_43,
input [18:0] Wgt_1_44,
input [18:0] Wgt_1_45,
input [18:0] Wgt_1_46,
input [18:0] Wgt_1_47,
input [18:0] Wgt_1_48,
input [18:0] Wgt_1_49,
input [18:0] Wgt_1_50,
input [18:0] Wgt_1_51,
input [18:0] Wgt_1_52,
input [18:0] Wgt_1_53,
input [18:0] Wgt_1_54,
input [18:0] Wgt_1_55,
input [18:0] Wgt_1_56,
input [18:0] Wgt_1_57,
input [18:0] Wgt_1_58,
input [18:0] Wgt_1_59,
input [18:0] Wgt_1_60,
input [18:0] Wgt_1_61,
input [18:0] Wgt_1_62,
input [18:0] Wgt_1_63,
input [18:0] Wgt_1_64,
input [18:0] Wgt_1_65,
input [18:0] Wgt_1_66,
input [18:0] Wgt_1_67,
input [18:0] Wgt_1_68,
input [18:0] Wgt_1_69,
input [18:0] Wgt_1_70,
input [18:0] Wgt_1_71,
input [18:0] Wgt_1_72,
input [18:0] Wgt_1_73,
input [18:0] Wgt_1_74,
input [18:0] Wgt_1_75,
input [18:0] Wgt_1_76,
input [18:0] Wgt_1_77,
input [18:0] Wgt_1_78,
input [18:0] Wgt_1_79,
input [18:0] Wgt_1_80,
input [18:0] Wgt_1_81,
input [18:0] Wgt_1_82,
input [18:0] Wgt_1_83,
input [18:0] Wgt_1_84,
input [18:0] Wgt_1_85,
input [18:0] Wgt_1_86,
input [18:0] Wgt_1_87,
input [18:0] Wgt_1_88,
input [18:0] Wgt_1_89,
input [18:0] Wgt_1_90,
input [18:0] Wgt_1_91,
input [18:0] Wgt_1_92,
input [18:0] Wgt_1_93,
input [18:0] Wgt_1_94,
input [18:0] Wgt_1_95,
input [18:0] Wgt_1_96,
input [18:0] Wgt_1_97,
input [18:0] Wgt_1_98,
input [18:0] Wgt_1_99,
input [18:0] Wgt_1_100,
input [18:0] Wgt_1_101,
input [18:0] Wgt_1_102,
input [18:0] Wgt_1_103,
input [18:0] Wgt_1_104,
input [18:0] Wgt_1_105,
input [18:0] Wgt_1_106,
input [18:0] Wgt_1_107,
input [18:0] Wgt_1_108,
input [18:0] Wgt_1_109,
input [18:0] Wgt_1_110,
input [18:0] Wgt_1_111,
input [18:0] Wgt_1_112,
input [18:0] Wgt_1_113,
input [18:0] Wgt_1_114,
input [18:0] Wgt_1_115,
input [18:0] Wgt_1_116,
input [18:0] Wgt_1_117,
input [18:0] Wgt_1_118,
input [18:0] Wgt_1_119,
input [18:0] Wgt_1_120,
input [18:0] Wgt_1_121,
input [18:0] Wgt_1_122,
input [18:0] Wgt_1_123,
input [18:0] Wgt_1_124,
input [18:0] Wgt_1_125,
input [18:0] Wgt_1_126,
input [18:0] Wgt_1_127,
input [18:0] Wgt_1_128,
input [18:0] Wgt_1_129,
input [18:0] Wgt_1_130,
input [18:0] Wgt_1_131,
input [18:0] Wgt_1_132,
input [18:0] Wgt_1_133,
input [18:0] Wgt_1_134,
input [18:0] Wgt_1_135,
input [18:0] Wgt_1_136,
input [18:0] Wgt_1_137,
input [18:0] Wgt_1_138,
input [18:0] Wgt_1_139,
input [18:0] Wgt_1_140,
input [18:0] Wgt_1_141,
input [18:0] Wgt_1_142,
input [18:0] Wgt_1_143,
input [18:0] Wgt_1_144,
input [18:0] Wgt_1_145,
input [18:0] Wgt_1_146,
input [18:0] Wgt_1_147,
input [18:0] Wgt_1_148,
input [18:0] Wgt_1_149,
input [18:0] Wgt_1_150,
input [18:0] Wgt_1_151,
input [18:0] Wgt_1_152,
input [18:0] Wgt_1_153,
input [18:0] Wgt_1_154,
input [18:0] Wgt_1_155,
input [18:0] Wgt_1_156,
input [18:0] Wgt_1_157,
input [18:0] Wgt_1_158,
input [18:0] Wgt_1_159,
input [18:0] Wgt_1_160,
input [18:0] Wgt_1_161,
input [18:0] Wgt_1_162,
input [18:0] Wgt_1_163,
input [18:0] Wgt_1_164,
input [18:0] Wgt_1_165,
input [18:0] Wgt_1_166,
input [18:0] Wgt_1_167,
input [18:0] Wgt_1_168,
input [18:0] Wgt_1_169,
input [18:0] Wgt_1_170,
input [18:0] Wgt_1_171,
input [18:0] Wgt_1_172,
input [18:0] Wgt_1_173,
input [18:0] Wgt_1_174,
input [18:0] Wgt_1_175,
input [18:0] Wgt_1_176,
input [18:0] Wgt_1_177,
input [18:0] Wgt_1_178,
input [18:0] Wgt_1_179,
input [18:0] Wgt_1_180,
input [18:0] Wgt_1_181,
input [18:0] Wgt_1_182,
input [18:0] Wgt_1_183,
input [18:0] Wgt_1_184,
input [18:0] Wgt_1_185,
input [18:0] Wgt_1_186,
input [18:0] Wgt_1_187,
input [18:0] Wgt_1_188,
input [18:0] Wgt_1_189,
input [18:0] Wgt_1_190,
input [18:0] Wgt_1_191,
input [18:0] Wgt_1_192,
input [18:0] Wgt_1_193,
input [18:0] Wgt_1_194,
input [18:0] Wgt_1_195,
input [18:0] Wgt_1_196,
input [18:0] Wgt_1_197,
input [18:0] Wgt_1_198,
input [18:0] Wgt_1_199,
input [18:0] Wgt_1_200,
input [18:0] Wgt_1_201,
input [18:0] Wgt_1_202,
input [18:0] Wgt_1_203,
input [18:0] Wgt_1_204,
input [18:0] Wgt_1_205,
input [18:0] Wgt_1_206,
input [18:0] Wgt_1_207,
input [18:0] Wgt_1_208,
input [18:0] Wgt_1_209,
input [18:0] Wgt_1_210,
input [18:0] Wgt_1_211,
input [18:0] Wgt_1_212,
input [18:0] Wgt_1_213,
input [18:0] Wgt_1_214,
input [18:0] Wgt_1_215,
input [18:0] Wgt_1_216,
input [18:0] Wgt_1_217,
input [18:0] Wgt_1_218,
input [18:0] Wgt_1_219,
input [18:0] Wgt_1_220,
input [18:0] Wgt_1_221,
input [18:0] Wgt_1_222,
input [18:0] Wgt_1_223,
input [18:0] Wgt_1_224,
input [18:0] Wgt_1_225,
input [18:0] Wgt_1_226,
input [18:0] Wgt_1_227,
input [18:0] Wgt_1_228,
input [18:0] Wgt_1_229,
input [18:0] Wgt_1_230,
input [18:0] Wgt_1_231,
input [18:0] Wgt_1_232,
input [18:0] Wgt_1_233,
input [18:0] Wgt_1_234,
input [18:0] Wgt_1_235,
input [18:0] Wgt_1_236,
input [18:0] Wgt_1_237,
input [18:0] Wgt_1_238,
input [18:0] Wgt_1_239,
input [18:0] Wgt_1_240,
input [18:0] Wgt_1_241,
input [18:0] Wgt_1_242,
input [18:0] Wgt_1_243,
input [18:0] Wgt_1_244,
input [18:0] Wgt_1_245,
input [18:0] Wgt_1_246,
input [18:0] Wgt_1_247,
input [18:0] Wgt_1_248,
input [18:0] Wgt_1_249,
input [18:0] Wgt_1_250,
input [18:0] Wgt_1_251,
input [18:0] Wgt_1_252,
input [18:0] Wgt_1_253,
input [18:0] Wgt_1_254,
input [18:0] Wgt_1_255,
input [18:0] Wgt_1_256,
input [18:0] Wgt_1_257,
input [18:0] Wgt_1_258,
input [18:0] Wgt_1_259,
input [18:0] Wgt_1_260,
input [18:0] Wgt_1_261,
input [18:0] Wgt_1_262,
input [18:0] Wgt_1_263,
input [18:0] Wgt_1_264,
input [18:0] Wgt_1_265,
input [18:0] Wgt_1_266,
input [18:0] Wgt_1_267,
input [18:0] Wgt_1_268,
input [18:0] Wgt_1_269,
input [18:0] Wgt_1_270,
input [18:0] Wgt_1_271,
input [18:0] Wgt_1_272,
input [18:0] Wgt_1_273,
input [18:0] Wgt_1_274,
input [18:0] Wgt_1_275,
input [18:0] Wgt_1_276,
input [18:0] Wgt_1_277,
input [18:0] Wgt_1_278,
input [18:0] Wgt_1_279,
input [18:0] Wgt_1_280,
input [18:0] Wgt_1_281,
input [18:0] Wgt_1_282,
input [18:0] Wgt_1_283,
input [18:0] Wgt_1_284,
input [18:0] Wgt_1_285,
input [18:0] Wgt_1_286,
input [18:0] Wgt_1_287,
input [18:0] Wgt_1_288,
input [18:0] Wgt_1_289,
input [18:0] Wgt_1_290,
input [18:0] Wgt_1_291,
input [18:0] Wgt_1_292,
input [18:0] Wgt_1_293,
input [18:0] Wgt_1_294,
input [18:0] Wgt_1_295,
input [18:0] Wgt_1_296,
input [18:0] Wgt_1_297,
input [18:0] Wgt_1_298,
input [18:0] Wgt_1_299,
input [18:0] Wgt_1_300,
input [18:0] Wgt_1_301,
input [18:0] Wgt_1_302,
input [18:0] Wgt_1_303,
input [18:0] Wgt_1_304,
input [18:0] Wgt_1_305,
input [18:0] Wgt_1_306,
input [18:0] Wgt_1_307,
input [18:0] Wgt_1_308,
input [18:0] Wgt_1_309,
input [18:0] Wgt_1_310,
input [18:0] Wgt_1_311,
input [18:0] Wgt_1_312,
input [18:0] Wgt_1_313,
input [18:0] Wgt_1_314,
input [18:0] Wgt_1_315,
input [18:0] Wgt_1_316,
input [18:0] Wgt_1_317,
input [18:0] Wgt_1_318,
input [18:0] Wgt_1_319,
input [18:0] Wgt_1_320,
input [18:0] Wgt_1_321,
input [18:0] Wgt_1_322,
input [18:0] Wgt_1_323,
input [18:0] Wgt_1_324,
input [18:0] Wgt_1_325,
input [18:0] Wgt_1_326,
input [18:0] Wgt_1_327,
input [18:0] Wgt_1_328,
input [18:0] Wgt_1_329,
input [18:0] Wgt_1_330,
input [18:0] Wgt_1_331,
input [18:0] Wgt_1_332,
input [18:0] Wgt_1_333,
input [18:0] Wgt_1_334,
input [18:0] Wgt_1_335,
input [18:0] Wgt_1_336,
input [18:0] Wgt_1_337,
input [18:0] Wgt_1_338,
input [18:0] Wgt_1_339,
input [18:0] Wgt_1_340,
input [18:0] Wgt_1_341,
input [18:0] Wgt_1_342,
input [18:0] Wgt_1_343,
input [18:0] Wgt_1_344,
input [18:0] Wgt_1_345,
input [18:0] Wgt_1_346,
input [18:0] Wgt_1_347,
input [18:0] Wgt_1_348,
input [18:0] Wgt_1_349,
input [18:0] Wgt_1_350,
input [18:0] Wgt_1_351,
input [18:0] Wgt_1_352,
input [18:0] Wgt_1_353,
input [18:0] Wgt_1_354,
input [18:0] Wgt_1_355,
input [18:0] Wgt_1_356,
input [18:0] Wgt_1_357,
input [18:0] Wgt_1_358,
input [18:0] Wgt_1_359,
input [18:0] Wgt_1_360,
input [18:0] Wgt_1_361,
input [18:0] Wgt_1_362,
input [18:0] Wgt_1_363,
input [18:0] Wgt_1_364,
input [18:0] Wgt_1_365,
input [18:0] Wgt_1_366,
input [18:0] Wgt_1_367,
input [18:0] Wgt_1_368,
input [18:0] Wgt_1_369,
input [18:0] Wgt_1_370,
input [18:0] Wgt_1_371,
input [18:0] Wgt_1_372,
input [18:0] Wgt_1_373,
input [18:0] Wgt_1_374,
input [18:0] Wgt_1_375,
input [18:0] Wgt_1_376,
input [18:0] Wgt_1_377,
input [18:0] Wgt_1_378,
input [18:0] Wgt_1_379,
input [18:0] Wgt_1_380,
input [18:0] Wgt_1_381,
input [18:0] Wgt_1_382,
input [18:0] Wgt_1_383,
input [18:0] Wgt_1_384,
input [18:0] Wgt_1_385,
input [18:0] Wgt_1_386,
input [18:0] Wgt_1_387,
input [18:0] Wgt_1_388,
input [18:0] Wgt_1_389,
input [18:0] Wgt_1_390,
input [18:0] Wgt_1_391,
input [18:0] Wgt_1_392,
input [18:0] Wgt_1_393,
input [18:0] Wgt_1_394,
input [18:0] Wgt_1_395,
input [18:0] Wgt_1_396,
input [18:0] Wgt_1_397,
input [18:0] Wgt_1_398,
input [18:0] Wgt_1_399,
input [18:0] Wgt_1_400,
input [18:0] Wgt_1_401,
input [18:0] Wgt_1_402,
input [18:0] Wgt_1_403,
input [18:0] Wgt_1_404,
input [18:0] Wgt_1_405,
input [18:0] Wgt_1_406,
input [18:0] Wgt_1_407,
input [18:0] Wgt_1_408,
input [18:0] Wgt_1_409,
input [18:0] Wgt_1_410,
input [18:0] Wgt_1_411,
input [18:0] Wgt_1_412,
input [18:0] Wgt_1_413,
input [18:0] Wgt_1_414,
input [18:0] Wgt_1_415,
input [18:0] Wgt_1_416,
input [18:0] Wgt_1_417,
input [18:0] Wgt_1_418,
input [18:0] Wgt_1_419,
input [18:0] Wgt_1_420,
input [18:0] Wgt_1_421,
input [18:0] Wgt_1_422,
input [18:0] Wgt_1_423,
input [18:0] Wgt_1_424,
input [18:0] Wgt_1_425,
input [18:0] Wgt_1_426,
input [18:0] Wgt_1_427,
input [18:0] Wgt_1_428,
input [18:0] Wgt_1_429,
input [18:0] Wgt_1_430,
input [18:0] Wgt_1_431,
input [18:0] Wgt_1_432,
input [18:0] Wgt_1_433,
input [18:0] Wgt_1_434,
input [18:0] Wgt_1_435,
input [18:0] Wgt_1_436,
input [18:0] Wgt_1_437,
input [18:0] Wgt_1_438,
input [18:0] Wgt_1_439,
input [18:0] Wgt_1_440,
input [18:0] Wgt_1_441,
input [18:0] Wgt_1_442,
input [18:0] Wgt_1_443,
input [18:0] Wgt_1_444,
input [18:0] Wgt_1_445,
input [18:0] Wgt_1_446,
input [18:0] Wgt_1_447,
input [18:0] Wgt_1_448,
input [18:0] Wgt_1_449,
input [18:0] Wgt_1_450,
input [18:0] Wgt_1_451,
input [18:0] Wgt_1_452,
input [18:0] Wgt_1_453,
input [18:0] Wgt_1_454,
input [18:0] Wgt_1_455,
input [18:0] Wgt_1_456,
input [18:0] Wgt_1_457,
input [18:0] Wgt_1_458,
input [18:0] Wgt_1_459,
input [18:0] Wgt_1_460,
input [18:0] Wgt_1_461,
input [18:0] Wgt_1_462,
input [18:0] Wgt_1_463,
input [18:0] Wgt_1_464,
input [18:0] Wgt_1_465,
input [18:0] Wgt_1_466,
input [18:0] Wgt_1_467,
input [18:0] Wgt_1_468,
input [18:0] Wgt_1_469,
input [18:0] Wgt_1_470,
input [18:0] Wgt_1_471,
input [18:0] Wgt_1_472,
input [18:0] Wgt_1_473,
input [18:0] Wgt_1_474,
input [18:0] Wgt_1_475,
input [18:0] Wgt_1_476,
input [18:0] Wgt_1_477,
input [18:0] Wgt_1_478,
input [18:0] Wgt_1_479,
input [18:0] Wgt_1_480,
input [18:0] Wgt_1_481,
input [18:0] Wgt_1_482,
input [18:0] Wgt_1_483,
input [18:0] Wgt_1_484,
input [18:0] Wgt_1_485,
input [18:0] Wgt_1_486,
input [18:0] Wgt_1_487,
input [18:0] Wgt_1_488,
input [18:0] Wgt_1_489,
input [18:0] Wgt_1_490,
input [18:0] Wgt_1_491,
input [18:0] Wgt_1_492,
input [18:0] Wgt_1_493,
input [18:0] Wgt_1_494,
input [18:0] Wgt_1_495,
input [18:0] Wgt_1_496,
input [18:0] Wgt_1_497,
input [18:0] Wgt_1_498,
input [18:0] Wgt_1_499,
input [18:0] Wgt_1_500,
input [18:0] Wgt_1_501,
input [18:0] Wgt_1_502,
input [18:0] Wgt_1_503,
input [18:0] Wgt_1_504,
input [18:0] Wgt_1_505,
input [18:0] Wgt_1_506,
input [18:0] Wgt_1_507,
input [18:0] Wgt_1_508,
input [18:0] Wgt_1_509,
input [18:0] Wgt_1_510,
input [18:0] Wgt_1_511,
input [18:0] Wgt_1_512,
input [18:0] Wgt_1_513,
input [18:0] Wgt_1_514,
input [18:0] Wgt_1_515,
input [18:0] Wgt_1_516,
input [18:0] Wgt_1_517,
input [18:0] Wgt_1_518,
input [18:0] Wgt_1_519,
input [18:0] Wgt_1_520,
input [18:0] Wgt_1_521,
input [18:0] Wgt_1_522,
input [18:0] Wgt_1_523,
input [18:0] Wgt_1_524,
input [18:0] Wgt_1_525,
input [18:0] Wgt_1_526,
input [18:0] Wgt_1_527,
input [18:0] Wgt_1_528,
input [18:0] Wgt_1_529,
input [18:0] Wgt_1_530,
input [18:0] Wgt_1_531,
input [18:0] Wgt_1_532,
input [18:0] Wgt_1_533,
input [18:0] Wgt_1_534,
input [18:0] Wgt_1_535,
input [18:0] Wgt_1_536,
input [18:0] Wgt_1_537,
input [18:0] Wgt_1_538,
input [18:0] Wgt_1_539,
input [18:0] Wgt_1_540,
input [18:0] Wgt_1_541,
input [18:0] Wgt_1_542,
input [18:0] Wgt_1_543,
input [18:0] Wgt_1_544,
input [18:0] Wgt_1_545,
input [18:0] Wgt_1_546,
input [18:0] Wgt_1_547,
input [18:0] Wgt_1_548,
input [18:0] Wgt_1_549,
input [18:0] Wgt_1_550,
input [18:0] Wgt_1_551,
input [18:0] Wgt_1_552,
input [18:0] Wgt_1_553,
input [18:0] Wgt_1_554,
input [18:0] Wgt_1_555,
input [18:0] Wgt_1_556,
input [18:0] Wgt_1_557,
input [18:0] Wgt_1_558,
input [18:0] Wgt_1_559,
input [18:0] Wgt_1_560,
input [18:0] Wgt_1_561,
input [18:0] Wgt_1_562,
input [18:0] Wgt_1_563,
input [18:0] Wgt_1_564,
input [18:0] Wgt_1_565,
input [18:0] Wgt_1_566,
input [18:0] Wgt_1_567,
input [18:0] Wgt_1_568,
input [18:0] Wgt_1_569,
input [18:0] Wgt_1_570,
input [18:0] Wgt_1_571,
input [18:0] Wgt_1_572,
input [18:0] Wgt_1_573,
input [18:0] Wgt_1_574,
input [18:0] Wgt_1_575,
input [18:0] Wgt_1_576,
input [18:0] Wgt_1_577,
input [18:0] Wgt_1_578,
input [18:0] Wgt_1_579,
input [18:0] Wgt_1_580,
input [18:0] Wgt_1_581,
input [18:0] Wgt_1_582,
input [18:0] Wgt_1_583,
input [18:0] Wgt_1_584,
input [18:0] Wgt_1_585,
input [18:0] Wgt_1_586,
input [18:0] Wgt_1_587,
input [18:0] Wgt_1_588,
input [18:0] Wgt_1_589,
input [18:0] Wgt_1_590,
input [18:0] Wgt_1_591,
input [18:0] Wgt_1_592,
input [18:0] Wgt_1_593,
input [18:0] Wgt_1_594,
input [18:0] Wgt_1_595,
input [18:0] Wgt_1_596,
input [18:0] Wgt_1_597,
input [18:0] Wgt_1_598,
input [18:0] Wgt_1_599,
input [18:0] Wgt_1_600,
input [18:0] Wgt_1_601,
input [18:0] Wgt_1_602,
input [18:0] Wgt_1_603,
input [18:0] Wgt_1_604,
input [18:0] Wgt_1_605,
input [18:0] Wgt_1_606,
input [18:0] Wgt_1_607,
input [18:0] Wgt_1_608,
input [18:0] Wgt_1_609,
input [18:0] Wgt_1_610,
input [18:0] Wgt_1_611,
input [18:0] Wgt_1_612,
input [18:0] Wgt_1_613,
input [18:0] Wgt_1_614,
input [18:0] Wgt_1_615,
input [18:0] Wgt_1_616,
input [18:0] Wgt_1_617,
input [18:0] Wgt_1_618,
input [18:0] Wgt_1_619,
input [18:0] Wgt_1_620,
input [18:0] Wgt_1_621,
input [18:0] Wgt_1_622,
input [18:0] Wgt_1_623,
input [18:0] Wgt_1_624,
input [18:0] Wgt_1_625,
input [18:0] Wgt_1_626,
input [18:0] Wgt_1_627,
input [18:0] Wgt_1_628,
input [18:0] Wgt_1_629,
input [18:0] Wgt_1_630,
input [18:0] Wgt_1_631,
input [18:0] Wgt_1_632,
input [18:0] Wgt_1_633,
input [18:0] Wgt_1_634,
input [18:0] Wgt_1_635,
input [18:0] Wgt_1_636,
input [18:0] Wgt_1_637,
input [18:0] Wgt_1_638,
input [18:0] Wgt_1_639,
input [18:0] Wgt_1_640,
input [18:0] Wgt_1_641,
input [18:0] Wgt_1_642,
input [18:0] Wgt_1_643,
input [18:0] Wgt_1_644,
input [18:0] Wgt_1_645,
input [18:0] Wgt_1_646,
input [18:0] Wgt_1_647,
input [18:0] Wgt_1_648,
input [18:0] Wgt_1_649,
input [18:0] Wgt_1_650,
input [18:0] Wgt_1_651,
input [18:0] Wgt_1_652,
input [18:0] Wgt_1_653,
input [18:0] Wgt_1_654,
input [18:0] Wgt_1_655,
input [18:0] Wgt_1_656,
input [18:0] Wgt_1_657,
input [18:0] Wgt_1_658,
input [18:0] Wgt_1_659,
input [18:0] Wgt_1_660,
input [18:0] Wgt_1_661,
input [18:0] Wgt_1_662,
input [18:0] Wgt_1_663,
input [18:0] Wgt_1_664,
input [18:0] Wgt_1_665,
input [18:0] Wgt_1_666,
input [18:0] Wgt_1_667,
input [18:0] Wgt_1_668,
input [18:0] Wgt_1_669,
input [18:0] Wgt_1_670,
input [18:0] Wgt_1_671,
input [18:0] Wgt_1_672,
input [18:0] Wgt_1_673,
input [18:0] Wgt_1_674,
input [18:0] Wgt_1_675,
input [18:0] Wgt_1_676,
input [18:0] Wgt_1_677,
input [18:0] Wgt_1_678,
input [18:0] Wgt_1_679,
input [18:0] Wgt_1_680,
input [18:0] Wgt_1_681,
input [18:0] Wgt_1_682,
input [18:0] Wgt_1_683,
input [18:0] Wgt_1_684,
input [18:0] Wgt_1_685,
input [18:0] Wgt_1_686,
input [18:0] Wgt_1_687,
input [18:0] Wgt_1_688,
input [18:0] Wgt_1_689,
input [18:0] Wgt_1_690,
input [18:0] Wgt_1_691,
input [18:0] Wgt_1_692,
input [18:0] Wgt_1_693,
input [18:0] Wgt_1_694,
input [18:0] Wgt_1_695,
input [18:0] Wgt_1_696,
input [18:0] Wgt_1_697,
input [18:0] Wgt_1_698,
input [18:0] Wgt_1_699,
input [18:0] Wgt_1_700,
input [18:0] Wgt_1_701,
input [18:0] Wgt_1_702,
input [18:0] Wgt_1_703,
input [18:0] Wgt_1_704,
input [18:0] Wgt_1_705,
input [18:0] Wgt_1_706,
input [18:0] Wgt_1_707,
input [18:0] Wgt_1_708,
input [18:0] Wgt_1_709,
input [18:0] Wgt_1_710,
input [18:0] Wgt_1_711,
input [18:0] Wgt_1_712,
input [18:0] Wgt_1_713,
input [18:0] Wgt_1_714,
input [18:0] Wgt_1_715,
input [18:0] Wgt_1_716,
input [18:0] Wgt_1_717,
input [18:0] Wgt_1_718,
input [18:0] Wgt_1_719,
input [18:0] Wgt_1_720,
input [18:0] Wgt_1_721,
input [18:0] Wgt_1_722,
input [18:0] Wgt_1_723,
input [18:0] Wgt_1_724,
input [18:0] Wgt_1_725,
input [18:0] Wgt_1_726,
input [18:0] Wgt_1_727,
input [18:0] Wgt_1_728,
input [18:0] Wgt_1_729,
input [18:0] Wgt_1_730,
input [18:0] Wgt_1_731,
input [18:0] Wgt_1_732,
input [18:0] Wgt_1_733,
input [18:0] Wgt_1_734,
input [18:0] Wgt_1_735,
input [18:0] Wgt_1_736,
input [18:0] Wgt_1_737,
input [18:0] Wgt_1_738,
input [18:0] Wgt_1_739,
input [18:0] Wgt_1_740,
input [18:0] Wgt_1_741,
input [18:0] Wgt_1_742,
input [18:0] Wgt_1_743,
input [18:0] Wgt_1_744,
input [18:0] Wgt_1_745,
input [18:0] Wgt_1_746,
input [18:0] Wgt_1_747,
input [18:0] Wgt_1_748,
input [18:0] Wgt_1_749,
input [18:0] Wgt_1_750,
input [18:0] Wgt_1_751,
input [18:0] Wgt_1_752,
input [18:0] Wgt_1_753,
input [18:0] Wgt_1_754,
input [18:0] Wgt_1_755,
input [18:0] Wgt_1_756,
input [18:0] Wgt_1_757,
input [18:0] Wgt_1_758,
input [18:0] Wgt_1_759,
input [18:0] Wgt_1_760,
input [18:0] Wgt_1_761,
input [18:0] Wgt_1_762,
input [18:0] Wgt_1_763,
input [18:0] Wgt_1_764,
input [18:0] Wgt_1_765,
input [18:0] Wgt_1_766,
input [18:0] Wgt_1_767,
input [18:0] Wgt_1_768,
input [18:0] Wgt_1_769,
input [18:0] Wgt_1_770,
input [18:0] Wgt_1_771,
input [18:0] Wgt_1_772,
input [18:0] Wgt_1_773,
input [18:0] Wgt_1_774,
input [18:0] Wgt_1_775,
input [18:0] Wgt_1_776,
input [18:0] Wgt_1_777,
input [18:0] Wgt_1_778,
input [18:0] Wgt_1_779,
input [18:0] Wgt_1_780,
input [18:0] Wgt_1_781,
input [18:0] Wgt_1_782,
input [18:0] Wgt_1_783,
input [18:0] Wgt_1_784,
input [18:0] Wgt_2_0,
input [18:0] Wgt_2_1,
input [18:0] Wgt_2_2,
input [18:0] Wgt_2_3,
input [18:0] Wgt_2_4,
input [18:0] Wgt_2_5,
input [18:0] Wgt_2_6,
input [18:0] Wgt_2_7,
input [18:0] Wgt_2_8,
input [18:0] Wgt_2_9,
input [18:0] Wgt_2_10,
input [18:0] Wgt_2_11,
input [18:0] Wgt_2_12,
input [18:0] Wgt_2_13,
input [18:0] Wgt_2_14,
input [18:0] Wgt_2_15,
input [18:0] Wgt_2_16,
input [18:0] Wgt_2_17,
input [18:0] Wgt_2_18,
input [18:0] Wgt_2_19,
input [18:0] Wgt_2_20,
input [18:0] Wgt_2_21,
input [18:0] Wgt_2_22,
input [18:0] Wgt_2_23,
input [18:0] Wgt_2_24,
input [18:0] Wgt_2_25,
input [18:0] Wgt_2_26,
input [18:0] Wgt_2_27,
input [18:0] Wgt_2_28,
input [18:0] Wgt_2_29,
input [18:0] Wgt_2_30,
input [18:0] Wgt_2_31,
input [18:0] Wgt_2_32,
input [18:0] Wgt_2_33,
input [18:0] Wgt_2_34,
input [18:0] Wgt_2_35,
input [18:0] Wgt_2_36,
input [18:0] Wgt_2_37,
input [18:0] Wgt_2_38,
input [18:0] Wgt_2_39,
input [18:0] Wgt_2_40,
input [18:0] Wgt_2_41,
input [18:0] Wgt_2_42,
input [18:0] Wgt_2_43,
input [18:0] Wgt_2_44,
input [18:0] Wgt_2_45,
input [18:0] Wgt_2_46,
input [18:0] Wgt_2_47,
input [18:0] Wgt_2_48,
input [18:0] Wgt_2_49,
input [18:0] Wgt_2_50,
input [18:0] Wgt_2_51,
input [18:0] Wgt_2_52,
input [18:0] Wgt_2_53,
input [18:0] Wgt_2_54,
input [18:0] Wgt_2_55,
input [18:0] Wgt_2_56,
input [18:0] Wgt_2_57,
input [18:0] Wgt_2_58,
input [18:0] Wgt_2_59,
input [18:0] Wgt_2_60,
input [18:0] Wgt_2_61,
input [18:0] Wgt_2_62,
input [18:0] Wgt_2_63,
input [18:0] Wgt_2_64,
input [18:0] Wgt_2_65,
input [18:0] Wgt_2_66,
input [18:0] Wgt_2_67,
input [18:0] Wgt_2_68,
input [18:0] Wgt_2_69,
input [18:0] Wgt_2_70,
input [18:0] Wgt_2_71,
input [18:0] Wgt_2_72,
input [18:0] Wgt_2_73,
input [18:0] Wgt_2_74,
input [18:0] Wgt_2_75,
input [18:0] Wgt_2_76,
input [18:0] Wgt_2_77,
input [18:0] Wgt_2_78,
input [18:0] Wgt_2_79,
input [18:0] Wgt_2_80,
input [18:0] Wgt_2_81,
input [18:0] Wgt_2_82,
input [18:0] Wgt_2_83,
input [18:0] Wgt_2_84,
input [18:0] Wgt_2_85,
input [18:0] Wgt_2_86,
input [18:0] Wgt_2_87,
input [18:0] Wgt_2_88,
input [18:0] Wgt_2_89,
input [18:0] Wgt_2_90,
input [18:0] Wgt_2_91,
input [18:0] Wgt_2_92,
input [18:0] Wgt_2_93,
input [18:0] Wgt_2_94,
input [18:0] Wgt_2_95,
input [18:0] Wgt_2_96,
input [18:0] Wgt_2_97,
input [18:0] Wgt_2_98,
input [18:0] Wgt_2_99,
input [18:0] Wgt_2_100,
input [18:0] Wgt_2_101,
input [18:0] Wgt_2_102,
input [18:0] Wgt_2_103,
input [18:0] Wgt_2_104,
input [18:0] Wgt_2_105,
input [18:0] Wgt_2_106,
input [18:0] Wgt_2_107,
input [18:0] Wgt_2_108,
input [18:0] Wgt_2_109,
input [18:0] Wgt_2_110,
input [18:0] Wgt_2_111,
input [18:0] Wgt_2_112,
input [18:0] Wgt_2_113,
input [18:0] Wgt_2_114,
input [18:0] Wgt_2_115,
input [18:0] Wgt_2_116,
input [18:0] Wgt_2_117,
input [18:0] Wgt_2_118,
input [18:0] Wgt_2_119,
input [18:0] Wgt_2_120,
input [18:0] Wgt_2_121,
input [18:0] Wgt_2_122,
input [18:0] Wgt_2_123,
input [18:0] Wgt_2_124,
input [18:0] Wgt_2_125,
input [18:0] Wgt_2_126,
input [18:0] Wgt_2_127,
input [18:0] Wgt_2_128,
input [18:0] Wgt_2_129,
input [18:0] Wgt_2_130,
input [18:0] Wgt_2_131,
input [18:0] Wgt_2_132,
input [18:0] Wgt_2_133,
input [18:0] Wgt_2_134,
input [18:0] Wgt_2_135,
input [18:0] Wgt_2_136,
input [18:0] Wgt_2_137,
input [18:0] Wgt_2_138,
input [18:0] Wgt_2_139,
input [18:0] Wgt_2_140,
input [18:0] Wgt_2_141,
input [18:0] Wgt_2_142,
input [18:0] Wgt_2_143,
input [18:0] Wgt_2_144,
input [18:0] Wgt_2_145,
input [18:0] Wgt_2_146,
input [18:0] Wgt_2_147,
input [18:0] Wgt_2_148,
input [18:0] Wgt_2_149,
input [18:0] Wgt_2_150,
input [18:0] Wgt_2_151,
input [18:0] Wgt_2_152,
input [18:0] Wgt_2_153,
input [18:0] Wgt_2_154,
input [18:0] Wgt_2_155,
input [18:0] Wgt_2_156,
input [18:0] Wgt_2_157,
input [18:0] Wgt_2_158,
input [18:0] Wgt_2_159,
input [18:0] Wgt_2_160,
input [18:0] Wgt_2_161,
input [18:0] Wgt_2_162,
input [18:0] Wgt_2_163,
input [18:0] Wgt_2_164,
input [18:0] Wgt_2_165,
input [18:0] Wgt_2_166,
input [18:0] Wgt_2_167,
input [18:0] Wgt_2_168,
input [18:0] Wgt_2_169,
input [18:0] Wgt_2_170,
input [18:0] Wgt_2_171,
input [18:0] Wgt_2_172,
input [18:0] Wgt_2_173,
input [18:0] Wgt_2_174,
input [18:0] Wgt_2_175,
input [18:0] Wgt_2_176,
input [18:0] Wgt_2_177,
input [18:0] Wgt_2_178,
input [18:0] Wgt_2_179,
input [18:0] Wgt_2_180,
input [18:0] Wgt_2_181,
input [18:0] Wgt_2_182,
input [18:0] Wgt_2_183,
input [18:0] Wgt_2_184,
input [18:0] Wgt_2_185,
input [18:0] Wgt_2_186,
input [18:0] Wgt_2_187,
input [18:0] Wgt_2_188,
input [18:0] Wgt_2_189,
input [18:0] Wgt_2_190,
input [18:0] Wgt_2_191,
input [18:0] Wgt_2_192,
input [18:0] Wgt_2_193,
input [18:0] Wgt_2_194,
input [18:0] Wgt_2_195,
input [18:0] Wgt_2_196,
input [18:0] Wgt_2_197,
input [18:0] Wgt_2_198,
input [18:0] Wgt_2_199,
input [18:0] Wgt_2_200,
input [18:0] Wgt_2_201,
input [18:0] Wgt_2_202,
input [18:0] Wgt_2_203,
input [18:0] Wgt_2_204,
input [18:0] Wgt_2_205,
input [18:0] Wgt_2_206,
input [18:0] Wgt_2_207,
input [18:0] Wgt_2_208,
input [18:0] Wgt_2_209,
input [18:0] Wgt_2_210,
input [18:0] Wgt_2_211,
input [18:0] Wgt_2_212,
input [18:0] Wgt_2_213,
input [18:0] Wgt_2_214,
input [18:0] Wgt_2_215,
input [18:0] Wgt_2_216,
input [18:0] Wgt_2_217,
input [18:0] Wgt_2_218,
input [18:0] Wgt_2_219,
input [18:0] Wgt_2_220,
input [18:0] Wgt_2_221,
input [18:0] Wgt_2_222,
input [18:0] Wgt_2_223,
input [18:0] Wgt_2_224,
input [18:0] Wgt_2_225,
input [18:0] Wgt_2_226,
input [18:0] Wgt_2_227,
input [18:0] Wgt_2_228,
input [18:0] Wgt_2_229,
input [18:0] Wgt_2_230,
input [18:0] Wgt_2_231,
input [18:0] Wgt_2_232,
input [18:0] Wgt_2_233,
input [18:0] Wgt_2_234,
input [18:0] Wgt_2_235,
input [18:0] Wgt_2_236,
input [18:0] Wgt_2_237,
input [18:0] Wgt_2_238,
input [18:0] Wgt_2_239,
input [18:0] Wgt_2_240,
input [18:0] Wgt_2_241,
input [18:0] Wgt_2_242,
input [18:0] Wgt_2_243,
input [18:0] Wgt_2_244,
input [18:0] Wgt_2_245,
input [18:0] Wgt_2_246,
input [18:0] Wgt_2_247,
input [18:0] Wgt_2_248,
input [18:0] Wgt_2_249,
input [18:0] Wgt_2_250,
input [18:0] Wgt_2_251,
input [18:0] Wgt_2_252,
input [18:0] Wgt_2_253,
input [18:0] Wgt_2_254,
input [18:0] Wgt_2_255,
input [18:0] Wgt_2_256,
input [18:0] Wgt_2_257,
input [18:0] Wgt_2_258,
input [18:0] Wgt_2_259,
input [18:0] Wgt_2_260,
input [18:0] Wgt_2_261,
input [18:0] Wgt_2_262,
input [18:0] Wgt_2_263,
input [18:0] Wgt_2_264,
input [18:0] Wgt_2_265,
input [18:0] Wgt_2_266,
input [18:0] Wgt_2_267,
input [18:0] Wgt_2_268,
input [18:0] Wgt_2_269,
input [18:0] Wgt_2_270,
input [18:0] Wgt_2_271,
input [18:0] Wgt_2_272,
input [18:0] Wgt_2_273,
input [18:0] Wgt_2_274,
input [18:0] Wgt_2_275,
input [18:0] Wgt_2_276,
input [18:0] Wgt_2_277,
input [18:0] Wgt_2_278,
input [18:0] Wgt_2_279,
input [18:0] Wgt_2_280,
input [18:0] Wgt_2_281,
input [18:0] Wgt_2_282,
input [18:0] Wgt_2_283,
input [18:0] Wgt_2_284,
input [18:0] Wgt_2_285,
input [18:0] Wgt_2_286,
input [18:0] Wgt_2_287,
input [18:0] Wgt_2_288,
input [18:0] Wgt_2_289,
input [18:0] Wgt_2_290,
input [18:0] Wgt_2_291,
input [18:0] Wgt_2_292,
input [18:0] Wgt_2_293,
input [18:0] Wgt_2_294,
input [18:0] Wgt_2_295,
input [18:0] Wgt_2_296,
input [18:0] Wgt_2_297,
input [18:0] Wgt_2_298,
input [18:0] Wgt_2_299,
input [18:0] Wgt_2_300,
input [18:0] Wgt_2_301,
input [18:0] Wgt_2_302,
input [18:0] Wgt_2_303,
input [18:0] Wgt_2_304,
input [18:0] Wgt_2_305,
input [18:0] Wgt_2_306,
input [18:0] Wgt_2_307,
input [18:0] Wgt_2_308,
input [18:0] Wgt_2_309,
input [18:0] Wgt_2_310,
input [18:0] Wgt_2_311,
input [18:0] Wgt_2_312,
input [18:0] Wgt_2_313,
input [18:0] Wgt_2_314,
input [18:0] Wgt_2_315,
input [18:0] Wgt_2_316,
input [18:0] Wgt_2_317,
input [18:0] Wgt_2_318,
input [18:0] Wgt_2_319,
input [18:0] Wgt_2_320,
input [18:0] Wgt_2_321,
input [18:0] Wgt_2_322,
input [18:0] Wgt_2_323,
input [18:0] Wgt_2_324,
input [18:0] Wgt_2_325,
input [18:0] Wgt_2_326,
input [18:0] Wgt_2_327,
input [18:0] Wgt_2_328,
input [18:0] Wgt_2_329,
input [18:0] Wgt_2_330,
input [18:0] Wgt_2_331,
input [18:0] Wgt_2_332,
input [18:0] Wgt_2_333,
input [18:0] Wgt_2_334,
input [18:0] Wgt_2_335,
input [18:0] Wgt_2_336,
input [18:0] Wgt_2_337,
input [18:0] Wgt_2_338,
input [18:0] Wgt_2_339,
input [18:0] Wgt_2_340,
input [18:0] Wgt_2_341,
input [18:0] Wgt_2_342,
input [18:0] Wgt_2_343,
input [18:0] Wgt_2_344,
input [18:0] Wgt_2_345,
input [18:0] Wgt_2_346,
input [18:0] Wgt_2_347,
input [18:0] Wgt_2_348,
input [18:0] Wgt_2_349,
input [18:0] Wgt_2_350,
input [18:0] Wgt_2_351,
input [18:0] Wgt_2_352,
input [18:0] Wgt_2_353,
input [18:0] Wgt_2_354,
input [18:0] Wgt_2_355,
input [18:0] Wgt_2_356,
input [18:0] Wgt_2_357,
input [18:0] Wgt_2_358,
input [18:0] Wgt_2_359,
input [18:0] Wgt_2_360,
input [18:0] Wgt_2_361,
input [18:0] Wgt_2_362,
input [18:0] Wgt_2_363,
input [18:0] Wgt_2_364,
input [18:0] Wgt_2_365,
input [18:0] Wgt_2_366,
input [18:0] Wgt_2_367,
input [18:0] Wgt_2_368,
input [18:0] Wgt_2_369,
input [18:0] Wgt_2_370,
input [18:0] Wgt_2_371,
input [18:0] Wgt_2_372,
input [18:0] Wgt_2_373,
input [18:0] Wgt_2_374,
input [18:0] Wgt_2_375,
input [18:0] Wgt_2_376,
input [18:0] Wgt_2_377,
input [18:0] Wgt_2_378,
input [18:0] Wgt_2_379,
input [18:0] Wgt_2_380,
input [18:0] Wgt_2_381,
input [18:0] Wgt_2_382,
input [18:0] Wgt_2_383,
input [18:0] Wgt_2_384,
input [18:0] Wgt_2_385,
input [18:0] Wgt_2_386,
input [18:0] Wgt_2_387,
input [18:0] Wgt_2_388,
input [18:0] Wgt_2_389,
input [18:0] Wgt_2_390,
input [18:0] Wgt_2_391,
input [18:0] Wgt_2_392,
input [18:0] Wgt_2_393,
input [18:0] Wgt_2_394,
input [18:0] Wgt_2_395,
input [18:0] Wgt_2_396,
input [18:0] Wgt_2_397,
input [18:0] Wgt_2_398,
input [18:0] Wgt_2_399,
input [18:0] Wgt_2_400,
input [18:0] Wgt_2_401,
input [18:0] Wgt_2_402,
input [18:0] Wgt_2_403,
input [18:0] Wgt_2_404,
input [18:0] Wgt_2_405,
input [18:0] Wgt_2_406,
input [18:0] Wgt_2_407,
input [18:0] Wgt_2_408,
input [18:0] Wgt_2_409,
input [18:0] Wgt_2_410,
input [18:0] Wgt_2_411,
input [18:0] Wgt_2_412,
input [18:0] Wgt_2_413,
input [18:0] Wgt_2_414,
input [18:0] Wgt_2_415,
input [18:0] Wgt_2_416,
input [18:0] Wgt_2_417,
input [18:0] Wgt_2_418,
input [18:0] Wgt_2_419,
input [18:0] Wgt_2_420,
input [18:0] Wgt_2_421,
input [18:0] Wgt_2_422,
input [18:0] Wgt_2_423,
input [18:0] Wgt_2_424,
input [18:0] Wgt_2_425,
input [18:0] Wgt_2_426,
input [18:0] Wgt_2_427,
input [18:0] Wgt_2_428,
input [18:0] Wgt_2_429,
input [18:0] Wgt_2_430,
input [18:0] Wgt_2_431,
input [18:0] Wgt_2_432,
input [18:0] Wgt_2_433,
input [18:0] Wgt_2_434,
input [18:0] Wgt_2_435,
input [18:0] Wgt_2_436,
input [18:0] Wgt_2_437,
input [18:0] Wgt_2_438,
input [18:0] Wgt_2_439,
input [18:0] Wgt_2_440,
input [18:0] Wgt_2_441,
input [18:0] Wgt_2_442,
input [18:0] Wgt_2_443,
input [18:0] Wgt_2_444,
input [18:0] Wgt_2_445,
input [18:0] Wgt_2_446,
input [18:0] Wgt_2_447,
input [18:0] Wgt_2_448,
input [18:0] Wgt_2_449,
input [18:0] Wgt_2_450,
input [18:0] Wgt_2_451,
input [18:0] Wgt_2_452,
input [18:0] Wgt_2_453,
input [18:0] Wgt_2_454,
input [18:0] Wgt_2_455,
input [18:0] Wgt_2_456,
input [18:0] Wgt_2_457,
input [18:0] Wgt_2_458,
input [18:0] Wgt_2_459,
input [18:0] Wgt_2_460,
input [18:0] Wgt_2_461,
input [18:0] Wgt_2_462,
input [18:0] Wgt_2_463,
input [18:0] Wgt_2_464,
input [18:0] Wgt_2_465,
input [18:0] Wgt_2_466,
input [18:0] Wgt_2_467,
input [18:0] Wgt_2_468,
input [18:0] Wgt_2_469,
input [18:0] Wgt_2_470,
input [18:0] Wgt_2_471,
input [18:0] Wgt_2_472,
input [18:0] Wgt_2_473,
input [18:0] Wgt_2_474,
input [18:0] Wgt_2_475,
input [18:0] Wgt_2_476,
input [18:0] Wgt_2_477,
input [18:0] Wgt_2_478,
input [18:0] Wgt_2_479,
input [18:0] Wgt_2_480,
input [18:0] Wgt_2_481,
input [18:0] Wgt_2_482,
input [18:0] Wgt_2_483,
input [18:0] Wgt_2_484,
input [18:0] Wgt_2_485,
input [18:0] Wgt_2_486,
input [18:0] Wgt_2_487,
input [18:0] Wgt_2_488,
input [18:0] Wgt_2_489,
input [18:0] Wgt_2_490,
input [18:0] Wgt_2_491,
input [18:0] Wgt_2_492,
input [18:0] Wgt_2_493,
input [18:0] Wgt_2_494,
input [18:0] Wgt_2_495,
input [18:0] Wgt_2_496,
input [18:0] Wgt_2_497,
input [18:0] Wgt_2_498,
input [18:0] Wgt_2_499,
input [18:0] Wgt_2_500,
input [18:0] Wgt_2_501,
input [18:0] Wgt_2_502,
input [18:0] Wgt_2_503,
input [18:0] Wgt_2_504,
input [18:0] Wgt_2_505,
input [18:0] Wgt_2_506,
input [18:0] Wgt_2_507,
input [18:0] Wgt_2_508,
input [18:0] Wgt_2_509,
input [18:0] Wgt_2_510,
input [18:0] Wgt_2_511,
input [18:0] Wgt_2_512,
input [18:0] Wgt_2_513,
input [18:0] Wgt_2_514,
input [18:0] Wgt_2_515,
input [18:0] Wgt_2_516,
input [18:0] Wgt_2_517,
input [18:0] Wgt_2_518,
input [18:0] Wgt_2_519,
input [18:0] Wgt_2_520,
input [18:0] Wgt_2_521,
input [18:0] Wgt_2_522,
input [18:0] Wgt_2_523,
input [18:0] Wgt_2_524,
input [18:0] Wgt_2_525,
input [18:0] Wgt_2_526,
input [18:0] Wgt_2_527,
input [18:0] Wgt_2_528,
input [18:0] Wgt_2_529,
input [18:0] Wgt_2_530,
input [18:0] Wgt_2_531,
input [18:0] Wgt_2_532,
input [18:0] Wgt_2_533,
input [18:0] Wgt_2_534,
input [18:0] Wgt_2_535,
input [18:0] Wgt_2_536,
input [18:0] Wgt_2_537,
input [18:0] Wgt_2_538,
input [18:0] Wgt_2_539,
input [18:0] Wgt_2_540,
input [18:0] Wgt_2_541,
input [18:0] Wgt_2_542,
input [18:0] Wgt_2_543,
input [18:0] Wgt_2_544,
input [18:0] Wgt_2_545,
input [18:0] Wgt_2_546,
input [18:0] Wgt_2_547,
input [18:0] Wgt_2_548,
input [18:0] Wgt_2_549,
input [18:0] Wgt_2_550,
input [18:0] Wgt_2_551,
input [18:0] Wgt_2_552,
input [18:0] Wgt_2_553,
input [18:0] Wgt_2_554,
input [18:0] Wgt_2_555,
input [18:0] Wgt_2_556,
input [18:0] Wgt_2_557,
input [18:0] Wgt_2_558,
input [18:0] Wgt_2_559,
input [18:0] Wgt_2_560,
input [18:0] Wgt_2_561,
input [18:0] Wgt_2_562,
input [18:0] Wgt_2_563,
input [18:0] Wgt_2_564,
input [18:0] Wgt_2_565,
input [18:0] Wgt_2_566,
input [18:0] Wgt_2_567,
input [18:0] Wgt_2_568,
input [18:0] Wgt_2_569,
input [18:0] Wgt_2_570,
input [18:0] Wgt_2_571,
input [18:0] Wgt_2_572,
input [18:0] Wgt_2_573,
input [18:0] Wgt_2_574,
input [18:0] Wgt_2_575,
input [18:0] Wgt_2_576,
input [18:0] Wgt_2_577,
input [18:0] Wgt_2_578,
input [18:0] Wgt_2_579,
input [18:0] Wgt_2_580,
input [18:0] Wgt_2_581,
input [18:0] Wgt_2_582,
input [18:0] Wgt_2_583,
input [18:0] Wgt_2_584,
input [18:0] Wgt_2_585,
input [18:0] Wgt_2_586,
input [18:0] Wgt_2_587,
input [18:0] Wgt_2_588,
input [18:0] Wgt_2_589,
input [18:0] Wgt_2_590,
input [18:0] Wgt_2_591,
input [18:0] Wgt_2_592,
input [18:0] Wgt_2_593,
input [18:0] Wgt_2_594,
input [18:0] Wgt_2_595,
input [18:0] Wgt_2_596,
input [18:0] Wgt_2_597,
input [18:0] Wgt_2_598,
input [18:0] Wgt_2_599,
input [18:0] Wgt_2_600,
input [18:0] Wgt_2_601,
input [18:0] Wgt_2_602,
input [18:0] Wgt_2_603,
input [18:0] Wgt_2_604,
input [18:0] Wgt_2_605,
input [18:0] Wgt_2_606,
input [18:0] Wgt_2_607,
input [18:0] Wgt_2_608,
input [18:0] Wgt_2_609,
input [18:0] Wgt_2_610,
input [18:0] Wgt_2_611,
input [18:0] Wgt_2_612,
input [18:0] Wgt_2_613,
input [18:0] Wgt_2_614,
input [18:0] Wgt_2_615,
input [18:0] Wgt_2_616,
input [18:0] Wgt_2_617,
input [18:0] Wgt_2_618,
input [18:0] Wgt_2_619,
input [18:0] Wgt_2_620,
input [18:0] Wgt_2_621,
input [18:0] Wgt_2_622,
input [18:0] Wgt_2_623,
input [18:0] Wgt_2_624,
input [18:0] Wgt_2_625,
input [18:0] Wgt_2_626,
input [18:0] Wgt_2_627,
input [18:0] Wgt_2_628,
input [18:0] Wgt_2_629,
input [18:0] Wgt_2_630,
input [18:0] Wgt_2_631,
input [18:0] Wgt_2_632,
input [18:0] Wgt_2_633,
input [18:0] Wgt_2_634,
input [18:0] Wgt_2_635,
input [18:0] Wgt_2_636,
input [18:0] Wgt_2_637,
input [18:0] Wgt_2_638,
input [18:0] Wgt_2_639,
input [18:0] Wgt_2_640,
input [18:0] Wgt_2_641,
input [18:0] Wgt_2_642,
input [18:0] Wgt_2_643,
input [18:0] Wgt_2_644,
input [18:0] Wgt_2_645,
input [18:0] Wgt_2_646,
input [18:0] Wgt_2_647,
input [18:0] Wgt_2_648,
input [18:0] Wgt_2_649,
input [18:0] Wgt_2_650,
input [18:0] Wgt_2_651,
input [18:0] Wgt_2_652,
input [18:0] Wgt_2_653,
input [18:0] Wgt_2_654,
input [18:0] Wgt_2_655,
input [18:0] Wgt_2_656,
input [18:0] Wgt_2_657,
input [18:0] Wgt_2_658,
input [18:0] Wgt_2_659,
input [18:0] Wgt_2_660,
input [18:0] Wgt_2_661,
input [18:0] Wgt_2_662,
input [18:0] Wgt_2_663,
input [18:0] Wgt_2_664,
input [18:0] Wgt_2_665,
input [18:0] Wgt_2_666,
input [18:0] Wgt_2_667,
input [18:0] Wgt_2_668,
input [18:0] Wgt_2_669,
input [18:0] Wgt_2_670,
input [18:0] Wgt_2_671,
input [18:0] Wgt_2_672,
input [18:0] Wgt_2_673,
input [18:0] Wgt_2_674,
input [18:0] Wgt_2_675,
input [18:0] Wgt_2_676,
input [18:0] Wgt_2_677,
input [18:0] Wgt_2_678,
input [18:0] Wgt_2_679,
input [18:0] Wgt_2_680,
input [18:0] Wgt_2_681,
input [18:0] Wgt_2_682,
input [18:0] Wgt_2_683,
input [18:0] Wgt_2_684,
input [18:0] Wgt_2_685,
input [18:0] Wgt_2_686,
input [18:0] Wgt_2_687,
input [18:0] Wgt_2_688,
input [18:0] Wgt_2_689,
input [18:0] Wgt_2_690,
input [18:0] Wgt_2_691,
input [18:0] Wgt_2_692,
input [18:0] Wgt_2_693,
input [18:0] Wgt_2_694,
input [18:0] Wgt_2_695,
input [18:0] Wgt_2_696,
input [18:0] Wgt_2_697,
input [18:0] Wgt_2_698,
input [18:0] Wgt_2_699,
input [18:0] Wgt_2_700,
input [18:0] Wgt_2_701,
input [18:0] Wgt_2_702,
input [18:0] Wgt_2_703,
input [18:0] Wgt_2_704,
input [18:0] Wgt_2_705,
input [18:0] Wgt_2_706,
input [18:0] Wgt_2_707,
input [18:0] Wgt_2_708,
input [18:0] Wgt_2_709,
input [18:0] Wgt_2_710,
input [18:0] Wgt_2_711,
input [18:0] Wgt_2_712,
input [18:0] Wgt_2_713,
input [18:0] Wgt_2_714,
input [18:0] Wgt_2_715,
input [18:0] Wgt_2_716,
input [18:0] Wgt_2_717,
input [18:0] Wgt_2_718,
input [18:0] Wgt_2_719,
input [18:0] Wgt_2_720,
input [18:0] Wgt_2_721,
input [18:0] Wgt_2_722,
input [18:0] Wgt_2_723,
input [18:0] Wgt_2_724,
input [18:0] Wgt_2_725,
input [18:0] Wgt_2_726,
input [18:0] Wgt_2_727,
input [18:0] Wgt_2_728,
input [18:0] Wgt_2_729,
input [18:0] Wgt_2_730,
input [18:0] Wgt_2_731,
input [18:0] Wgt_2_732,
input [18:0] Wgt_2_733,
input [18:0] Wgt_2_734,
input [18:0] Wgt_2_735,
input [18:0] Wgt_2_736,
input [18:0] Wgt_2_737,
input [18:0] Wgt_2_738,
input [18:0] Wgt_2_739,
input [18:0] Wgt_2_740,
input [18:0] Wgt_2_741,
input [18:0] Wgt_2_742,
input [18:0] Wgt_2_743,
input [18:0] Wgt_2_744,
input [18:0] Wgt_2_745,
input [18:0] Wgt_2_746,
input [18:0] Wgt_2_747,
input [18:0] Wgt_2_748,
input [18:0] Wgt_2_749,
input [18:0] Wgt_2_750,
input [18:0] Wgt_2_751,
input [18:0] Wgt_2_752,
input [18:0] Wgt_2_753,
input [18:0] Wgt_2_754,
input [18:0] Wgt_2_755,
input [18:0] Wgt_2_756,
input [18:0] Wgt_2_757,
input [18:0] Wgt_2_758,
input [18:0] Wgt_2_759,
input [18:0] Wgt_2_760,
input [18:0] Wgt_2_761,
input [18:0] Wgt_2_762,
input [18:0] Wgt_2_763,
input [18:0] Wgt_2_764,
input [18:0] Wgt_2_765,
input [18:0] Wgt_2_766,
input [18:0] Wgt_2_767,
input [18:0] Wgt_2_768,
input [18:0] Wgt_2_769,
input [18:0] Wgt_2_770,
input [18:0] Wgt_2_771,
input [18:0] Wgt_2_772,
input [18:0] Wgt_2_773,
input [18:0] Wgt_2_774,
input [18:0] Wgt_2_775,
input [18:0] Wgt_2_776,
input [18:0] Wgt_2_777,
input [18:0] Wgt_2_778,
input [18:0] Wgt_2_779,
input [18:0] Wgt_2_780,
input [18:0] Wgt_2_781,
input [18:0] Wgt_2_782,
input [18:0] Wgt_2_783,
input [18:0] Wgt_2_784,
input [18:0] Wgt_3_0,
input [18:0] Wgt_3_1,
input [18:0] Wgt_3_2,
input [18:0] Wgt_3_3,
input [18:0] Wgt_3_4,
input [18:0] Wgt_3_5,
input [18:0] Wgt_3_6,
input [18:0] Wgt_3_7,
input [18:0] Wgt_3_8,
input [18:0] Wgt_3_9,
input [18:0] Wgt_3_10,
input [18:0] Wgt_3_11,
input [18:0] Wgt_3_12,
input [18:0] Wgt_3_13,
input [18:0] Wgt_3_14,
input [18:0] Wgt_3_15,
input [18:0] Wgt_3_16,
input [18:0] Wgt_3_17,
input [18:0] Wgt_3_18,
input [18:0] Wgt_3_19,
input [18:0] Wgt_3_20,
input [18:0] Wgt_3_21,
input [18:0] Wgt_3_22,
input [18:0] Wgt_3_23,
input [18:0] Wgt_3_24,
input [18:0] Wgt_3_25,
input [18:0] Wgt_3_26,
input [18:0] Wgt_3_27,
input [18:0] Wgt_3_28,
input [18:0] Wgt_3_29,
input [18:0] Wgt_3_30,
input [18:0] Wgt_3_31,
input [18:0] Wgt_3_32,
input [18:0] Wgt_3_33,
input [18:0] Wgt_3_34,
input [18:0] Wgt_3_35,
input [18:0] Wgt_3_36,
input [18:0] Wgt_3_37,
input [18:0] Wgt_3_38,
input [18:0] Wgt_3_39,
input [18:0] Wgt_3_40,
input [18:0] Wgt_3_41,
input [18:0] Wgt_3_42,
input [18:0] Wgt_3_43,
input [18:0] Wgt_3_44,
input [18:0] Wgt_3_45,
input [18:0] Wgt_3_46,
input [18:0] Wgt_3_47,
input [18:0] Wgt_3_48,
input [18:0] Wgt_3_49,
input [18:0] Wgt_3_50,
input [18:0] Wgt_3_51,
input [18:0] Wgt_3_52,
input [18:0] Wgt_3_53,
input [18:0] Wgt_3_54,
input [18:0] Wgt_3_55,
input [18:0] Wgt_3_56,
input [18:0] Wgt_3_57,
input [18:0] Wgt_3_58,
input [18:0] Wgt_3_59,
input [18:0] Wgt_3_60,
input [18:0] Wgt_3_61,
input [18:0] Wgt_3_62,
input [18:0] Wgt_3_63,
input [18:0] Wgt_3_64,
input [18:0] Wgt_3_65,
input [18:0] Wgt_3_66,
input [18:0] Wgt_3_67,
input [18:0] Wgt_3_68,
input [18:0] Wgt_3_69,
input [18:0] Wgt_3_70,
input [18:0] Wgt_3_71,
input [18:0] Wgt_3_72,
input [18:0] Wgt_3_73,
input [18:0] Wgt_3_74,
input [18:0] Wgt_3_75,
input [18:0] Wgt_3_76,
input [18:0] Wgt_3_77,
input [18:0] Wgt_3_78,
input [18:0] Wgt_3_79,
input [18:0] Wgt_3_80,
input [18:0] Wgt_3_81,
input [18:0] Wgt_3_82,
input [18:0] Wgt_3_83,
input [18:0] Wgt_3_84,
input [18:0] Wgt_3_85,
input [18:0] Wgt_3_86,
input [18:0] Wgt_3_87,
input [18:0] Wgt_3_88,
input [18:0] Wgt_3_89,
input [18:0] Wgt_3_90,
input [18:0] Wgt_3_91,
input [18:0] Wgt_3_92,
input [18:0] Wgt_3_93,
input [18:0] Wgt_3_94,
input [18:0] Wgt_3_95,
input [18:0] Wgt_3_96,
input [18:0] Wgt_3_97,
input [18:0] Wgt_3_98,
input [18:0] Wgt_3_99,
input [18:0] Wgt_3_100,
input [18:0] Wgt_3_101,
input [18:0] Wgt_3_102,
input [18:0] Wgt_3_103,
input [18:0] Wgt_3_104,
input [18:0] Wgt_3_105,
input [18:0] Wgt_3_106,
input [18:0] Wgt_3_107,
input [18:0] Wgt_3_108,
input [18:0] Wgt_3_109,
input [18:0] Wgt_3_110,
input [18:0] Wgt_3_111,
input [18:0] Wgt_3_112,
input [18:0] Wgt_3_113,
input [18:0] Wgt_3_114,
input [18:0] Wgt_3_115,
input [18:0] Wgt_3_116,
input [18:0] Wgt_3_117,
input [18:0] Wgt_3_118,
input [18:0] Wgt_3_119,
input [18:0] Wgt_3_120,
input [18:0] Wgt_3_121,
input [18:0] Wgt_3_122,
input [18:0] Wgt_3_123,
input [18:0] Wgt_3_124,
input [18:0] Wgt_3_125,
input [18:0] Wgt_3_126,
input [18:0] Wgt_3_127,
input [18:0] Wgt_3_128,
input [18:0] Wgt_3_129,
input [18:0] Wgt_3_130,
input [18:0] Wgt_3_131,
input [18:0] Wgt_3_132,
input [18:0] Wgt_3_133,
input [18:0] Wgt_3_134,
input [18:0] Wgt_3_135,
input [18:0] Wgt_3_136,
input [18:0] Wgt_3_137,
input [18:0] Wgt_3_138,
input [18:0] Wgt_3_139,
input [18:0] Wgt_3_140,
input [18:0] Wgt_3_141,
input [18:0] Wgt_3_142,
input [18:0] Wgt_3_143,
input [18:0] Wgt_3_144,
input [18:0] Wgt_3_145,
input [18:0] Wgt_3_146,
input [18:0] Wgt_3_147,
input [18:0] Wgt_3_148,
input [18:0] Wgt_3_149,
input [18:0] Wgt_3_150,
input [18:0] Wgt_3_151,
input [18:0] Wgt_3_152,
input [18:0] Wgt_3_153,
input [18:0] Wgt_3_154,
input [18:0] Wgt_3_155,
input [18:0] Wgt_3_156,
input [18:0] Wgt_3_157,
input [18:0] Wgt_3_158,
input [18:0] Wgt_3_159,
input [18:0] Wgt_3_160,
input [18:0] Wgt_3_161,
input [18:0] Wgt_3_162,
input [18:0] Wgt_3_163,
input [18:0] Wgt_3_164,
input [18:0] Wgt_3_165,
input [18:0] Wgt_3_166,
input [18:0] Wgt_3_167,
input [18:0] Wgt_3_168,
input [18:0] Wgt_3_169,
input [18:0] Wgt_3_170,
input [18:0] Wgt_3_171,
input [18:0] Wgt_3_172,
input [18:0] Wgt_3_173,
input [18:0] Wgt_3_174,
input [18:0] Wgt_3_175,
input [18:0] Wgt_3_176,
input [18:0] Wgt_3_177,
input [18:0] Wgt_3_178,
input [18:0] Wgt_3_179,
input [18:0] Wgt_3_180,
input [18:0] Wgt_3_181,
input [18:0] Wgt_3_182,
input [18:0] Wgt_3_183,
input [18:0] Wgt_3_184,
input [18:0] Wgt_3_185,
input [18:0] Wgt_3_186,
input [18:0] Wgt_3_187,
input [18:0] Wgt_3_188,
input [18:0] Wgt_3_189,
input [18:0] Wgt_3_190,
input [18:0] Wgt_3_191,
input [18:0] Wgt_3_192,
input [18:0] Wgt_3_193,
input [18:0] Wgt_3_194,
input [18:0] Wgt_3_195,
input [18:0] Wgt_3_196,
input [18:0] Wgt_3_197,
input [18:0] Wgt_3_198,
input [18:0] Wgt_3_199,
input [18:0] Wgt_3_200,
input [18:0] Wgt_3_201,
input [18:0] Wgt_3_202,
input [18:0] Wgt_3_203,
input [18:0] Wgt_3_204,
input [18:0] Wgt_3_205,
input [18:0] Wgt_3_206,
input [18:0] Wgt_3_207,
input [18:0] Wgt_3_208,
input [18:0] Wgt_3_209,
input [18:0] Wgt_3_210,
input [18:0] Wgt_3_211,
input [18:0] Wgt_3_212,
input [18:0] Wgt_3_213,
input [18:0] Wgt_3_214,
input [18:0] Wgt_3_215,
input [18:0] Wgt_3_216,
input [18:0] Wgt_3_217,
input [18:0] Wgt_3_218,
input [18:0] Wgt_3_219,
input [18:0] Wgt_3_220,
input [18:0] Wgt_3_221,
input [18:0] Wgt_3_222,
input [18:0] Wgt_3_223,
input [18:0] Wgt_3_224,
input [18:0] Wgt_3_225,
input [18:0] Wgt_3_226,
input [18:0] Wgt_3_227,
input [18:0] Wgt_3_228,
input [18:0] Wgt_3_229,
input [18:0] Wgt_3_230,
input [18:0] Wgt_3_231,
input [18:0] Wgt_3_232,
input [18:0] Wgt_3_233,
input [18:0] Wgt_3_234,
input [18:0] Wgt_3_235,
input [18:0] Wgt_3_236,
input [18:0] Wgt_3_237,
input [18:0] Wgt_3_238,
input [18:0] Wgt_3_239,
input [18:0] Wgt_3_240,
input [18:0] Wgt_3_241,
input [18:0] Wgt_3_242,
input [18:0] Wgt_3_243,
input [18:0] Wgt_3_244,
input [18:0] Wgt_3_245,
input [18:0] Wgt_3_246,
input [18:0] Wgt_3_247,
input [18:0] Wgt_3_248,
input [18:0] Wgt_3_249,
input [18:0] Wgt_3_250,
input [18:0] Wgt_3_251,
input [18:0] Wgt_3_252,
input [18:0] Wgt_3_253,
input [18:0] Wgt_3_254,
input [18:0] Wgt_3_255,
input [18:0] Wgt_3_256,
input [18:0] Wgt_3_257,
input [18:0] Wgt_3_258,
input [18:0] Wgt_3_259,
input [18:0] Wgt_3_260,
input [18:0] Wgt_3_261,
input [18:0] Wgt_3_262,
input [18:0] Wgt_3_263,
input [18:0] Wgt_3_264,
input [18:0] Wgt_3_265,
input [18:0] Wgt_3_266,
input [18:0] Wgt_3_267,
input [18:0] Wgt_3_268,
input [18:0] Wgt_3_269,
input [18:0] Wgt_3_270,
input [18:0] Wgt_3_271,
input [18:0] Wgt_3_272,
input [18:0] Wgt_3_273,
input [18:0] Wgt_3_274,
input [18:0] Wgt_3_275,
input [18:0] Wgt_3_276,
input [18:0] Wgt_3_277,
input [18:0] Wgt_3_278,
input [18:0] Wgt_3_279,
input [18:0] Wgt_3_280,
input [18:0] Wgt_3_281,
input [18:0] Wgt_3_282,
input [18:0] Wgt_3_283,
input [18:0] Wgt_3_284,
input [18:0] Wgt_3_285,
input [18:0] Wgt_3_286,
input [18:0] Wgt_3_287,
input [18:0] Wgt_3_288,
input [18:0] Wgt_3_289,
input [18:0] Wgt_3_290,
input [18:0] Wgt_3_291,
input [18:0] Wgt_3_292,
input [18:0] Wgt_3_293,
input [18:0] Wgt_3_294,
input [18:0] Wgt_3_295,
input [18:0] Wgt_3_296,
input [18:0] Wgt_3_297,
input [18:0] Wgt_3_298,
input [18:0] Wgt_3_299,
input [18:0] Wgt_3_300,
input [18:0] Wgt_3_301,
input [18:0] Wgt_3_302,
input [18:0] Wgt_3_303,
input [18:0] Wgt_3_304,
input [18:0] Wgt_3_305,
input [18:0] Wgt_3_306,
input [18:0] Wgt_3_307,
input [18:0] Wgt_3_308,
input [18:0] Wgt_3_309,
input [18:0] Wgt_3_310,
input [18:0] Wgt_3_311,
input [18:0] Wgt_3_312,
input [18:0] Wgt_3_313,
input [18:0] Wgt_3_314,
input [18:0] Wgt_3_315,
input [18:0] Wgt_3_316,
input [18:0] Wgt_3_317,
input [18:0] Wgt_3_318,
input [18:0] Wgt_3_319,
input [18:0] Wgt_3_320,
input [18:0] Wgt_3_321,
input [18:0] Wgt_3_322,
input [18:0] Wgt_3_323,
input [18:0] Wgt_3_324,
input [18:0] Wgt_3_325,
input [18:0] Wgt_3_326,
input [18:0] Wgt_3_327,
input [18:0] Wgt_3_328,
input [18:0] Wgt_3_329,
input [18:0] Wgt_3_330,
input [18:0] Wgt_3_331,
input [18:0] Wgt_3_332,
input [18:0] Wgt_3_333,
input [18:0] Wgt_3_334,
input [18:0] Wgt_3_335,
input [18:0] Wgt_3_336,
input [18:0] Wgt_3_337,
input [18:0] Wgt_3_338,
input [18:0] Wgt_3_339,
input [18:0] Wgt_3_340,
input [18:0] Wgt_3_341,
input [18:0] Wgt_3_342,
input [18:0] Wgt_3_343,
input [18:0] Wgt_3_344,
input [18:0] Wgt_3_345,
input [18:0] Wgt_3_346,
input [18:0] Wgt_3_347,
input [18:0] Wgt_3_348,
input [18:0] Wgt_3_349,
input [18:0] Wgt_3_350,
input [18:0] Wgt_3_351,
input [18:0] Wgt_3_352,
input [18:0] Wgt_3_353,
input [18:0] Wgt_3_354,
input [18:0] Wgt_3_355,
input [18:0] Wgt_3_356,
input [18:0] Wgt_3_357,
input [18:0] Wgt_3_358,
input [18:0] Wgt_3_359,
input [18:0] Wgt_3_360,
input [18:0] Wgt_3_361,
input [18:0] Wgt_3_362,
input [18:0] Wgt_3_363,
input [18:0] Wgt_3_364,
input [18:0] Wgt_3_365,
input [18:0] Wgt_3_366,
input [18:0] Wgt_3_367,
input [18:0] Wgt_3_368,
input [18:0] Wgt_3_369,
input [18:0] Wgt_3_370,
input [18:0] Wgt_3_371,
input [18:0] Wgt_3_372,
input [18:0] Wgt_3_373,
input [18:0] Wgt_3_374,
input [18:0] Wgt_3_375,
input [18:0] Wgt_3_376,
input [18:0] Wgt_3_377,
input [18:0] Wgt_3_378,
input [18:0] Wgt_3_379,
input [18:0] Wgt_3_380,
input [18:0] Wgt_3_381,
input [18:0] Wgt_3_382,
input [18:0] Wgt_3_383,
input [18:0] Wgt_3_384,
input [18:0] Wgt_3_385,
input [18:0] Wgt_3_386,
input [18:0] Wgt_3_387,
input [18:0] Wgt_3_388,
input [18:0] Wgt_3_389,
input [18:0] Wgt_3_390,
input [18:0] Wgt_3_391,
input [18:0] Wgt_3_392,
input [18:0] Wgt_3_393,
input [18:0] Wgt_3_394,
input [18:0] Wgt_3_395,
input [18:0] Wgt_3_396,
input [18:0] Wgt_3_397,
input [18:0] Wgt_3_398,
input [18:0] Wgt_3_399,
input [18:0] Wgt_3_400,
input [18:0] Wgt_3_401,
input [18:0] Wgt_3_402,
input [18:0] Wgt_3_403,
input [18:0] Wgt_3_404,
input [18:0] Wgt_3_405,
input [18:0] Wgt_3_406,
input [18:0] Wgt_3_407,
input [18:0] Wgt_3_408,
input [18:0] Wgt_3_409,
input [18:0] Wgt_3_410,
input [18:0] Wgt_3_411,
input [18:0] Wgt_3_412,
input [18:0] Wgt_3_413,
input [18:0] Wgt_3_414,
input [18:0] Wgt_3_415,
input [18:0] Wgt_3_416,
input [18:0] Wgt_3_417,
input [18:0] Wgt_3_418,
input [18:0] Wgt_3_419,
input [18:0] Wgt_3_420,
input [18:0] Wgt_3_421,
input [18:0] Wgt_3_422,
input [18:0] Wgt_3_423,
input [18:0] Wgt_3_424,
input [18:0] Wgt_3_425,
input [18:0] Wgt_3_426,
input [18:0] Wgt_3_427,
input [18:0] Wgt_3_428,
input [18:0] Wgt_3_429,
input [18:0] Wgt_3_430,
input [18:0] Wgt_3_431,
input [18:0] Wgt_3_432,
input [18:0] Wgt_3_433,
input [18:0] Wgt_3_434,
input [18:0] Wgt_3_435,
input [18:0] Wgt_3_436,
input [18:0] Wgt_3_437,
input [18:0] Wgt_3_438,
input [18:0] Wgt_3_439,
input [18:0] Wgt_3_440,
input [18:0] Wgt_3_441,
input [18:0] Wgt_3_442,
input [18:0] Wgt_3_443,
input [18:0] Wgt_3_444,
input [18:0] Wgt_3_445,
input [18:0] Wgt_3_446,
input [18:0] Wgt_3_447,
input [18:0] Wgt_3_448,
input [18:0] Wgt_3_449,
input [18:0] Wgt_3_450,
input [18:0] Wgt_3_451,
input [18:0] Wgt_3_452,
input [18:0] Wgt_3_453,
input [18:0] Wgt_3_454,
input [18:0] Wgt_3_455,
input [18:0] Wgt_3_456,
input [18:0] Wgt_3_457,
input [18:0] Wgt_3_458,
input [18:0] Wgt_3_459,
input [18:0] Wgt_3_460,
input [18:0] Wgt_3_461,
input [18:0] Wgt_3_462,
input [18:0] Wgt_3_463,
input [18:0] Wgt_3_464,
input [18:0] Wgt_3_465,
input [18:0] Wgt_3_466,
input [18:0] Wgt_3_467,
input [18:0] Wgt_3_468,
input [18:0] Wgt_3_469,
input [18:0] Wgt_3_470,
input [18:0] Wgt_3_471,
input [18:0] Wgt_3_472,
input [18:0] Wgt_3_473,
input [18:0] Wgt_3_474,
input [18:0] Wgt_3_475,
input [18:0] Wgt_3_476,
input [18:0] Wgt_3_477,
input [18:0] Wgt_3_478,
input [18:0] Wgt_3_479,
input [18:0] Wgt_3_480,
input [18:0] Wgt_3_481,
input [18:0] Wgt_3_482,
input [18:0] Wgt_3_483,
input [18:0] Wgt_3_484,
input [18:0] Wgt_3_485,
input [18:0] Wgt_3_486,
input [18:0] Wgt_3_487,
input [18:0] Wgt_3_488,
input [18:0] Wgt_3_489,
input [18:0] Wgt_3_490,
input [18:0] Wgt_3_491,
input [18:0] Wgt_3_492,
input [18:0] Wgt_3_493,
input [18:0] Wgt_3_494,
input [18:0] Wgt_3_495,
input [18:0] Wgt_3_496,
input [18:0] Wgt_3_497,
input [18:0] Wgt_3_498,
input [18:0] Wgt_3_499,
input [18:0] Wgt_3_500,
input [18:0] Wgt_3_501,
input [18:0] Wgt_3_502,
input [18:0] Wgt_3_503,
input [18:0] Wgt_3_504,
input [18:0] Wgt_3_505,
input [18:0] Wgt_3_506,
input [18:0] Wgt_3_507,
input [18:0] Wgt_3_508,
input [18:0] Wgt_3_509,
input [18:0] Wgt_3_510,
input [18:0] Wgt_3_511,
input [18:0] Wgt_3_512,
input [18:0] Wgt_3_513,
input [18:0] Wgt_3_514,
input [18:0] Wgt_3_515,
input [18:0] Wgt_3_516,
input [18:0] Wgt_3_517,
input [18:0] Wgt_3_518,
input [18:0] Wgt_3_519,
input [18:0] Wgt_3_520,
input [18:0] Wgt_3_521,
input [18:0] Wgt_3_522,
input [18:0] Wgt_3_523,
input [18:0] Wgt_3_524,
input [18:0] Wgt_3_525,
input [18:0] Wgt_3_526,
input [18:0] Wgt_3_527,
input [18:0] Wgt_3_528,
input [18:0] Wgt_3_529,
input [18:0] Wgt_3_530,
input [18:0] Wgt_3_531,
input [18:0] Wgt_3_532,
input [18:0] Wgt_3_533,
input [18:0] Wgt_3_534,
input [18:0] Wgt_3_535,
input [18:0] Wgt_3_536,
input [18:0] Wgt_3_537,
input [18:0] Wgt_3_538,
input [18:0] Wgt_3_539,
input [18:0] Wgt_3_540,
input [18:0] Wgt_3_541,
input [18:0] Wgt_3_542,
input [18:0] Wgt_3_543,
input [18:0] Wgt_3_544,
input [18:0] Wgt_3_545,
input [18:0] Wgt_3_546,
input [18:0] Wgt_3_547,
input [18:0] Wgt_3_548,
input [18:0] Wgt_3_549,
input [18:0] Wgt_3_550,
input [18:0] Wgt_3_551,
input [18:0] Wgt_3_552,
input [18:0] Wgt_3_553,
input [18:0] Wgt_3_554,
input [18:0] Wgt_3_555,
input [18:0] Wgt_3_556,
input [18:0] Wgt_3_557,
input [18:0] Wgt_3_558,
input [18:0] Wgt_3_559,
input [18:0] Wgt_3_560,
input [18:0] Wgt_3_561,
input [18:0] Wgt_3_562,
input [18:0] Wgt_3_563,
input [18:0] Wgt_3_564,
input [18:0] Wgt_3_565,
input [18:0] Wgt_3_566,
input [18:0] Wgt_3_567,
input [18:0] Wgt_3_568,
input [18:0] Wgt_3_569,
input [18:0] Wgt_3_570,
input [18:0] Wgt_3_571,
input [18:0] Wgt_3_572,
input [18:0] Wgt_3_573,
input [18:0] Wgt_3_574,
input [18:0] Wgt_3_575,
input [18:0] Wgt_3_576,
input [18:0] Wgt_3_577,
input [18:0] Wgt_3_578,
input [18:0] Wgt_3_579,
input [18:0] Wgt_3_580,
input [18:0] Wgt_3_581,
input [18:0] Wgt_3_582,
input [18:0] Wgt_3_583,
input [18:0] Wgt_3_584,
input [18:0] Wgt_3_585,
input [18:0] Wgt_3_586,
input [18:0] Wgt_3_587,
input [18:0] Wgt_3_588,
input [18:0] Wgt_3_589,
input [18:0] Wgt_3_590,
input [18:0] Wgt_3_591,
input [18:0] Wgt_3_592,
input [18:0] Wgt_3_593,
input [18:0] Wgt_3_594,
input [18:0] Wgt_3_595,
input [18:0] Wgt_3_596,
input [18:0] Wgt_3_597,
input [18:0] Wgt_3_598,
input [18:0] Wgt_3_599,
input [18:0] Wgt_3_600,
input [18:0] Wgt_3_601,
input [18:0] Wgt_3_602,
input [18:0] Wgt_3_603,
input [18:0] Wgt_3_604,
input [18:0] Wgt_3_605,
input [18:0] Wgt_3_606,
input [18:0] Wgt_3_607,
input [18:0] Wgt_3_608,
input [18:0] Wgt_3_609,
input [18:0] Wgt_3_610,
input [18:0] Wgt_3_611,
input [18:0] Wgt_3_612,
input [18:0] Wgt_3_613,
input [18:0] Wgt_3_614,
input [18:0] Wgt_3_615,
input [18:0] Wgt_3_616,
input [18:0] Wgt_3_617,
input [18:0] Wgt_3_618,
input [18:0] Wgt_3_619,
input [18:0] Wgt_3_620,
input [18:0] Wgt_3_621,
input [18:0] Wgt_3_622,
input [18:0] Wgt_3_623,
input [18:0] Wgt_3_624,
input [18:0] Wgt_3_625,
input [18:0] Wgt_3_626,
input [18:0] Wgt_3_627,
input [18:0] Wgt_3_628,
input [18:0] Wgt_3_629,
input [18:0] Wgt_3_630,
input [18:0] Wgt_3_631,
input [18:0] Wgt_3_632,
input [18:0] Wgt_3_633,
input [18:0] Wgt_3_634,
input [18:0] Wgt_3_635,
input [18:0] Wgt_3_636,
input [18:0] Wgt_3_637,
input [18:0] Wgt_3_638,
input [18:0] Wgt_3_639,
input [18:0] Wgt_3_640,
input [18:0] Wgt_3_641,
input [18:0] Wgt_3_642,
input [18:0] Wgt_3_643,
input [18:0] Wgt_3_644,
input [18:0] Wgt_3_645,
input [18:0] Wgt_3_646,
input [18:0] Wgt_3_647,
input [18:0] Wgt_3_648,
input [18:0] Wgt_3_649,
input [18:0] Wgt_3_650,
input [18:0] Wgt_3_651,
input [18:0] Wgt_3_652,
input [18:0] Wgt_3_653,
input [18:0] Wgt_3_654,
input [18:0] Wgt_3_655,
input [18:0] Wgt_3_656,
input [18:0] Wgt_3_657,
input [18:0] Wgt_3_658,
input [18:0] Wgt_3_659,
input [18:0] Wgt_3_660,
input [18:0] Wgt_3_661,
input [18:0] Wgt_3_662,
input [18:0] Wgt_3_663,
input [18:0] Wgt_3_664,
input [18:0] Wgt_3_665,
input [18:0] Wgt_3_666,
input [18:0] Wgt_3_667,
input [18:0] Wgt_3_668,
input [18:0] Wgt_3_669,
input [18:0] Wgt_3_670,
input [18:0] Wgt_3_671,
input [18:0] Wgt_3_672,
input [18:0] Wgt_3_673,
input [18:0] Wgt_3_674,
input [18:0] Wgt_3_675,
input [18:0] Wgt_3_676,
input [18:0] Wgt_3_677,
input [18:0] Wgt_3_678,
input [18:0] Wgt_3_679,
input [18:0] Wgt_3_680,
input [18:0] Wgt_3_681,
input [18:0] Wgt_3_682,
input [18:0] Wgt_3_683,
input [18:0] Wgt_3_684,
input [18:0] Wgt_3_685,
input [18:0] Wgt_3_686,
input [18:0] Wgt_3_687,
input [18:0] Wgt_3_688,
input [18:0] Wgt_3_689,
input [18:0] Wgt_3_690,
input [18:0] Wgt_3_691,
input [18:0] Wgt_3_692,
input [18:0] Wgt_3_693,
input [18:0] Wgt_3_694,
input [18:0] Wgt_3_695,
input [18:0] Wgt_3_696,
input [18:0] Wgt_3_697,
input [18:0] Wgt_3_698,
input [18:0] Wgt_3_699,
input [18:0] Wgt_3_700,
input [18:0] Wgt_3_701,
input [18:0] Wgt_3_702,
input [18:0] Wgt_3_703,
input [18:0] Wgt_3_704,
input [18:0] Wgt_3_705,
input [18:0] Wgt_3_706,
input [18:0] Wgt_3_707,
input [18:0] Wgt_3_708,
input [18:0] Wgt_3_709,
input [18:0] Wgt_3_710,
input [18:0] Wgt_3_711,
input [18:0] Wgt_3_712,
input [18:0] Wgt_3_713,
input [18:0] Wgt_3_714,
input [18:0] Wgt_3_715,
input [18:0] Wgt_3_716,
input [18:0] Wgt_3_717,
input [18:0] Wgt_3_718,
input [18:0] Wgt_3_719,
input [18:0] Wgt_3_720,
input [18:0] Wgt_3_721,
input [18:0] Wgt_3_722,
input [18:0] Wgt_3_723,
input [18:0] Wgt_3_724,
input [18:0] Wgt_3_725,
input [18:0] Wgt_3_726,
input [18:0] Wgt_3_727,
input [18:0] Wgt_3_728,
input [18:0] Wgt_3_729,
input [18:0] Wgt_3_730,
input [18:0] Wgt_3_731,
input [18:0] Wgt_3_732,
input [18:0] Wgt_3_733,
input [18:0] Wgt_3_734,
input [18:0] Wgt_3_735,
input [18:0] Wgt_3_736,
input [18:0] Wgt_3_737,
input [18:0] Wgt_3_738,
input [18:0] Wgt_3_739,
input [18:0] Wgt_3_740,
input [18:0] Wgt_3_741,
input [18:0] Wgt_3_742,
input [18:0] Wgt_3_743,
input [18:0] Wgt_3_744,
input [18:0] Wgt_3_745,
input [18:0] Wgt_3_746,
input [18:0] Wgt_3_747,
input [18:0] Wgt_3_748,
input [18:0] Wgt_3_749,
input [18:0] Wgt_3_750,
input [18:0] Wgt_3_751,
input [18:0] Wgt_3_752,
input [18:0] Wgt_3_753,
input [18:0] Wgt_3_754,
input [18:0] Wgt_3_755,
input [18:0] Wgt_3_756,
input [18:0] Wgt_3_757,
input [18:0] Wgt_3_758,
input [18:0] Wgt_3_759,
input [18:0] Wgt_3_760,
input [18:0] Wgt_3_761,
input [18:0] Wgt_3_762,
input [18:0] Wgt_3_763,
input [18:0] Wgt_3_764,
input [18:0] Wgt_3_765,
input [18:0] Wgt_3_766,
input [18:0] Wgt_3_767,
input [18:0] Wgt_3_768,
input [18:0] Wgt_3_769,
input [18:0] Wgt_3_770,
input [18:0] Wgt_3_771,
input [18:0] Wgt_3_772,
input [18:0] Wgt_3_773,
input [18:0] Wgt_3_774,
input [18:0] Wgt_3_775,
input [18:0] Wgt_3_776,
input [18:0] Wgt_3_777,
input [18:0] Wgt_3_778,
input [18:0] Wgt_3_779,
input [18:0] Wgt_3_780,
input [18:0] Wgt_3_781,
input [18:0] Wgt_3_782,
input [18:0] Wgt_3_783,
input [18:0] Wgt_3_784,
input [18:0] Wgt_4_0,
input [18:0] Wgt_4_1,
input [18:0] Wgt_4_2,
input [18:0] Wgt_4_3,
input [18:0] Wgt_4_4,
input [18:0] Wgt_4_5,
input [18:0] Wgt_4_6,
input [18:0] Wgt_4_7,
input [18:0] Wgt_4_8,
input [18:0] Wgt_4_9,
input [18:0] Wgt_4_10,
input [18:0] Wgt_4_11,
input [18:0] Wgt_4_12,
input [18:0] Wgt_4_13,
input [18:0] Wgt_4_14,
input [18:0] Wgt_4_15,
input [18:0] Wgt_4_16,
input [18:0] Wgt_4_17,
input [18:0] Wgt_4_18,
input [18:0] Wgt_4_19,
input [18:0] Wgt_4_20,
input [18:0] Wgt_4_21,
input [18:0] Wgt_4_22,
input [18:0] Wgt_4_23,
input [18:0] Wgt_4_24,
input [18:0] Wgt_4_25,
input [18:0] Wgt_4_26,
input [18:0] Wgt_4_27,
input [18:0] Wgt_4_28,
input [18:0] Wgt_4_29,
input [18:0] Wgt_4_30,
input [18:0] Wgt_4_31,
input [18:0] Wgt_4_32,
input [18:0] Wgt_4_33,
input [18:0] Wgt_4_34,
input [18:0] Wgt_4_35,
input [18:0] Wgt_4_36,
input [18:0] Wgt_4_37,
input [18:0] Wgt_4_38,
input [18:0] Wgt_4_39,
input [18:0] Wgt_4_40,
input [18:0] Wgt_4_41,
input [18:0] Wgt_4_42,
input [18:0] Wgt_4_43,
input [18:0] Wgt_4_44,
input [18:0] Wgt_4_45,
input [18:0] Wgt_4_46,
input [18:0] Wgt_4_47,
input [18:0] Wgt_4_48,
input [18:0] Wgt_4_49,
input [18:0] Wgt_4_50,
input [18:0] Wgt_4_51,
input [18:0] Wgt_4_52,
input [18:0] Wgt_4_53,
input [18:0] Wgt_4_54,
input [18:0] Wgt_4_55,
input [18:0] Wgt_4_56,
input [18:0] Wgt_4_57,
input [18:0] Wgt_4_58,
input [18:0] Wgt_4_59,
input [18:0] Wgt_4_60,
input [18:0] Wgt_4_61,
input [18:0] Wgt_4_62,
input [18:0] Wgt_4_63,
input [18:0] Wgt_4_64,
input [18:0] Wgt_4_65,
input [18:0] Wgt_4_66,
input [18:0] Wgt_4_67,
input [18:0] Wgt_4_68,
input [18:0] Wgt_4_69,
input [18:0] Wgt_4_70,
input [18:0] Wgt_4_71,
input [18:0] Wgt_4_72,
input [18:0] Wgt_4_73,
input [18:0] Wgt_4_74,
input [18:0] Wgt_4_75,
input [18:0] Wgt_4_76,
input [18:0] Wgt_4_77,
input [18:0] Wgt_4_78,
input [18:0] Wgt_4_79,
input [18:0] Wgt_4_80,
input [18:0] Wgt_4_81,
input [18:0] Wgt_4_82,
input [18:0] Wgt_4_83,
input [18:0] Wgt_4_84,
input [18:0] Wgt_4_85,
input [18:0] Wgt_4_86,
input [18:0] Wgt_4_87,
input [18:0] Wgt_4_88,
input [18:0] Wgt_4_89,
input [18:0] Wgt_4_90,
input [18:0] Wgt_4_91,
input [18:0] Wgt_4_92,
input [18:0] Wgt_4_93,
input [18:0] Wgt_4_94,
input [18:0] Wgt_4_95,
input [18:0] Wgt_4_96,
input [18:0] Wgt_4_97,
input [18:0] Wgt_4_98,
input [18:0] Wgt_4_99,
input [18:0] Wgt_4_100,
input [18:0] Wgt_4_101,
input [18:0] Wgt_4_102,
input [18:0] Wgt_4_103,
input [18:0] Wgt_4_104,
input [18:0] Wgt_4_105,
input [18:0] Wgt_4_106,
input [18:0] Wgt_4_107,
input [18:0] Wgt_4_108,
input [18:0] Wgt_4_109,
input [18:0] Wgt_4_110,
input [18:0] Wgt_4_111,
input [18:0] Wgt_4_112,
input [18:0] Wgt_4_113,
input [18:0] Wgt_4_114,
input [18:0] Wgt_4_115,
input [18:0] Wgt_4_116,
input [18:0] Wgt_4_117,
input [18:0] Wgt_4_118,
input [18:0] Wgt_4_119,
input [18:0] Wgt_4_120,
input [18:0] Wgt_4_121,
input [18:0] Wgt_4_122,
input [18:0] Wgt_4_123,
input [18:0] Wgt_4_124,
input [18:0] Wgt_4_125,
input [18:0] Wgt_4_126,
input [18:0] Wgt_4_127,
input [18:0] Wgt_4_128,
input [18:0] Wgt_4_129,
input [18:0] Wgt_4_130,
input [18:0] Wgt_4_131,
input [18:0] Wgt_4_132,
input [18:0] Wgt_4_133,
input [18:0] Wgt_4_134,
input [18:0] Wgt_4_135,
input [18:0] Wgt_4_136,
input [18:0] Wgt_4_137,
input [18:0] Wgt_4_138,
input [18:0] Wgt_4_139,
input [18:0] Wgt_4_140,
input [18:0] Wgt_4_141,
input [18:0] Wgt_4_142,
input [18:0] Wgt_4_143,
input [18:0] Wgt_4_144,
input [18:0] Wgt_4_145,
input [18:0] Wgt_4_146,
input [18:0] Wgt_4_147,
input [18:0] Wgt_4_148,
input [18:0] Wgt_4_149,
input [18:0] Wgt_4_150,
input [18:0] Wgt_4_151,
input [18:0] Wgt_4_152,
input [18:0] Wgt_4_153,
input [18:0] Wgt_4_154,
input [18:0] Wgt_4_155,
input [18:0] Wgt_4_156,
input [18:0] Wgt_4_157,
input [18:0] Wgt_4_158,
input [18:0] Wgt_4_159,
input [18:0] Wgt_4_160,
input [18:0] Wgt_4_161,
input [18:0] Wgt_4_162,
input [18:0] Wgt_4_163,
input [18:0] Wgt_4_164,
input [18:0] Wgt_4_165,
input [18:0] Wgt_4_166,
input [18:0] Wgt_4_167,
input [18:0] Wgt_4_168,
input [18:0] Wgt_4_169,
input [18:0] Wgt_4_170,
input [18:0] Wgt_4_171,
input [18:0] Wgt_4_172,
input [18:0] Wgt_4_173,
input [18:0] Wgt_4_174,
input [18:0] Wgt_4_175,
input [18:0] Wgt_4_176,
input [18:0] Wgt_4_177,
input [18:0] Wgt_4_178,
input [18:0] Wgt_4_179,
input [18:0] Wgt_4_180,
input [18:0] Wgt_4_181,
input [18:0] Wgt_4_182,
input [18:0] Wgt_4_183,
input [18:0] Wgt_4_184,
input [18:0] Wgt_4_185,
input [18:0] Wgt_4_186,
input [18:0] Wgt_4_187,
input [18:0] Wgt_4_188,
input [18:0] Wgt_4_189,
input [18:0] Wgt_4_190,
input [18:0] Wgt_4_191,
input [18:0] Wgt_4_192,
input [18:0] Wgt_4_193,
input [18:0] Wgt_4_194,
input [18:0] Wgt_4_195,
input [18:0] Wgt_4_196,
input [18:0] Wgt_4_197,
input [18:0] Wgt_4_198,
input [18:0] Wgt_4_199,
input [18:0] Wgt_4_200,
input [18:0] Wgt_4_201,
input [18:0] Wgt_4_202,
input [18:0] Wgt_4_203,
input [18:0] Wgt_4_204,
input [18:0] Wgt_4_205,
input [18:0] Wgt_4_206,
input [18:0] Wgt_4_207,
input [18:0] Wgt_4_208,
input [18:0] Wgt_4_209,
input [18:0] Wgt_4_210,
input [18:0] Wgt_4_211,
input [18:0] Wgt_4_212,
input [18:0] Wgt_4_213,
input [18:0] Wgt_4_214,
input [18:0] Wgt_4_215,
input [18:0] Wgt_4_216,
input [18:0] Wgt_4_217,
input [18:0] Wgt_4_218,
input [18:0] Wgt_4_219,
input [18:0] Wgt_4_220,
input [18:0] Wgt_4_221,
input [18:0] Wgt_4_222,
input [18:0] Wgt_4_223,
input [18:0] Wgt_4_224,
input [18:0] Wgt_4_225,
input [18:0] Wgt_4_226,
input [18:0] Wgt_4_227,
input [18:0] Wgt_4_228,
input [18:0] Wgt_4_229,
input [18:0] Wgt_4_230,
input [18:0] Wgt_4_231,
input [18:0] Wgt_4_232,
input [18:0] Wgt_4_233,
input [18:0] Wgt_4_234,
input [18:0] Wgt_4_235,
input [18:0] Wgt_4_236,
input [18:0] Wgt_4_237,
input [18:0] Wgt_4_238,
input [18:0] Wgt_4_239,
input [18:0] Wgt_4_240,
input [18:0] Wgt_4_241,
input [18:0] Wgt_4_242,
input [18:0] Wgt_4_243,
input [18:0] Wgt_4_244,
input [18:0] Wgt_4_245,
input [18:0] Wgt_4_246,
input [18:0] Wgt_4_247,
input [18:0] Wgt_4_248,
input [18:0] Wgt_4_249,
input [18:0] Wgt_4_250,
input [18:0] Wgt_4_251,
input [18:0] Wgt_4_252,
input [18:0] Wgt_4_253,
input [18:0] Wgt_4_254,
input [18:0] Wgt_4_255,
input [18:0] Wgt_4_256,
input [18:0] Wgt_4_257,
input [18:0] Wgt_4_258,
input [18:0] Wgt_4_259,
input [18:0] Wgt_4_260,
input [18:0] Wgt_4_261,
input [18:0] Wgt_4_262,
input [18:0] Wgt_4_263,
input [18:0] Wgt_4_264,
input [18:0] Wgt_4_265,
input [18:0] Wgt_4_266,
input [18:0] Wgt_4_267,
input [18:0] Wgt_4_268,
input [18:0] Wgt_4_269,
input [18:0] Wgt_4_270,
input [18:0] Wgt_4_271,
input [18:0] Wgt_4_272,
input [18:0] Wgt_4_273,
input [18:0] Wgt_4_274,
input [18:0] Wgt_4_275,
input [18:0] Wgt_4_276,
input [18:0] Wgt_4_277,
input [18:0] Wgt_4_278,
input [18:0] Wgt_4_279,
input [18:0] Wgt_4_280,
input [18:0] Wgt_4_281,
input [18:0] Wgt_4_282,
input [18:0] Wgt_4_283,
input [18:0] Wgt_4_284,
input [18:0] Wgt_4_285,
input [18:0] Wgt_4_286,
input [18:0] Wgt_4_287,
input [18:0] Wgt_4_288,
input [18:0] Wgt_4_289,
input [18:0] Wgt_4_290,
input [18:0] Wgt_4_291,
input [18:0] Wgt_4_292,
input [18:0] Wgt_4_293,
input [18:0] Wgt_4_294,
input [18:0] Wgt_4_295,
input [18:0] Wgt_4_296,
input [18:0] Wgt_4_297,
input [18:0] Wgt_4_298,
input [18:0] Wgt_4_299,
input [18:0] Wgt_4_300,
input [18:0] Wgt_4_301,
input [18:0] Wgt_4_302,
input [18:0] Wgt_4_303,
input [18:0] Wgt_4_304,
input [18:0] Wgt_4_305,
input [18:0] Wgt_4_306,
input [18:0] Wgt_4_307,
input [18:0] Wgt_4_308,
input [18:0] Wgt_4_309,
input [18:0] Wgt_4_310,
input [18:0] Wgt_4_311,
input [18:0] Wgt_4_312,
input [18:0] Wgt_4_313,
input [18:0] Wgt_4_314,
input [18:0] Wgt_4_315,
input [18:0] Wgt_4_316,
input [18:0] Wgt_4_317,
input [18:0] Wgt_4_318,
input [18:0] Wgt_4_319,
input [18:0] Wgt_4_320,
input [18:0] Wgt_4_321,
input [18:0] Wgt_4_322,
input [18:0] Wgt_4_323,
input [18:0] Wgt_4_324,
input [18:0] Wgt_4_325,
input [18:0] Wgt_4_326,
input [18:0] Wgt_4_327,
input [18:0] Wgt_4_328,
input [18:0] Wgt_4_329,
input [18:0] Wgt_4_330,
input [18:0] Wgt_4_331,
input [18:0] Wgt_4_332,
input [18:0] Wgt_4_333,
input [18:0] Wgt_4_334,
input [18:0] Wgt_4_335,
input [18:0] Wgt_4_336,
input [18:0] Wgt_4_337,
input [18:0] Wgt_4_338,
input [18:0] Wgt_4_339,
input [18:0] Wgt_4_340,
input [18:0] Wgt_4_341,
input [18:0] Wgt_4_342,
input [18:0] Wgt_4_343,
input [18:0] Wgt_4_344,
input [18:0] Wgt_4_345,
input [18:0] Wgt_4_346,
input [18:0] Wgt_4_347,
input [18:0] Wgt_4_348,
input [18:0] Wgt_4_349,
input [18:0] Wgt_4_350,
input [18:0] Wgt_4_351,
input [18:0] Wgt_4_352,
input [18:0] Wgt_4_353,
input [18:0] Wgt_4_354,
input [18:0] Wgt_4_355,
input [18:0] Wgt_4_356,
input [18:0] Wgt_4_357,
input [18:0] Wgt_4_358,
input [18:0] Wgt_4_359,
input [18:0] Wgt_4_360,
input [18:0] Wgt_4_361,
input [18:0] Wgt_4_362,
input [18:0] Wgt_4_363,
input [18:0] Wgt_4_364,
input [18:0] Wgt_4_365,
input [18:0] Wgt_4_366,
input [18:0] Wgt_4_367,
input [18:0] Wgt_4_368,
input [18:0] Wgt_4_369,
input [18:0] Wgt_4_370,
input [18:0] Wgt_4_371,
input [18:0] Wgt_4_372,
input [18:0] Wgt_4_373,
input [18:0] Wgt_4_374,
input [18:0] Wgt_4_375,
input [18:0] Wgt_4_376,
input [18:0] Wgt_4_377,
input [18:0] Wgt_4_378,
input [18:0] Wgt_4_379,
input [18:0] Wgt_4_380,
input [18:0] Wgt_4_381,
input [18:0] Wgt_4_382,
input [18:0] Wgt_4_383,
input [18:0] Wgt_4_384,
input [18:0] Wgt_4_385,
input [18:0] Wgt_4_386,
input [18:0] Wgt_4_387,
input [18:0] Wgt_4_388,
input [18:0] Wgt_4_389,
input [18:0] Wgt_4_390,
input [18:0] Wgt_4_391,
input [18:0] Wgt_4_392,
input [18:0] Wgt_4_393,
input [18:0] Wgt_4_394,
input [18:0] Wgt_4_395,
input [18:0] Wgt_4_396,
input [18:0] Wgt_4_397,
input [18:0] Wgt_4_398,
input [18:0] Wgt_4_399,
input [18:0] Wgt_4_400,
input [18:0] Wgt_4_401,
input [18:0] Wgt_4_402,
input [18:0] Wgt_4_403,
input [18:0] Wgt_4_404,
input [18:0] Wgt_4_405,
input [18:0] Wgt_4_406,
input [18:0] Wgt_4_407,
input [18:0] Wgt_4_408,
input [18:0] Wgt_4_409,
input [18:0] Wgt_4_410,
input [18:0] Wgt_4_411,
input [18:0] Wgt_4_412,
input [18:0] Wgt_4_413,
input [18:0] Wgt_4_414,
input [18:0] Wgt_4_415,
input [18:0] Wgt_4_416,
input [18:0] Wgt_4_417,
input [18:0] Wgt_4_418,
input [18:0] Wgt_4_419,
input [18:0] Wgt_4_420,
input [18:0] Wgt_4_421,
input [18:0] Wgt_4_422,
input [18:0] Wgt_4_423,
input [18:0] Wgt_4_424,
input [18:0] Wgt_4_425,
input [18:0] Wgt_4_426,
input [18:0] Wgt_4_427,
input [18:0] Wgt_4_428,
input [18:0] Wgt_4_429,
input [18:0] Wgt_4_430,
input [18:0] Wgt_4_431,
input [18:0] Wgt_4_432,
input [18:0] Wgt_4_433,
input [18:0] Wgt_4_434,
input [18:0] Wgt_4_435,
input [18:0] Wgt_4_436,
input [18:0] Wgt_4_437,
input [18:0] Wgt_4_438,
input [18:0] Wgt_4_439,
input [18:0] Wgt_4_440,
input [18:0] Wgt_4_441,
input [18:0] Wgt_4_442,
input [18:0] Wgt_4_443,
input [18:0] Wgt_4_444,
input [18:0] Wgt_4_445,
input [18:0] Wgt_4_446,
input [18:0] Wgt_4_447,
input [18:0] Wgt_4_448,
input [18:0] Wgt_4_449,
input [18:0] Wgt_4_450,
input [18:0] Wgt_4_451,
input [18:0] Wgt_4_452,
input [18:0] Wgt_4_453,
input [18:0] Wgt_4_454,
input [18:0] Wgt_4_455,
input [18:0] Wgt_4_456,
input [18:0] Wgt_4_457,
input [18:0] Wgt_4_458,
input [18:0] Wgt_4_459,
input [18:0] Wgt_4_460,
input [18:0] Wgt_4_461,
input [18:0] Wgt_4_462,
input [18:0] Wgt_4_463,
input [18:0] Wgt_4_464,
input [18:0] Wgt_4_465,
input [18:0] Wgt_4_466,
input [18:0] Wgt_4_467,
input [18:0] Wgt_4_468,
input [18:0] Wgt_4_469,
input [18:0] Wgt_4_470,
input [18:0] Wgt_4_471,
input [18:0] Wgt_4_472,
input [18:0] Wgt_4_473,
input [18:0] Wgt_4_474,
input [18:0] Wgt_4_475,
input [18:0] Wgt_4_476,
input [18:0] Wgt_4_477,
input [18:0] Wgt_4_478,
input [18:0] Wgt_4_479,
input [18:0] Wgt_4_480,
input [18:0] Wgt_4_481,
input [18:0] Wgt_4_482,
input [18:0] Wgt_4_483,
input [18:0] Wgt_4_484,
input [18:0] Wgt_4_485,
input [18:0] Wgt_4_486,
input [18:0] Wgt_4_487,
input [18:0] Wgt_4_488,
input [18:0] Wgt_4_489,
input [18:0] Wgt_4_490,
input [18:0] Wgt_4_491,
input [18:0] Wgt_4_492,
input [18:0] Wgt_4_493,
input [18:0] Wgt_4_494,
input [18:0] Wgt_4_495,
input [18:0] Wgt_4_496,
input [18:0] Wgt_4_497,
input [18:0] Wgt_4_498,
input [18:0] Wgt_4_499,
input [18:0] Wgt_4_500,
input [18:0] Wgt_4_501,
input [18:0] Wgt_4_502,
input [18:0] Wgt_4_503,
input [18:0] Wgt_4_504,
input [18:0] Wgt_4_505,
input [18:0] Wgt_4_506,
input [18:0] Wgt_4_507,
input [18:0] Wgt_4_508,
input [18:0] Wgt_4_509,
input [18:0] Wgt_4_510,
input [18:0] Wgt_4_511,
input [18:0] Wgt_4_512,
input [18:0] Wgt_4_513,
input [18:0] Wgt_4_514,
input [18:0] Wgt_4_515,
input [18:0] Wgt_4_516,
input [18:0] Wgt_4_517,
input [18:0] Wgt_4_518,
input [18:0] Wgt_4_519,
input [18:0] Wgt_4_520,
input [18:0] Wgt_4_521,
input [18:0] Wgt_4_522,
input [18:0] Wgt_4_523,
input [18:0] Wgt_4_524,
input [18:0] Wgt_4_525,
input [18:0] Wgt_4_526,
input [18:0] Wgt_4_527,
input [18:0] Wgt_4_528,
input [18:0] Wgt_4_529,
input [18:0] Wgt_4_530,
input [18:0] Wgt_4_531,
input [18:0] Wgt_4_532,
input [18:0] Wgt_4_533,
input [18:0] Wgt_4_534,
input [18:0] Wgt_4_535,
input [18:0] Wgt_4_536,
input [18:0] Wgt_4_537,
input [18:0] Wgt_4_538,
input [18:0] Wgt_4_539,
input [18:0] Wgt_4_540,
input [18:0] Wgt_4_541,
input [18:0] Wgt_4_542,
input [18:0] Wgt_4_543,
input [18:0] Wgt_4_544,
input [18:0] Wgt_4_545,
input [18:0] Wgt_4_546,
input [18:0] Wgt_4_547,
input [18:0] Wgt_4_548,
input [18:0] Wgt_4_549,
input [18:0] Wgt_4_550,
input [18:0] Wgt_4_551,
input [18:0] Wgt_4_552,
input [18:0] Wgt_4_553,
input [18:0] Wgt_4_554,
input [18:0] Wgt_4_555,
input [18:0] Wgt_4_556,
input [18:0] Wgt_4_557,
input [18:0] Wgt_4_558,
input [18:0] Wgt_4_559,
input [18:0] Wgt_4_560,
input [18:0] Wgt_4_561,
input [18:0] Wgt_4_562,
input [18:0] Wgt_4_563,
input [18:0] Wgt_4_564,
input [18:0] Wgt_4_565,
input [18:0] Wgt_4_566,
input [18:0] Wgt_4_567,
input [18:0] Wgt_4_568,
input [18:0] Wgt_4_569,
input [18:0] Wgt_4_570,
input [18:0] Wgt_4_571,
input [18:0] Wgt_4_572,
input [18:0] Wgt_4_573,
input [18:0] Wgt_4_574,
input [18:0] Wgt_4_575,
input [18:0] Wgt_4_576,
input [18:0] Wgt_4_577,
input [18:0] Wgt_4_578,
input [18:0] Wgt_4_579,
input [18:0] Wgt_4_580,
input [18:0] Wgt_4_581,
input [18:0] Wgt_4_582,
input [18:0] Wgt_4_583,
input [18:0] Wgt_4_584,
input [18:0] Wgt_4_585,
input [18:0] Wgt_4_586,
input [18:0] Wgt_4_587,
input [18:0] Wgt_4_588,
input [18:0] Wgt_4_589,
input [18:0] Wgt_4_590,
input [18:0] Wgt_4_591,
input [18:0] Wgt_4_592,
input [18:0] Wgt_4_593,
input [18:0] Wgt_4_594,
input [18:0] Wgt_4_595,
input [18:0] Wgt_4_596,
input [18:0] Wgt_4_597,
input [18:0] Wgt_4_598,
input [18:0] Wgt_4_599,
input [18:0] Wgt_4_600,
input [18:0] Wgt_4_601,
input [18:0] Wgt_4_602,
input [18:0] Wgt_4_603,
input [18:0] Wgt_4_604,
input [18:0] Wgt_4_605,
input [18:0] Wgt_4_606,
input [18:0] Wgt_4_607,
input [18:0] Wgt_4_608,
input [18:0] Wgt_4_609,
input [18:0] Wgt_4_610,
input [18:0] Wgt_4_611,
input [18:0] Wgt_4_612,
input [18:0] Wgt_4_613,
input [18:0] Wgt_4_614,
input [18:0] Wgt_4_615,
input [18:0] Wgt_4_616,
input [18:0] Wgt_4_617,
input [18:0] Wgt_4_618,
input [18:0] Wgt_4_619,
input [18:0] Wgt_4_620,
input [18:0] Wgt_4_621,
input [18:0] Wgt_4_622,
input [18:0] Wgt_4_623,
input [18:0] Wgt_4_624,
input [18:0] Wgt_4_625,
input [18:0] Wgt_4_626,
input [18:0] Wgt_4_627,
input [18:0] Wgt_4_628,
input [18:0] Wgt_4_629,
input [18:0] Wgt_4_630,
input [18:0] Wgt_4_631,
input [18:0] Wgt_4_632,
input [18:0] Wgt_4_633,
input [18:0] Wgt_4_634,
input [18:0] Wgt_4_635,
input [18:0] Wgt_4_636,
input [18:0] Wgt_4_637,
input [18:0] Wgt_4_638,
input [18:0] Wgt_4_639,
input [18:0] Wgt_4_640,
input [18:0] Wgt_4_641,
input [18:0] Wgt_4_642,
input [18:0] Wgt_4_643,
input [18:0] Wgt_4_644,
input [18:0] Wgt_4_645,
input [18:0] Wgt_4_646,
input [18:0] Wgt_4_647,
input [18:0] Wgt_4_648,
input [18:0] Wgt_4_649,
input [18:0] Wgt_4_650,
input [18:0] Wgt_4_651,
input [18:0] Wgt_4_652,
input [18:0] Wgt_4_653,
input [18:0] Wgt_4_654,
input [18:0] Wgt_4_655,
input [18:0] Wgt_4_656,
input [18:0] Wgt_4_657,
input [18:0] Wgt_4_658,
input [18:0] Wgt_4_659,
input [18:0] Wgt_4_660,
input [18:0] Wgt_4_661,
input [18:0] Wgt_4_662,
input [18:0] Wgt_4_663,
input [18:0] Wgt_4_664,
input [18:0] Wgt_4_665,
input [18:0] Wgt_4_666,
input [18:0] Wgt_4_667,
input [18:0] Wgt_4_668,
input [18:0] Wgt_4_669,
input [18:0] Wgt_4_670,
input [18:0] Wgt_4_671,
input [18:0] Wgt_4_672,
input [18:0] Wgt_4_673,
input [18:0] Wgt_4_674,
input [18:0] Wgt_4_675,
input [18:0] Wgt_4_676,
input [18:0] Wgt_4_677,
input [18:0] Wgt_4_678,
input [18:0] Wgt_4_679,
input [18:0] Wgt_4_680,
input [18:0] Wgt_4_681,
input [18:0] Wgt_4_682,
input [18:0] Wgt_4_683,
input [18:0] Wgt_4_684,
input [18:0] Wgt_4_685,
input [18:0] Wgt_4_686,
input [18:0] Wgt_4_687,
input [18:0] Wgt_4_688,
input [18:0] Wgt_4_689,
input [18:0] Wgt_4_690,
input [18:0] Wgt_4_691,
input [18:0] Wgt_4_692,
input [18:0] Wgt_4_693,
input [18:0] Wgt_4_694,
input [18:0] Wgt_4_695,
input [18:0] Wgt_4_696,
input [18:0] Wgt_4_697,
input [18:0] Wgt_4_698,
input [18:0] Wgt_4_699,
input [18:0] Wgt_4_700,
input [18:0] Wgt_4_701,
input [18:0] Wgt_4_702,
input [18:0] Wgt_4_703,
input [18:0] Wgt_4_704,
input [18:0] Wgt_4_705,
input [18:0] Wgt_4_706,
input [18:0] Wgt_4_707,
input [18:0] Wgt_4_708,
input [18:0] Wgt_4_709,
input [18:0] Wgt_4_710,
input [18:0] Wgt_4_711,
input [18:0] Wgt_4_712,
input [18:0] Wgt_4_713,
input [18:0] Wgt_4_714,
input [18:0] Wgt_4_715,
input [18:0] Wgt_4_716,
input [18:0] Wgt_4_717,
input [18:0] Wgt_4_718,
input [18:0] Wgt_4_719,
input [18:0] Wgt_4_720,
input [18:0] Wgt_4_721,
input [18:0] Wgt_4_722,
input [18:0] Wgt_4_723,
input [18:0] Wgt_4_724,
input [18:0] Wgt_4_725,
input [18:0] Wgt_4_726,
input [18:0] Wgt_4_727,
input [18:0] Wgt_4_728,
input [18:0] Wgt_4_729,
input [18:0] Wgt_4_730,
input [18:0] Wgt_4_731,
input [18:0] Wgt_4_732,
input [18:0] Wgt_4_733,
input [18:0] Wgt_4_734,
input [18:0] Wgt_4_735,
input [18:0] Wgt_4_736,
input [18:0] Wgt_4_737,
input [18:0] Wgt_4_738,
input [18:0] Wgt_4_739,
input [18:0] Wgt_4_740,
input [18:0] Wgt_4_741,
input [18:0] Wgt_4_742,
input [18:0] Wgt_4_743,
input [18:0] Wgt_4_744,
input [18:0] Wgt_4_745,
input [18:0] Wgt_4_746,
input [18:0] Wgt_4_747,
input [18:0] Wgt_4_748,
input [18:0] Wgt_4_749,
input [18:0] Wgt_4_750,
input [18:0] Wgt_4_751,
input [18:0] Wgt_4_752,
input [18:0] Wgt_4_753,
input [18:0] Wgt_4_754,
input [18:0] Wgt_4_755,
input [18:0] Wgt_4_756,
input [18:0] Wgt_4_757,
input [18:0] Wgt_4_758,
input [18:0] Wgt_4_759,
input [18:0] Wgt_4_760,
input [18:0] Wgt_4_761,
input [18:0] Wgt_4_762,
input [18:0] Wgt_4_763,
input [18:0] Wgt_4_764,
input [18:0] Wgt_4_765,
input [18:0] Wgt_4_766,
input [18:0] Wgt_4_767,
input [18:0] Wgt_4_768,
input [18:0] Wgt_4_769,
input [18:0] Wgt_4_770,
input [18:0] Wgt_4_771,
input [18:0] Wgt_4_772,
input [18:0] Wgt_4_773,
input [18:0] Wgt_4_774,
input [18:0] Wgt_4_775,
input [18:0] Wgt_4_776,
input [18:0] Wgt_4_777,
input [18:0] Wgt_4_778,
input [18:0] Wgt_4_779,
input [18:0] Wgt_4_780,
input [18:0] Wgt_4_781,
input [18:0] Wgt_4_782,
input [18:0] Wgt_4_783,
input [18:0] Wgt_4_784,
input [18:0] Wgt_5_0,
input [18:0] Wgt_5_1,
input [18:0] Wgt_5_2,
input [18:0] Wgt_5_3,
input [18:0] Wgt_5_4,
input [18:0] Wgt_5_5,
input [18:0] Wgt_5_6,
input [18:0] Wgt_5_7,
input [18:0] Wgt_5_8,
input [18:0] Wgt_5_9,
input [18:0] Wgt_5_10,
input [18:0] Wgt_5_11,
input [18:0] Wgt_5_12,
input [18:0] Wgt_5_13,
input [18:0] Wgt_5_14,
input [18:0] Wgt_5_15,
input [18:0] Wgt_5_16,
input [18:0] Wgt_5_17,
input [18:0] Wgt_5_18,
input [18:0] Wgt_5_19,
input [18:0] Wgt_5_20,
input [18:0] Wgt_5_21,
input [18:0] Wgt_5_22,
input [18:0] Wgt_5_23,
input [18:0] Wgt_5_24,
input [18:0] Wgt_5_25,
input [18:0] Wgt_5_26,
input [18:0] Wgt_5_27,
input [18:0] Wgt_5_28,
input [18:0] Wgt_5_29,
input [18:0] Wgt_5_30,
input [18:0] Wgt_5_31,
input [18:0] Wgt_5_32,
input [18:0] Wgt_5_33,
input [18:0] Wgt_5_34,
input [18:0] Wgt_5_35,
input [18:0] Wgt_5_36,
input [18:0] Wgt_5_37,
input [18:0] Wgt_5_38,
input [18:0] Wgt_5_39,
input [18:0] Wgt_5_40,
input [18:0] Wgt_5_41,
input [18:0] Wgt_5_42,
input [18:0] Wgt_5_43,
input [18:0] Wgt_5_44,
input [18:0] Wgt_5_45,
input [18:0] Wgt_5_46,
input [18:0] Wgt_5_47,
input [18:0] Wgt_5_48,
input [18:0] Wgt_5_49,
input [18:0] Wgt_5_50,
input [18:0] Wgt_5_51,
input [18:0] Wgt_5_52,
input [18:0] Wgt_5_53,
input [18:0] Wgt_5_54,
input [18:0] Wgt_5_55,
input [18:0] Wgt_5_56,
input [18:0] Wgt_5_57,
input [18:0] Wgt_5_58,
input [18:0] Wgt_5_59,
input [18:0] Wgt_5_60,
input [18:0] Wgt_5_61,
input [18:0] Wgt_5_62,
input [18:0] Wgt_5_63,
input [18:0] Wgt_5_64,
input [18:0] Wgt_5_65,
input [18:0] Wgt_5_66,
input [18:0] Wgt_5_67,
input [18:0] Wgt_5_68,
input [18:0] Wgt_5_69,
input [18:0] Wgt_5_70,
input [18:0] Wgt_5_71,
input [18:0] Wgt_5_72,
input [18:0] Wgt_5_73,
input [18:0] Wgt_5_74,
input [18:0] Wgt_5_75,
input [18:0] Wgt_5_76,
input [18:0] Wgt_5_77,
input [18:0] Wgt_5_78,
input [18:0] Wgt_5_79,
input [18:0] Wgt_5_80,
input [18:0] Wgt_5_81,
input [18:0] Wgt_5_82,
input [18:0] Wgt_5_83,
input [18:0] Wgt_5_84,
input [18:0] Wgt_5_85,
input [18:0] Wgt_5_86,
input [18:0] Wgt_5_87,
input [18:0] Wgt_5_88,
input [18:0] Wgt_5_89,
input [18:0] Wgt_5_90,
input [18:0] Wgt_5_91,
input [18:0] Wgt_5_92,
input [18:0] Wgt_5_93,
input [18:0] Wgt_5_94,
input [18:0] Wgt_5_95,
input [18:0] Wgt_5_96,
input [18:0] Wgt_5_97,
input [18:0] Wgt_5_98,
input [18:0] Wgt_5_99,
input [18:0] Wgt_5_100,
input [18:0] Wgt_5_101,
input [18:0] Wgt_5_102,
input [18:0] Wgt_5_103,
input [18:0] Wgt_5_104,
input [18:0] Wgt_5_105,
input [18:0] Wgt_5_106,
input [18:0] Wgt_5_107,
input [18:0] Wgt_5_108,
input [18:0] Wgt_5_109,
input [18:0] Wgt_5_110,
input [18:0] Wgt_5_111,
input [18:0] Wgt_5_112,
input [18:0] Wgt_5_113,
input [18:0] Wgt_5_114,
input [18:0] Wgt_5_115,
input [18:0] Wgt_5_116,
input [18:0] Wgt_5_117,
input [18:0] Wgt_5_118,
input [18:0] Wgt_5_119,
input [18:0] Wgt_5_120,
input [18:0] Wgt_5_121,
input [18:0] Wgt_5_122,
input [18:0] Wgt_5_123,
input [18:0] Wgt_5_124,
input [18:0] Wgt_5_125,
input [18:0] Wgt_5_126,
input [18:0] Wgt_5_127,
input [18:0] Wgt_5_128,
input [18:0] Wgt_5_129,
input [18:0] Wgt_5_130,
input [18:0] Wgt_5_131,
input [18:0] Wgt_5_132,
input [18:0] Wgt_5_133,
input [18:0] Wgt_5_134,
input [18:0] Wgt_5_135,
input [18:0] Wgt_5_136,
input [18:0] Wgt_5_137,
input [18:0] Wgt_5_138,
input [18:0] Wgt_5_139,
input [18:0] Wgt_5_140,
input [18:0] Wgt_5_141,
input [18:0] Wgt_5_142,
input [18:0] Wgt_5_143,
input [18:0] Wgt_5_144,
input [18:0] Wgt_5_145,
input [18:0] Wgt_5_146,
input [18:0] Wgt_5_147,
input [18:0] Wgt_5_148,
input [18:0] Wgt_5_149,
input [18:0] Wgt_5_150,
input [18:0] Wgt_5_151,
input [18:0] Wgt_5_152,
input [18:0] Wgt_5_153,
input [18:0] Wgt_5_154,
input [18:0] Wgt_5_155,
input [18:0] Wgt_5_156,
input [18:0] Wgt_5_157,
input [18:0] Wgt_5_158,
input [18:0] Wgt_5_159,
input [18:0] Wgt_5_160,
input [18:0] Wgt_5_161,
input [18:0] Wgt_5_162,
input [18:0] Wgt_5_163,
input [18:0] Wgt_5_164,
input [18:0] Wgt_5_165,
input [18:0] Wgt_5_166,
input [18:0] Wgt_5_167,
input [18:0] Wgt_5_168,
input [18:0] Wgt_5_169,
input [18:0] Wgt_5_170,
input [18:0] Wgt_5_171,
input [18:0] Wgt_5_172,
input [18:0] Wgt_5_173,
input [18:0] Wgt_5_174,
input [18:0] Wgt_5_175,
input [18:0] Wgt_5_176,
input [18:0] Wgt_5_177,
input [18:0] Wgt_5_178,
input [18:0] Wgt_5_179,
input [18:0] Wgt_5_180,
input [18:0] Wgt_5_181,
input [18:0] Wgt_5_182,
input [18:0] Wgt_5_183,
input [18:0] Wgt_5_184,
input [18:0] Wgt_5_185,
input [18:0] Wgt_5_186,
input [18:0] Wgt_5_187,
input [18:0] Wgt_5_188,
input [18:0] Wgt_5_189,
input [18:0] Wgt_5_190,
input [18:0] Wgt_5_191,
input [18:0] Wgt_5_192,
input [18:0] Wgt_5_193,
input [18:0] Wgt_5_194,
input [18:0] Wgt_5_195,
input [18:0] Wgt_5_196,
input [18:0] Wgt_5_197,
input [18:0] Wgt_5_198,
input [18:0] Wgt_5_199,
input [18:0] Wgt_5_200,
input [18:0] Wgt_5_201,
input [18:0] Wgt_5_202,
input [18:0] Wgt_5_203,
input [18:0] Wgt_5_204,
input [18:0] Wgt_5_205,
input [18:0] Wgt_5_206,
input [18:0] Wgt_5_207,
input [18:0] Wgt_5_208,
input [18:0] Wgt_5_209,
input [18:0] Wgt_5_210,
input [18:0] Wgt_5_211,
input [18:0] Wgt_5_212,
input [18:0] Wgt_5_213,
input [18:0] Wgt_5_214,
input [18:0] Wgt_5_215,
input [18:0] Wgt_5_216,
input [18:0] Wgt_5_217,
input [18:0] Wgt_5_218,
input [18:0] Wgt_5_219,
input [18:0] Wgt_5_220,
input [18:0] Wgt_5_221,
input [18:0] Wgt_5_222,
input [18:0] Wgt_5_223,
input [18:0] Wgt_5_224,
input [18:0] Wgt_5_225,
input [18:0] Wgt_5_226,
input [18:0] Wgt_5_227,
input [18:0] Wgt_5_228,
input [18:0] Wgt_5_229,
input [18:0] Wgt_5_230,
input [18:0] Wgt_5_231,
input [18:0] Wgt_5_232,
input [18:0] Wgt_5_233,
input [18:0] Wgt_5_234,
input [18:0] Wgt_5_235,
input [18:0] Wgt_5_236,
input [18:0] Wgt_5_237,
input [18:0] Wgt_5_238,
input [18:0] Wgt_5_239,
input [18:0] Wgt_5_240,
input [18:0] Wgt_5_241,
input [18:0] Wgt_5_242,
input [18:0] Wgt_5_243,
input [18:0] Wgt_5_244,
input [18:0] Wgt_5_245,
input [18:0] Wgt_5_246,
input [18:0] Wgt_5_247,
input [18:0] Wgt_5_248,
input [18:0] Wgt_5_249,
input [18:0] Wgt_5_250,
input [18:0] Wgt_5_251,
input [18:0] Wgt_5_252,
input [18:0] Wgt_5_253,
input [18:0] Wgt_5_254,
input [18:0] Wgt_5_255,
input [18:0] Wgt_5_256,
input [18:0] Wgt_5_257,
input [18:0] Wgt_5_258,
input [18:0] Wgt_5_259,
input [18:0] Wgt_5_260,
input [18:0] Wgt_5_261,
input [18:0] Wgt_5_262,
input [18:0] Wgt_5_263,
input [18:0] Wgt_5_264,
input [18:0] Wgt_5_265,
input [18:0] Wgt_5_266,
input [18:0] Wgt_5_267,
input [18:0] Wgt_5_268,
input [18:0] Wgt_5_269,
input [18:0] Wgt_5_270,
input [18:0] Wgt_5_271,
input [18:0] Wgt_5_272,
input [18:0] Wgt_5_273,
input [18:0] Wgt_5_274,
input [18:0] Wgt_5_275,
input [18:0] Wgt_5_276,
input [18:0] Wgt_5_277,
input [18:0] Wgt_5_278,
input [18:0] Wgt_5_279,
input [18:0] Wgt_5_280,
input [18:0] Wgt_5_281,
input [18:0] Wgt_5_282,
input [18:0] Wgt_5_283,
input [18:0] Wgt_5_284,
input [18:0] Wgt_5_285,
input [18:0] Wgt_5_286,
input [18:0] Wgt_5_287,
input [18:0] Wgt_5_288,
input [18:0] Wgt_5_289,
input [18:0] Wgt_5_290,
input [18:0] Wgt_5_291,
input [18:0] Wgt_5_292,
input [18:0] Wgt_5_293,
input [18:0] Wgt_5_294,
input [18:0] Wgt_5_295,
input [18:0] Wgt_5_296,
input [18:0] Wgt_5_297,
input [18:0] Wgt_5_298,
input [18:0] Wgt_5_299,
input [18:0] Wgt_5_300,
input [18:0] Wgt_5_301,
input [18:0] Wgt_5_302,
input [18:0] Wgt_5_303,
input [18:0] Wgt_5_304,
input [18:0] Wgt_5_305,
input [18:0] Wgt_5_306,
input [18:0] Wgt_5_307,
input [18:0] Wgt_5_308,
input [18:0] Wgt_5_309,
input [18:0] Wgt_5_310,
input [18:0] Wgt_5_311,
input [18:0] Wgt_5_312,
input [18:0] Wgt_5_313,
input [18:0] Wgt_5_314,
input [18:0] Wgt_5_315,
input [18:0] Wgt_5_316,
input [18:0] Wgt_5_317,
input [18:0] Wgt_5_318,
input [18:0] Wgt_5_319,
input [18:0] Wgt_5_320,
input [18:0] Wgt_5_321,
input [18:0] Wgt_5_322,
input [18:0] Wgt_5_323,
input [18:0] Wgt_5_324,
input [18:0] Wgt_5_325,
input [18:0] Wgt_5_326,
input [18:0] Wgt_5_327,
input [18:0] Wgt_5_328,
input [18:0] Wgt_5_329,
input [18:0] Wgt_5_330,
input [18:0] Wgt_5_331,
input [18:0] Wgt_5_332,
input [18:0] Wgt_5_333,
input [18:0] Wgt_5_334,
input [18:0] Wgt_5_335,
input [18:0] Wgt_5_336,
input [18:0] Wgt_5_337,
input [18:0] Wgt_5_338,
input [18:0] Wgt_5_339,
input [18:0] Wgt_5_340,
input [18:0] Wgt_5_341,
input [18:0] Wgt_5_342,
input [18:0] Wgt_5_343,
input [18:0] Wgt_5_344,
input [18:0] Wgt_5_345,
input [18:0] Wgt_5_346,
input [18:0] Wgt_5_347,
input [18:0] Wgt_5_348,
input [18:0] Wgt_5_349,
input [18:0] Wgt_5_350,
input [18:0] Wgt_5_351,
input [18:0] Wgt_5_352,
input [18:0] Wgt_5_353,
input [18:0] Wgt_5_354,
input [18:0] Wgt_5_355,
input [18:0] Wgt_5_356,
input [18:0] Wgt_5_357,
input [18:0] Wgt_5_358,
input [18:0] Wgt_5_359,
input [18:0] Wgt_5_360,
input [18:0] Wgt_5_361,
input [18:0] Wgt_5_362,
input [18:0] Wgt_5_363,
input [18:0] Wgt_5_364,
input [18:0] Wgt_5_365,
input [18:0] Wgt_5_366,
input [18:0] Wgt_5_367,
input [18:0] Wgt_5_368,
input [18:0] Wgt_5_369,
input [18:0] Wgt_5_370,
input [18:0] Wgt_5_371,
input [18:0] Wgt_5_372,
input [18:0] Wgt_5_373,
input [18:0] Wgt_5_374,
input [18:0] Wgt_5_375,
input [18:0] Wgt_5_376,
input [18:0] Wgt_5_377,
input [18:0] Wgt_5_378,
input [18:0] Wgt_5_379,
input [18:0] Wgt_5_380,
input [18:0] Wgt_5_381,
input [18:0] Wgt_5_382,
input [18:0] Wgt_5_383,
input [18:0] Wgt_5_384,
input [18:0] Wgt_5_385,
input [18:0] Wgt_5_386,
input [18:0] Wgt_5_387,
input [18:0] Wgt_5_388,
input [18:0] Wgt_5_389,
input [18:0] Wgt_5_390,
input [18:0] Wgt_5_391,
input [18:0] Wgt_5_392,
input [18:0] Wgt_5_393,
input [18:0] Wgt_5_394,
input [18:0] Wgt_5_395,
input [18:0] Wgt_5_396,
input [18:0] Wgt_5_397,
input [18:0] Wgt_5_398,
input [18:0] Wgt_5_399,
input [18:0] Wgt_5_400,
input [18:0] Wgt_5_401,
input [18:0] Wgt_5_402,
input [18:0] Wgt_5_403,
input [18:0] Wgt_5_404,
input [18:0] Wgt_5_405,
input [18:0] Wgt_5_406,
input [18:0] Wgt_5_407,
input [18:0] Wgt_5_408,
input [18:0] Wgt_5_409,
input [18:0] Wgt_5_410,
input [18:0] Wgt_5_411,
input [18:0] Wgt_5_412,
input [18:0] Wgt_5_413,
input [18:0] Wgt_5_414,
input [18:0] Wgt_5_415,
input [18:0] Wgt_5_416,
input [18:0] Wgt_5_417,
input [18:0] Wgt_5_418,
input [18:0] Wgt_5_419,
input [18:0] Wgt_5_420,
input [18:0] Wgt_5_421,
input [18:0] Wgt_5_422,
input [18:0] Wgt_5_423,
input [18:0] Wgt_5_424,
input [18:0] Wgt_5_425,
input [18:0] Wgt_5_426,
input [18:0] Wgt_5_427,
input [18:0] Wgt_5_428,
input [18:0] Wgt_5_429,
input [18:0] Wgt_5_430,
input [18:0] Wgt_5_431,
input [18:0] Wgt_5_432,
input [18:0] Wgt_5_433,
input [18:0] Wgt_5_434,
input [18:0] Wgt_5_435,
input [18:0] Wgt_5_436,
input [18:0] Wgt_5_437,
input [18:0] Wgt_5_438,
input [18:0] Wgt_5_439,
input [18:0] Wgt_5_440,
input [18:0] Wgt_5_441,
input [18:0] Wgt_5_442,
input [18:0] Wgt_5_443,
input [18:0] Wgt_5_444,
input [18:0] Wgt_5_445,
input [18:0] Wgt_5_446,
input [18:0] Wgt_5_447,
input [18:0] Wgt_5_448,
input [18:0] Wgt_5_449,
input [18:0] Wgt_5_450,
input [18:0] Wgt_5_451,
input [18:0] Wgt_5_452,
input [18:0] Wgt_5_453,
input [18:0] Wgt_5_454,
input [18:0] Wgt_5_455,
input [18:0] Wgt_5_456,
input [18:0] Wgt_5_457,
input [18:0] Wgt_5_458,
input [18:0] Wgt_5_459,
input [18:0] Wgt_5_460,
input [18:0] Wgt_5_461,
input [18:0] Wgt_5_462,
input [18:0] Wgt_5_463,
input [18:0] Wgt_5_464,
input [18:0] Wgt_5_465,
input [18:0] Wgt_5_466,
input [18:0] Wgt_5_467,
input [18:0] Wgt_5_468,
input [18:0] Wgt_5_469,
input [18:0] Wgt_5_470,
input [18:0] Wgt_5_471,
input [18:0] Wgt_5_472,
input [18:0] Wgt_5_473,
input [18:0] Wgt_5_474,
input [18:0] Wgt_5_475,
input [18:0] Wgt_5_476,
input [18:0] Wgt_5_477,
input [18:0] Wgt_5_478,
input [18:0] Wgt_5_479,
input [18:0] Wgt_5_480,
input [18:0] Wgt_5_481,
input [18:0] Wgt_5_482,
input [18:0] Wgt_5_483,
input [18:0] Wgt_5_484,
input [18:0] Wgt_5_485,
input [18:0] Wgt_5_486,
input [18:0] Wgt_5_487,
input [18:0] Wgt_5_488,
input [18:0] Wgt_5_489,
input [18:0] Wgt_5_490,
input [18:0] Wgt_5_491,
input [18:0] Wgt_5_492,
input [18:0] Wgt_5_493,
input [18:0] Wgt_5_494,
input [18:0] Wgt_5_495,
input [18:0] Wgt_5_496,
input [18:0] Wgt_5_497,
input [18:0] Wgt_5_498,
input [18:0] Wgt_5_499,
input [18:0] Wgt_5_500,
input [18:0] Wgt_5_501,
input [18:0] Wgt_5_502,
input [18:0] Wgt_5_503,
input [18:0] Wgt_5_504,
input [18:0] Wgt_5_505,
input [18:0] Wgt_5_506,
input [18:0] Wgt_5_507,
input [18:0] Wgt_5_508,
input [18:0] Wgt_5_509,
input [18:0] Wgt_5_510,
input [18:0] Wgt_5_511,
input [18:0] Wgt_5_512,
input [18:0] Wgt_5_513,
input [18:0] Wgt_5_514,
input [18:0] Wgt_5_515,
input [18:0] Wgt_5_516,
input [18:0] Wgt_5_517,
input [18:0] Wgt_5_518,
input [18:0] Wgt_5_519,
input [18:0] Wgt_5_520,
input [18:0] Wgt_5_521,
input [18:0] Wgt_5_522,
input [18:0] Wgt_5_523,
input [18:0] Wgt_5_524,
input [18:0] Wgt_5_525,
input [18:0] Wgt_5_526,
input [18:0] Wgt_5_527,
input [18:0] Wgt_5_528,
input [18:0] Wgt_5_529,
input [18:0] Wgt_5_530,
input [18:0] Wgt_5_531,
input [18:0] Wgt_5_532,
input [18:0] Wgt_5_533,
input [18:0] Wgt_5_534,
input [18:0] Wgt_5_535,
input [18:0] Wgt_5_536,
input [18:0] Wgt_5_537,
input [18:0] Wgt_5_538,
input [18:0] Wgt_5_539,
input [18:0] Wgt_5_540,
input [18:0] Wgt_5_541,
input [18:0] Wgt_5_542,
input [18:0] Wgt_5_543,
input [18:0] Wgt_5_544,
input [18:0] Wgt_5_545,
input [18:0] Wgt_5_546,
input [18:0] Wgt_5_547,
input [18:0] Wgt_5_548,
input [18:0] Wgt_5_549,
input [18:0] Wgt_5_550,
input [18:0] Wgt_5_551,
input [18:0] Wgt_5_552,
input [18:0] Wgt_5_553,
input [18:0] Wgt_5_554,
input [18:0] Wgt_5_555,
input [18:0] Wgt_5_556,
input [18:0] Wgt_5_557,
input [18:0] Wgt_5_558,
input [18:0] Wgt_5_559,
input [18:0] Wgt_5_560,
input [18:0] Wgt_5_561,
input [18:0] Wgt_5_562,
input [18:0] Wgt_5_563,
input [18:0] Wgt_5_564,
input [18:0] Wgt_5_565,
input [18:0] Wgt_5_566,
input [18:0] Wgt_5_567,
input [18:0] Wgt_5_568,
input [18:0] Wgt_5_569,
input [18:0] Wgt_5_570,
input [18:0] Wgt_5_571,
input [18:0] Wgt_5_572,
input [18:0] Wgt_5_573,
input [18:0] Wgt_5_574,
input [18:0] Wgt_5_575,
input [18:0] Wgt_5_576,
input [18:0] Wgt_5_577,
input [18:0] Wgt_5_578,
input [18:0] Wgt_5_579,
input [18:0] Wgt_5_580,
input [18:0] Wgt_5_581,
input [18:0] Wgt_5_582,
input [18:0] Wgt_5_583,
input [18:0] Wgt_5_584,
input [18:0] Wgt_5_585,
input [18:0] Wgt_5_586,
input [18:0] Wgt_5_587,
input [18:0] Wgt_5_588,
input [18:0] Wgt_5_589,
input [18:0] Wgt_5_590,
input [18:0] Wgt_5_591,
input [18:0] Wgt_5_592,
input [18:0] Wgt_5_593,
input [18:0] Wgt_5_594,
input [18:0] Wgt_5_595,
input [18:0] Wgt_5_596,
input [18:0] Wgt_5_597,
input [18:0] Wgt_5_598,
input [18:0] Wgt_5_599,
input [18:0] Wgt_5_600,
input [18:0] Wgt_5_601,
input [18:0] Wgt_5_602,
input [18:0] Wgt_5_603,
input [18:0] Wgt_5_604,
input [18:0] Wgt_5_605,
input [18:0] Wgt_5_606,
input [18:0] Wgt_5_607,
input [18:0] Wgt_5_608,
input [18:0] Wgt_5_609,
input [18:0] Wgt_5_610,
input [18:0] Wgt_5_611,
input [18:0] Wgt_5_612,
input [18:0] Wgt_5_613,
input [18:0] Wgt_5_614,
input [18:0] Wgt_5_615,
input [18:0] Wgt_5_616,
input [18:0] Wgt_5_617,
input [18:0] Wgt_5_618,
input [18:0] Wgt_5_619,
input [18:0] Wgt_5_620,
input [18:0] Wgt_5_621,
input [18:0] Wgt_5_622,
input [18:0] Wgt_5_623,
input [18:0] Wgt_5_624,
input [18:0] Wgt_5_625,
input [18:0] Wgt_5_626,
input [18:0] Wgt_5_627,
input [18:0] Wgt_5_628,
input [18:0] Wgt_5_629,
input [18:0] Wgt_5_630,
input [18:0] Wgt_5_631,
input [18:0] Wgt_5_632,
input [18:0] Wgt_5_633,
input [18:0] Wgt_5_634,
input [18:0] Wgt_5_635,
input [18:0] Wgt_5_636,
input [18:0] Wgt_5_637,
input [18:0] Wgt_5_638,
input [18:0] Wgt_5_639,
input [18:0] Wgt_5_640,
input [18:0] Wgt_5_641,
input [18:0] Wgt_5_642,
input [18:0] Wgt_5_643,
input [18:0] Wgt_5_644,
input [18:0] Wgt_5_645,
input [18:0] Wgt_5_646,
input [18:0] Wgt_5_647,
input [18:0] Wgt_5_648,
input [18:0] Wgt_5_649,
input [18:0] Wgt_5_650,
input [18:0] Wgt_5_651,
input [18:0] Wgt_5_652,
input [18:0] Wgt_5_653,
input [18:0] Wgt_5_654,
input [18:0] Wgt_5_655,
input [18:0] Wgt_5_656,
input [18:0] Wgt_5_657,
input [18:0] Wgt_5_658,
input [18:0] Wgt_5_659,
input [18:0] Wgt_5_660,
input [18:0] Wgt_5_661,
input [18:0] Wgt_5_662,
input [18:0] Wgt_5_663,
input [18:0] Wgt_5_664,
input [18:0] Wgt_5_665,
input [18:0] Wgt_5_666,
input [18:0] Wgt_5_667,
input [18:0] Wgt_5_668,
input [18:0] Wgt_5_669,
input [18:0] Wgt_5_670,
input [18:0] Wgt_5_671,
input [18:0] Wgt_5_672,
input [18:0] Wgt_5_673,
input [18:0] Wgt_5_674,
input [18:0] Wgt_5_675,
input [18:0] Wgt_5_676,
input [18:0] Wgt_5_677,
input [18:0] Wgt_5_678,
input [18:0] Wgt_5_679,
input [18:0] Wgt_5_680,
input [18:0] Wgt_5_681,
input [18:0] Wgt_5_682,
input [18:0] Wgt_5_683,
input [18:0] Wgt_5_684,
input [18:0] Wgt_5_685,
input [18:0] Wgt_5_686,
input [18:0] Wgt_5_687,
input [18:0] Wgt_5_688,
input [18:0] Wgt_5_689,
input [18:0] Wgt_5_690,
input [18:0] Wgt_5_691,
input [18:0] Wgt_5_692,
input [18:0] Wgt_5_693,
input [18:0] Wgt_5_694,
input [18:0] Wgt_5_695,
input [18:0] Wgt_5_696,
input [18:0] Wgt_5_697,
input [18:0] Wgt_5_698,
input [18:0] Wgt_5_699,
input [18:0] Wgt_5_700,
input [18:0] Wgt_5_701,
input [18:0] Wgt_5_702,
input [18:0] Wgt_5_703,
input [18:0] Wgt_5_704,
input [18:0] Wgt_5_705,
input [18:0] Wgt_5_706,
input [18:0] Wgt_5_707,
input [18:0] Wgt_5_708,
input [18:0] Wgt_5_709,
input [18:0] Wgt_5_710,
input [18:0] Wgt_5_711,
input [18:0] Wgt_5_712,
input [18:0] Wgt_5_713,
input [18:0] Wgt_5_714,
input [18:0] Wgt_5_715,
input [18:0] Wgt_5_716,
input [18:0] Wgt_5_717,
input [18:0] Wgt_5_718,
input [18:0] Wgt_5_719,
input [18:0] Wgt_5_720,
input [18:0] Wgt_5_721,
input [18:0] Wgt_5_722,
input [18:0] Wgt_5_723,
input [18:0] Wgt_5_724,
input [18:0] Wgt_5_725,
input [18:0] Wgt_5_726,
input [18:0] Wgt_5_727,
input [18:0] Wgt_5_728,
input [18:0] Wgt_5_729,
input [18:0] Wgt_5_730,
input [18:0] Wgt_5_731,
input [18:0] Wgt_5_732,
input [18:0] Wgt_5_733,
input [18:0] Wgt_5_734,
input [18:0] Wgt_5_735,
input [18:0] Wgt_5_736,
input [18:0] Wgt_5_737,
input [18:0] Wgt_5_738,
input [18:0] Wgt_5_739,
input [18:0] Wgt_5_740,
input [18:0] Wgt_5_741,
input [18:0] Wgt_5_742,
input [18:0] Wgt_5_743,
input [18:0] Wgt_5_744,
input [18:0] Wgt_5_745,
input [18:0] Wgt_5_746,
input [18:0] Wgt_5_747,
input [18:0] Wgt_5_748,
input [18:0] Wgt_5_749,
input [18:0] Wgt_5_750,
input [18:0] Wgt_5_751,
input [18:0] Wgt_5_752,
input [18:0] Wgt_5_753,
input [18:0] Wgt_5_754,
input [18:0] Wgt_5_755,
input [18:0] Wgt_5_756,
input [18:0] Wgt_5_757,
input [18:0] Wgt_5_758,
input [18:0] Wgt_5_759,
input [18:0] Wgt_5_760,
input [18:0] Wgt_5_761,
input [18:0] Wgt_5_762,
input [18:0] Wgt_5_763,
input [18:0] Wgt_5_764,
input [18:0] Wgt_5_765,
input [18:0] Wgt_5_766,
input [18:0] Wgt_5_767,
input [18:0] Wgt_5_768,
input [18:0] Wgt_5_769,
input [18:0] Wgt_5_770,
input [18:0] Wgt_5_771,
input [18:0] Wgt_5_772,
input [18:0] Wgt_5_773,
input [18:0] Wgt_5_774,
input [18:0] Wgt_5_775,
input [18:0] Wgt_5_776,
input [18:0] Wgt_5_777,
input [18:0] Wgt_5_778,
input [18:0] Wgt_5_779,
input [18:0] Wgt_5_780,
input [18:0] Wgt_5_781,
input [18:0] Wgt_5_782,
input [18:0] Wgt_5_783,
input [18:0] Wgt_5_784,
input [18:0] Wgt_6_0,
input [18:0] Wgt_6_1,
input [18:0] Wgt_6_2,
input [18:0] Wgt_6_3,
input [18:0] Wgt_6_4,
input [18:0] Wgt_6_5,
input [18:0] Wgt_6_6,
input [18:0] Wgt_6_7,
input [18:0] Wgt_6_8,
input [18:0] Wgt_6_9,
input [18:0] Wgt_6_10,
input [18:0] Wgt_6_11,
input [18:0] Wgt_6_12,
input [18:0] Wgt_6_13,
input [18:0] Wgt_6_14,
input [18:0] Wgt_6_15,
input [18:0] Wgt_6_16,
input [18:0] Wgt_6_17,
input [18:0] Wgt_6_18,
input [18:0] Wgt_6_19,
input [18:0] Wgt_6_20,
input [18:0] Wgt_6_21,
input [18:0] Wgt_6_22,
input [18:0] Wgt_6_23,
input [18:0] Wgt_6_24,
input [18:0] Wgt_6_25,
input [18:0] Wgt_6_26,
input [18:0] Wgt_6_27,
input [18:0] Wgt_6_28,
input [18:0] Wgt_6_29,
input [18:0] Wgt_6_30,
input [18:0] Wgt_6_31,
input [18:0] Wgt_6_32,
input [18:0] Wgt_6_33,
input [18:0] Wgt_6_34,
input [18:0] Wgt_6_35,
input [18:0] Wgt_6_36,
input [18:0] Wgt_6_37,
input [18:0] Wgt_6_38,
input [18:0] Wgt_6_39,
input [18:0] Wgt_6_40,
input [18:0] Wgt_6_41,
input [18:0] Wgt_6_42,
input [18:0] Wgt_6_43,
input [18:0] Wgt_6_44,
input [18:0] Wgt_6_45,
input [18:0] Wgt_6_46,
input [18:0] Wgt_6_47,
input [18:0] Wgt_6_48,
input [18:0] Wgt_6_49,
input [18:0] Wgt_6_50,
input [18:0] Wgt_6_51,
input [18:0] Wgt_6_52,
input [18:0] Wgt_6_53,
input [18:0] Wgt_6_54,
input [18:0] Wgt_6_55,
input [18:0] Wgt_6_56,
input [18:0] Wgt_6_57,
input [18:0] Wgt_6_58,
input [18:0] Wgt_6_59,
input [18:0] Wgt_6_60,
input [18:0] Wgt_6_61,
input [18:0] Wgt_6_62,
input [18:0] Wgt_6_63,
input [18:0] Wgt_6_64,
input [18:0] Wgt_6_65,
input [18:0] Wgt_6_66,
input [18:0] Wgt_6_67,
input [18:0] Wgt_6_68,
input [18:0] Wgt_6_69,
input [18:0] Wgt_6_70,
input [18:0] Wgt_6_71,
input [18:0] Wgt_6_72,
input [18:0] Wgt_6_73,
input [18:0] Wgt_6_74,
input [18:0] Wgt_6_75,
input [18:0] Wgt_6_76,
input [18:0] Wgt_6_77,
input [18:0] Wgt_6_78,
input [18:0] Wgt_6_79,
input [18:0] Wgt_6_80,
input [18:0] Wgt_6_81,
input [18:0] Wgt_6_82,
input [18:0] Wgt_6_83,
input [18:0] Wgt_6_84,
input [18:0] Wgt_6_85,
input [18:0] Wgt_6_86,
input [18:0] Wgt_6_87,
input [18:0] Wgt_6_88,
input [18:0] Wgt_6_89,
input [18:0] Wgt_6_90,
input [18:0] Wgt_6_91,
input [18:0] Wgt_6_92,
input [18:0] Wgt_6_93,
input [18:0] Wgt_6_94,
input [18:0] Wgt_6_95,
input [18:0] Wgt_6_96,
input [18:0] Wgt_6_97,
input [18:0] Wgt_6_98,
input [18:0] Wgt_6_99,
input [18:0] Wgt_6_100,
input [18:0] Wgt_6_101,
input [18:0] Wgt_6_102,
input [18:0] Wgt_6_103,
input [18:0] Wgt_6_104,
input [18:0] Wgt_6_105,
input [18:0] Wgt_6_106,
input [18:0] Wgt_6_107,
input [18:0] Wgt_6_108,
input [18:0] Wgt_6_109,
input [18:0] Wgt_6_110,
input [18:0] Wgt_6_111,
input [18:0] Wgt_6_112,
input [18:0] Wgt_6_113,
input [18:0] Wgt_6_114,
input [18:0] Wgt_6_115,
input [18:0] Wgt_6_116,
input [18:0] Wgt_6_117,
input [18:0] Wgt_6_118,
input [18:0] Wgt_6_119,
input [18:0] Wgt_6_120,
input [18:0] Wgt_6_121,
input [18:0] Wgt_6_122,
input [18:0] Wgt_6_123,
input [18:0] Wgt_6_124,
input [18:0] Wgt_6_125,
input [18:0] Wgt_6_126,
input [18:0] Wgt_6_127,
input [18:0] Wgt_6_128,
input [18:0] Wgt_6_129,
input [18:0] Wgt_6_130,
input [18:0] Wgt_6_131,
input [18:0] Wgt_6_132,
input [18:0] Wgt_6_133,
input [18:0] Wgt_6_134,
input [18:0] Wgt_6_135,
input [18:0] Wgt_6_136,
input [18:0] Wgt_6_137,
input [18:0] Wgt_6_138,
input [18:0] Wgt_6_139,
input [18:0] Wgt_6_140,
input [18:0] Wgt_6_141,
input [18:0] Wgt_6_142,
input [18:0] Wgt_6_143,
input [18:0] Wgt_6_144,
input [18:0] Wgt_6_145,
input [18:0] Wgt_6_146,
input [18:0] Wgt_6_147,
input [18:0] Wgt_6_148,
input [18:0] Wgt_6_149,
input [18:0] Wgt_6_150,
input [18:0] Wgt_6_151,
input [18:0] Wgt_6_152,
input [18:0] Wgt_6_153,
input [18:0] Wgt_6_154,
input [18:0] Wgt_6_155,
input [18:0] Wgt_6_156,
input [18:0] Wgt_6_157,
input [18:0] Wgt_6_158,
input [18:0] Wgt_6_159,
input [18:0] Wgt_6_160,
input [18:0] Wgt_6_161,
input [18:0] Wgt_6_162,
input [18:0] Wgt_6_163,
input [18:0] Wgt_6_164,
input [18:0] Wgt_6_165,
input [18:0] Wgt_6_166,
input [18:0] Wgt_6_167,
input [18:0] Wgt_6_168,
input [18:0] Wgt_6_169,
input [18:0] Wgt_6_170,
input [18:0] Wgt_6_171,
input [18:0] Wgt_6_172,
input [18:0] Wgt_6_173,
input [18:0] Wgt_6_174,
input [18:0] Wgt_6_175,
input [18:0] Wgt_6_176,
input [18:0] Wgt_6_177,
input [18:0] Wgt_6_178,
input [18:0] Wgt_6_179,
input [18:0] Wgt_6_180,
input [18:0] Wgt_6_181,
input [18:0] Wgt_6_182,
input [18:0] Wgt_6_183,
input [18:0] Wgt_6_184,
input [18:0] Wgt_6_185,
input [18:0] Wgt_6_186,
input [18:0] Wgt_6_187,
input [18:0] Wgt_6_188,
input [18:0] Wgt_6_189,
input [18:0] Wgt_6_190,
input [18:0] Wgt_6_191,
input [18:0] Wgt_6_192,
input [18:0] Wgt_6_193,
input [18:0] Wgt_6_194,
input [18:0] Wgt_6_195,
input [18:0] Wgt_6_196,
input [18:0] Wgt_6_197,
input [18:0] Wgt_6_198,
input [18:0] Wgt_6_199,
input [18:0] Wgt_6_200,
input [18:0] Wgt_6_201,
input [18:0] Wgt_6_202,
input [18:0] Wgt_6_203,
input [18:0] Wgt_6_204,
input [18:0] Wgt_6_205,
input [18:0] Wgt_6_206,
input [18:0] Wgt_6_207,
input [18:0] Wgt_6_208,
input [18:0] Wgt_6_209,
input [18:0] Wgt_6_210,
input [18:0] Wgt_6_211,
input [18:0] Wgt_6_212,
input [18:0] Wgt_6_213,
input [18:0] Wgt_6_214,
input [18:0] Wgt_6_215,
input [18:0] Wgt_6_216,
input [18:0] Wgt_6_217,
input [18:0] Wgt_6_218,
input [18:0] Wgt_6_219,
input [18:0] Wgt_6_220,
input [18:0] Wgt_6_221,
input [18:0] Wgt_6_222,
input [18:0] Wgt_6_223,
input [18:0] Wgt_6_224,
input [18:0] Wgt_6_225,
input [18:0] Wgt_6_226,
input [18:0] Wgt_6_227,
input [18:0] Wgt_6_228,
input [18:0] Wgt_6_229,
input [18:0] Wgt_6_230,
input [18:0] Wgt_6_231,
input [18:0] Wgt_6_232,
input [18:0] Wgt_6_233,
input [18:0] Wgt_6_234,
input [18:0] Wgt_6_235,
input [18:0] Wgt_6_236,
input [18:0] Wgt_6_237,
input [18:0] Wgt_6_238,
input [18:0] Wgt_6_239,
input [18:0] Wgt_6_240,
input [18:0] Wgt_6_241,
input [18:0] Wgt_6_242,
input [18:0] Wgt_6_243,
input [18:0] Wgt_6_244,
input [18:0] Wgt_6_245,
input [18:0] Wgt_6_246,
input [18:0] Wgt_6_247,
input [18:0] Wgt_6_248,
input [18:0] Wgt_6_249,
input [18:0] Wgt_6_250,
input [18:0] Wgt_6_251,
input [18:0] Wgt_6_252,
input [18:0] Wgt_6_253,
input [18:0] Wgt_6_254,
input [18:0] Wgt_6_255,
input [18:0] Wgt_6_256,
input [18:0] Wgt_6_257,
input [18:0] Wgt_6_258,
input [18:0] Wgt_6_259,
input [18:0] Wgt_6_260,
input [18:0] Wgt_6_261,
input [18:0] Wgt_6_262,
input [18:0] Wgt_6_263,
input [18:0] Wgt_6_264,
input [18:0] Wgt_6_265,
input [18:0] Wgt_6_266,
input [18:0] Wgt_6_267,
input [18:0] Wgt_6_268,
input [18:0] Wgt_6_269,
input [18:0] Wgt_6_270,
input [18:0] Wgt_6_271,
input [18:0] Wgt_6_272,
input [18:0] Wgt_6_273,
input [18:0] Wgt_6_274,
input [18:0] Wgt_6_275,
input [18:0] Wgt_6_276,
input [18:0] Wgt_6_277,
input [18:0] Wgt_6_278,
input [18:0] Wgt_6_279,
input [18:0] Wgt_6_280,
input [18:0] Wgt_6_281,
input [18:0] Wgt_6_282,
input [18:0] Wgt_6_283,
input [18:0] Wgt_6_284,
input [18:0] Wgt_6_285,
input [18:0] Wgt_6_286,
input [18:0] Wgt_6_287,
input [18:0] Wgt_6_288,
input [18:0] Wgt_6_289,
input [18:0] Wgt_6_290,
input [18:0] Wgt_6_291,
input [18:0] Wgt_6_292,
input [18:0] Wgt_6_293,
input [18:0] Wgt_6_294,
input [18:0] Wgt_6_295,
input [18:0] Wgt_6_296,
input [18:0] Wgt_6_297,
input [18:0] Wgt_6_298,
input [18:0] Wgt_6_299,
input [18:0] Wgt_6_300,
input [18:0] Wgt_6_301,
input [18:0] Wgt_6_302,
input [18:0] Wgt_6_303,
input [18:0] Wgt_6_304,
input [18:0] Wgt_6_305,
input [18:0] Wgt_6_306,
input [18:0] Wgt_6_307,
input [18:0] Wgt_6_308,
input [18:0] Wgt_6_309,
input [18:0] Wgt_6_310,
input [18:0] Wgt_6_311,
input [18:0] Wgt_6_312,
input [18:0] Wgt_6_313,
input [18:0] Wgt_6_314,
input [18:0] Wgt_6_315,
input [18:0] Wgt_6_316,
input [18:0] Wgt_6_317,
input [18:0] Wgt_6_318,
input [18:0] Wgt_6_319,
input [18:0] Wgt_6_320,
input [18:0] Wgt_6_321,
input [18:0] Wgt_6_322,
input [18:0] Wgt_6_323,
input [18:0] Wgt_6_324,
input [18:0] Wgt_6_325,
input [18:0] Wgt_6_326,
input [18:0] Wgt_6_327,
input [18:0] Wgt_6_328,
input [18:0] Wgt_6_329,
input [18:0] Wgt_6_330,
input [18:0] Wgt_6_331,
input [18:0] Wgt_6_332,
input [18:0] Wgt_6_333,
input [18:0] Wgt_6_334,
input [18:0] Wgt_6_335,
input [18:0] Wgt_6_336,
input [18:0] Wgt_6_337,
input [18:0] Wgt_6_338,
input [18:0] Wgt_6_339,
input [18:0] Wgt_6_340,
input [18:0] Wgt_6_341,
input [18:0] Wgt_6_342,
input [18:0] Wgt_6_343,
input [18:0] Wgt_6_344,
input [18:0] Wgt_6_345,
input [18:0] Wgt_6_346,
input [18:0] Wgt_6_347,
input [18:0] Wgt_6_348,
input [18:0] Wgt_6_349,
input [18:0] Wgt_6_350,
input [18:0] Wgt_6_351,
input [18:0] Wgt_6_352,
input [18:0] Wgt_6_353,
input [18:0] Wgt_6_354,
input [18:0] Wgt_6_355,
input [18:0] Wgt_6_356,
input [18:0] Wgt_6_357,
input [18:0] Wgt_6_358,
input [18:0] Wgt_6_359,
input [18:0] Wgt_6_360,
input [18:0] Wgt_6_361,
input [18:0] Wgt_6_362,
input [18:0] Wgt_6_363,
input [18:0] Wgt_6_364,
input [18:0] Wgt_6_365,
input [18:0] Wgt_6_366,
input [18:0] Wgt_6_367,
input [18:0] Wgt_6_368,
input [18:0] Wgt_6_369,
input [18:0] Wgt_6_370,
input [18:0] Wgt_6_371,
input [18:0] Wgt_6_372,
input [18:0] Wgt_6_373,
input [18:0] Wgt_6_374,
input [18:0] Wgt_6_375,
input [18:0] Wgt_6_376,
input [18:0] Wgt_6_377,
input [18:0] Wgt_6_378,
input [18:0] Wgt_6_379,
input [18:0] Wgt_6_380,
input [18:0] Wgt_6_381,
input [18:0] Wgt_6_382,
input [18:0] Wgt_6_383,
input [18:0] Wgt_6_384,
input [18:0] Wgt_6_385,
input [18:0] Wgt_6_386,
input [18:0] Wgt_6_387,
input [18:0] Wgt_6_388,
input [18:0] Wgt_6_389,
input [18:0] Wgt_6_390,
input [18:0] Wgt_6_391,
input [18:0] Wgt_6_392,
input [18:0] Wgt_6_393,
input [18:0] Wgt_6_394,
input [18:0] Wgt_6_395,
input [18:0] Wgt_6_396,
input [18:0] Wgt_6_397,
input [18:0] Wgt_6_398,
input [18:0] Wgt_6_399,
input [18:0] Wgt_6_400,
input [18:0] Wgt_6_401,
input [18:0] Wgt_6_402,
input [18:0] Wgt_6_403,
input [18:0] Wgt_6_404,
input [18:0] Wgt_6_405,
input [18:0] Wgt_6_406,
input [18:0] Wgt_6_407,
input [18:0] Wgt_6_408,
input [18:0] Wgt_6_409,
input [18:0] Wgt_6_410,
input [18:0] Wgt_6_411,
input [18:0] Wgt_6_412,
input [18:0] Wgt_6_413,
input [18:0] Wgt_6_414,
input [18:0] Wgt_6_415,
input [18:0] Wgt_6_416,
input [18:0] Wgt_6_417,
input [18:0] Wgt_6_418,
input [18:0] Wgt_6_419,
input [18:0] Wgt_6_420,
input [18:0] Wgt_6_421,
input [18:0] Wgt_6_422,
input [18:0] Wgt_6_423,
input [18:0] Wgt_6_424,
input [18:0] Wgt_6_425,
input [18:0] Wgt_6_426,
input [18:0] Wgt_6_427,
input [18:0] Wgt_6_428,
input [18:0] Wgt_6_429,
input [18:0] Wgt_6_430,
input [18:0] Wgt_6_431,
input [18:0] Wgt_6_432,
input [18:0] Wgt_6_433,
input [18:0] Wgt_6_434,
input [18:0] Wgt_6_435,
input [18:0] Wgt_6_436,
input [18:0] Wgt_6_437,
input [18:0] Wgt_6_438,
input [18:0] Wgt_6_439,
input [18:0] Wgt_6_440,
input [18:0] Wgt_6_441,
input [18:0] Wgt_6_442,
input [18:0] Wgt_6_443,
input [18:0] Wgt_6_444,
input [18:0] Wgt_6_445,
input [18:0] Wgt_6_446,
input [18:0] Wgt_6_447,
input [18:0] Wgt_6_448,
input [18:0] Wgt_6_449,
input [18:0] Wgt_6_450,
input [18:0] Wgt_6_451,
input [18:0] Wgt_6_452,
input [18:0] Wgt_6_453,
input [18:0] Wgt_6_454,
input [18:0] Wgt_6_455,
input [18:0] Wgt_6_456,
input [18:0] Wgt_6_457,
input [18:0] Wgt_6_458,
input [18:0] Wgt_6_459,
input [18:0] Wgt_6_460,
input [18:0] Wgt_6_461,
input [18:0] Wgt_6_462,
input [18:0] Wgt_6_463,
input [18:0] Wgt_6_464,
input [18:0] Wgt_6_465,
input [18:0] Wgt_6_466,
input [18:0] Wgt_6_467,
input [18:0] Wgt_6_468,
input [18:0] Wgt_6_469,
input [18:0] Wgt_6_470,
input [18:0] Wgt_6_471,
input [18:0] Wgt_6_472,
input [18:0] Wgt_6_473,
input [18:0] Wgt_6_474,
input [18:0] Wgt_6_475,
input [18:0] Wgt_6_476,
input [18:0] Wgt_6_477,
input [18:0] Wgt_6_478,
input [18:0] Wgt_6_479,
input [18:0] Wgt_6_480,
input [18:0] Wgt_6_481,
input [18:0] Wgt_6_482,
input [18:0] Wgt_6_483,
input [18:0] Wgt_6_484,
input [18:0] Wgt_6_485,
input [18:0] Wgt_6_486,
input [18:0] Wgt_6_487,
input [18:0] Wgt_6_488,
input [18:0] Wgt_6_489,
input [18:0] Wgt_6_490,
input [18:0] Wgt_6_491,
input [18:0] Wgt_6_492,
input [18:0] Wgt_6_493,
input [18:0] Wgt_6_494,
input [18:0] Wgt_6_495,
input [18:0] Wgt_6_496,
input [18:0] Wgt_6_497,
input [18:0] Wgt_6_498,
input [18:0] Wgt_6_499,
input [18:0] Wgt_6_500,
input [18:0] Wgt_6_501,
input [18:0] Wgt_6_502,
input [18:0] Wgt_6_503,
input [18:0] Wgt_6_504,
input [18:0] Wgt_6_505,
input [18:0] Wgt_6_506,
input [18:0] Wgt_6_507,
input [18:0] Wgt_6_508,
input [18:0] Wgt_6_509,
input [18:0] Wgt_6_510,
input [18:0] Wgt_6_511,
input [18:0] Wgt_6_512,
input [18:0] Wgt_6_513,
input [18:0] Wgt_6_514,
input [18:0] Wgt_6_515,
input [18:0] Wgt_6_516,
input [18:0] Wgt_6_517,
input [18:0] Wgt_6_518,
input [18:0] Wgt_6_519,
input [18:0] Wgt_6_520,
input [18:0] Wgt_6_521,
input [18:0] Wgt_6_522,
input [18:0] Wgt_6_523,
input [18:0] Wgt_6_524,
input [18:0] Wgt_6_525,
input [18:0] Wgt_6_526,
input [18:0] Wgt_6_527,
input [18:0] Wgt_6_528,
input [18:0] Wgt_6_529,
input [18:0] Wgt_6_530,
input [18:0] Wgt_6_531,
input [18:0] Wgt_6_532,
input [18:0] Wgt_6_533,
input [18:0] Wgt_6_534,
input [18:0] Wgt_6_535,
input [18:0] Wgt_6_536,
input [18:0] Wgt_6_537,
input [18:0] Wgt_6_538,
input [18:0] Wgt_6_539,
input [18:0] Wgt_6_540,
input [18:0] Wgt_6_541,
input [18:0] Wgt_6_542,
input [18:0] Wgt_6_543,
input [18:0] Wgt_6_544,
input [18:0] Wgt_6_545,
input [18:0] Wgt_6_546,
input [18:0] Wgt_6_547,
input [18:0] Wgt_6_548,
input [18:0] Wgt_6_549,
input [18:0] Wgt_6_550,
input [18:0] Wgt_6_551,
input [18:0] Wgt_6_552,
input [18:0] Wgt_6_553,
input [18:0] Wgt_6_554,
input [18:0] Wgt_6_555,
input [18:0] Wgt_6_556,
input [18:0] Wgt_6_557,
input [18:0] Wgt_6_558,
input [18:0] Wgt_6_559,
input [18:0] Wgt_6_560,
input [18:0] Wgt_6_561,
input [18:0] Wgt_6_562,
input [18:0] Wgt_6_563,
input [18:0] Wgt_6_564,
input [18:0] Wgt_6_565,
input [18:0] Wgt_6_566,
input [18:0] Wgt_6_567,
input [18:0] Wgt_6_568,
input [18:0] Wgt_6_569,
input [18:0] Wgt_6_570,
input [18:0] Wgt_6_571,
input [18:0] Wgt_6_572,
input [18:0] Wgt_6_573,
input [18:0] Wgt_6_574,
input [18:0] Wgt_6_575,
input [18:0] Wgt_6_576,
input [18:0] Wgt_6_577,
input [18:0] Wgt_6_578,
input [18:0] Wgt_6_579,
input [18:0] Wgt_6_580,
input [18:0] Wgt_6_581,
input [18:0] Wgt_6_582,
input [18:0] Wgt_6_583,
input [18:0] Wgt_6_584,
input [18:0] Wgt_6_585,
input [18:0] Wgt_6_586,
input [18:0] Wgt_6_587,
input [18:0] Wgt_6_588,
input [18:0] Wgt_6_589,
input [18:0] Wgt_6_590,
input [18:0] Wgt_6_591,
input [18:0] Wgt_6_592,
input [18:0] Wgt_6_593,
input [18:0] Wgt_6_594,
input [18:0] Wgt_6_595,
input [18:0] Wgt_6_596,
input [18:0] Wgt_6_597,
input [18:0] Wgt_6_598,
input [18:0] Wgt_6_599,
input [18:0] Wgt_6_600,
input [18:0] Wgt_6_601,
input [18:0] Wgt_6_602,
input [18:0] Wgt_6_603,
input [18:0] Wgt_6_604,
input [18:0] Wgt_6_605,
input [18:0] Wgt_6_606,
input [18:0] Wgt_6_607,
input [18:0] Wgt_6_608,
input [18:0] Wgt_6_609,
input [18:0] Wgt_6_610,
input [18:0] Wgt_6_611,
input [18:0] Wgt_6_612,
input [18:0] Wgt_6_613,
input [18:0] Wgt_6_614,
input [18:0] Wgt_6_615,
input [18:0] Wgt_6_616,
input [18:0] Wgt_6_617,
input [18:0] Wgt_6_618,
input [18:0] Wgt_6_619,
input [18:0] Wgt_6_620,
input [18:0] Wgt_6_621,
input [18:0] Wgt_6_622,
input [18:0] Wgt_6_623,
input [18:0] Wgt_6_624,
input [18:0] Wgt_6_625,
input [18:0] Wgt_6_626,
input [18:0] Wgt_6_627,
input [18:0] Wgt_6_628,
input [18:0] Wgt_6_629,
input [18:0] Wgt_6_630,
input [18:0] Wgt_6_631,
input [18:0] Wgt_6_632,
input [18:0] Wgt_6_633,
input [18:0] Wgt_6_634,
input [18:0] Wgt_6_635,
input [18:0] Wgt_6_636,
input [18:0] Wgt_6_637,
input [18:0] Wgt_6_638,
input [18:0] Wgt_6_639,
input [18:0] Wgt_6_640,
input [18:0] Wgt_6_641,
input [18:0] Wgt_6_642,
input [18:0] Wgt_6_643,
input [18:0] Wgt_6_644,
input [18:0] Wgt_6_645,
input [18:0] Wgt_6_646,
input [18:0] Wgt_6_647,
input [18:0] Wgt_6_648,
input [18:0] Wgt_6_649,
input [18:0] Wgt_6_650,
input [18:0] Wgt_6_651,
input [18:0] Wgt_6_652,
input [18:0] Wgt_6_653,
input [18:0] Wgt_6_654,
input [18:0] Wgt_6_655,
input [18:0] Wgt_6_656,
input [18:0] Wgt_6_657,
input [18:0] Wgt_6_658,
input [18:0] Wgt_6_659,
input [18:0] Wgt_6_660,
input [18:0] Wgt_6_661,
input [18:0] Wgt_6_662,
input [18:0] Wgt_6_663,
input [18:0] Wgt_6_664,
input [18:0] Wgt_6_665,
input [18:0] Wgt_6_666,
input [18:0] Wgt_6_667,
input [18:0] Wgt_6_668,
input [18:0] Wgt_6_669,
input [18:0] Wgt_6_670,
input [18:0] Wgt_6_671,
input [18:0] Wgt_6_672,
input [18:0] Wgt_6_673,
input [18:0] Wgt_6_674,
input [18:0] Wgt_6_675,
input [18:0] Wgt_6_676,
input [18:0] Wgt_6_677,
input [18:0] Wgt_6_678,
input [18:0] Wgt_6_679,
input [18:0] Wgt_6_680,
input [18:0] Wgt_6_681,
input [18:0] Wgt_6_682,
input [18:0] Wgt_6_683,
input [18:0] Wgt_6_684,
input [18:0] Wgt_6_685,
input [18:0] Wgt_6_686,
input [18:0] Wgt_6_687,
input [18:0] Wgt_6_688,
input [18:0] Wgt_6_689,
input [18:0] Wgt_6_690,
input [18:0] Wgt_6_691,
input [18:0] Wgt_6_692,
input [18:0] Wgt_6_693,
input [18:0] Wgt_6_694,
input [18:0] Wgt_6_695,
input [18:0] Wgt_6_696,
input [18:0] Wgt_6_697,
input [18:0] Wgt_6_698,
input [18:0] Wgt_6_699,
input [18:0] Wgt_6_700,
input [18:0] Wgt_6_701,
input [18:0] Wgt_6_702,
input [18:0] Wgt_6_703,
input [18:0] Wgt_6_704,
input [18:0] Wgt_6_705,
input [18:0] Wgt_6_706,
input [18:0] Wgt_6_707,
input [18:0] Wgt_6_708,
input [18:0] Wgt_6_709,
input [18:0] Wgt_6_710,
input [18:0] Wgt_6_711,
input [18:0] Wgt_6_712,
input [18:0] Wgt_6_713,
input [18:0] Wgt_6_714,
input [18:0] Wgt_6_715,
input [18:0] Wgt_6_716,
input [18:0] Wgt_6_717,
input [18:0] Wgt_6_718,
input [18:0] Wgt_6_719,
input [18:0] Wgt_6_720,
input [18:0] Wgt_6_721,
input [18:0] Wgt_6_722,
input [18:0] Wgt_6_723,
input [18:0] Wgt_6_724,
input [18:0] Wgt_6_725,
input [18:0] Wgt_6_726,
input [18:0] Wgt_6_727,
input [18:0] Wgt_6_728,
input [18:0] Wgt_6_729,
input [18:0] Wgt_6_730,
input [18:0] Wgt_6_731,
input [18:0] Wgt_6_732,
input [18:0] Wgt_6_733,
input [18:0] Wgt_6_734,
input [18:0] Wgt_6_735,
input [18:0] Wgt_6_736,
input [18:0] Wgt_6_737,
input [18:0] Wgt_6_738,
input [18:0] Wgt_6_739,
input [18:0] Wgt_6_740,
input [18:0] Wgt_6_741,
input [18:0] Wgt_6_742,
input [18:0] Wgt_6_743,
input [18:0] Wgt_6_744,
input [18:0] Wgt_6_745,
input [18:0] Wgt_6_746,
input [18:0] Wgt_6_747,
input [18:0] Wgt_6_748,
input [18:0] Wgt_6_749,
input [18:0] Wgt_6_750,
input [18:0] Wgt_6_751,
input [18:0] Wgt_6_752,
input [18:0] Wgt_6_753,
input [18:0] Wgt_6_754,
input [18:0] Wgt_6_755,
input [18:0] Wgt_6_756,
input [18:0] Wgt_6_757,
input [18:0] Wgt_6_758,
input [18:0] Wgt_6_759,
input [18:0] Wgt_6_760,
input [18:0] Wgt_6_761,
input [18:0] Wgt_6_762,
input [18:0] Wgt_6_763,
input [18:0] Wgt_6_764,
input [18:0] Wgt_6_765,
input [18:0] Wgt_6_766,
input [18:0] Wgt_6_767,
input [18:0] Wgt_6_768,
input [18:0] Wgt_6_769,
input [18:0] Wgt_6_770,
input [18:0] Wgt_6_771,
input [18:0] Wgt_6_772,
input [18:0] Wgt_6_773,
input [18:0] Wgt_6_774,
input [18:0] Wgt_6_775,
input [18:0] Wgt_6_776,
input [18:0] Wgt_6_777,
input [18:0] Wgt_6_778,
input [18:0] Wgt_6_779,
input [18:0] Wgt_6_780,
input [18:0] Wgt_6_781,
input [18:0] Wgt_6_782,
input [18:0] Wgt_6_783,
input [18:0] Wgt_6_784,
input [18:0] Wgt_7_0,
input [18:0] Wgt_7_1,
input [18:0] Wgt_7_2,
input [18:0] Wgt_7_3,
input [18:0] Wgt_7_4,
input [18:0] Wgt_7_5,
input [18:0] Wgt_7_6,
input [18:0] Wgt_7_7,
input [18:0] Wgt_7_8,
input [18:0] Wgt_7_9,
input [18:0] Wgt_7_10,
input [18:0] Wgt_7_11,
input [18:0] Wgt_7_12,
input [18:0] Wgt_7_13,
input [18:0] Wgt_7_14,
input [18:0] Wgt_7_15,
input [18:0] Wgt_7_16,
input [18:0] Wgt_7_17,
input [18:0] Wgt_7_18,
input [18:0] Wgt_7_19,
input [18:0] Wgt_7_20,
input [18:0] Wgt_7_21,
input [18:0] Wgt_7_22,
input [18:0] Wgt_7_23,
input [18:0] Wgt_7_24,
input [18:0] Wgt_7_25,
input [18:0] Wgt_7_26,
input [18:0] Wgt_7_27,
input [18:0] Wgt_7_28,
input [18:0] Wgt_7_29,
input [18:0] Wgt_7_30,
input [18:0] Wgt_7_31,
input [18:0] Wgt_7_32,
input [18:0] Wgt_7_33,
input [18:0] Wgt_7_34,
input [18:0] Wgt_7_35,
input [18:0] Wgt_7_36,
input [18:0] Wgt_7_37,
input [18:0] Wgt_7_38,
input [18:0] Wgt_7_39,
input [18:0] Wgt_7_40,
input [18:0] Wgt_7_41,
input [18:0] Wgt_7_42,
input [18:0] Wgt_7_43,
input [18:0] Wgt_7_44,
input [18:0] Wgt_7_45,
input [18:0] Wgt_7_46,
input [18:0] Wgt_7_47,
input [18:0] Wgt_7_48,
input [18:0] Wgt_7_49,
input [18:0] Wgt_7_50,
input [18:0] Wgt_7_51,
input [18:0] Wgt_7_52,
input [18:0] Wgt_7_53,
input [18:0] Wgt_7_54,
input [18:0] Wgt_7_55,
input [18:0] Wgt_7_56,
input [18:0] Wgt_7_57,
input [18:0] Wgt_7_58,
input [18:0] Wgt_7_59,
input [18:0] Wgt_7_60,
input [18:0] Wgt_7_61,
input [18:0] Wgt_7_62,
input [18:0] Wgt_7_63,
input [18:0] Wgt_7_64,
input [18:0] Wgt_7_65,
input [18:0] Wgt_7_66,
input [18:0] Wgt_7_67,
input [18:0] Wgt_7_68,
input [18:0] Wgt_7_69,
input [18:0] Wgt_7_70,
input [18:0] Wgt_7_71,
input [18:0] Wgt_7_72,
input [18:0] Wgt_7_73,
input [18:0] Wgt_7_74,
input [18:0] Wgt_7_75,
input [18:0] Wgt_7_76,
input [18:0] Wgt_7_77,
input [18:0] Wgt_7_78,
input [18:0] Wgt_7_79,
input [18:0] Wgt_7_80,
input [18:0] Wgt_7_81,
input [18:0] Wgt_7_82,
input [18:0] Wgt_7_83,
input [18:0] Wgt_7_84,
input [18:0] Wgt_7_85,
input [18:0] Wgt_7_86,
input [18:0] Wgt_7_87,
input [18:0] Wgt_7_88,
input [18:0] Wgt_7_89,
input [18:0] Wgt_7_90,
input [18:0] Wgt_7_91,
input [18:0] Wgt_7_92,
input [18:0] Wgt_7_93,
input [18:0] Wgt_7_94,
input [18:0] Wgt_7_95,
input [18:0] Wgt_7_96,
input [18:0] Wgt_7_97,
input [18:0] Wgt_7_98,
input [18:0] Wgt_7_99,
input [18:0] Wgt_7_100,
input [18:0] Wgt_7_101,
input [18:0] Wgt_7_102,
input [18:0] Wgt_7_103,
input [18:0] Wgt_7_104,
input [18:0] Wgt_7_105,
input [18:0] Wgt_7_106,
input [18:0] Wgt_7_107,
input [18:0] Wgt_7_108,
input [18:0] Wgt_7_109,
input [18:0] Wgt_7_110,
input [18:0] Wgt_7_111,
input [18:0] Wgt_7_112,
input [18:0] Wgt_7_113,
input [18:0] Wgt_7_114,
input [18:0] Wgt_7_115,
input [18:0] Wgt_7_116,
input [18:0] Wgt_7_117,
input [18:0] Wgt_7_118,
input [18:0] Wgt_7_119,
input [18:0] Wgt_7_120,
input [18:0] Wgt_7_121,
input [18:0] Wgt_7_122,
input [18:0] Wgt_7_123,
input [18:0] Wgt_7_124,
input [18:0] Wgt_7_125,
input [18:0] Wgt_7_126,
input [18:0] Wgt_7_127,
input [18:0] Wgt_7_128,
input [18:0] Wgt_7_129,
input [18:0] Wgt_7_130,
input [18:0] Wgt_7_131,
input [18:0] Wgt_7_132,
input [18:0] Wgt_7_133,
input [18:0] Wgt_7_134,
input [18:0] Wgt_7_135,
input [18:0] Wgt_7_136,
input [18:0] Wgt_7_137,
input [18:0] Wgt_7_138,
input [18:0] Wgt_7_139,
input [18:0] Wgt_7_140,
input [18:0] Wgt_7_141,
input [18:0] Wgt_7_142,
input [18:0] Wgt_7_143,
input [18:0] Wgt_7_144,
input [18:0] Wgt_7_145,
input [18:0] Wgt_7_146,
input [18:0] Wgt_7_147,
input [18:0] Wgt_7_148,
input [18:0] Wgt_7_149,
input [18:0] Wgt_7_150,
input [18:0] Wgt_7_151,
input [18:0] Wgt_7_152,
input [18:0] Wgt_7_153,
input [18:0] Wgt_7_154,
input [18:0] Wgt_7_155,
input [18:0] Wgt_7_156,
input [18:0] Wgt_7_157,
input [18:0] Wgt_7_158,
input [18:0] Wgt_7_159,
input [18:0] Wgt_7_160,
input [18:0] Wgt_7_161,
input [18:0] Wgt_7_162,
input [18:0] Wgt_7_163,
input [18:0] Wgt_7_164,
input [18:0] Wgt_7_165,
input [18:0] Wgt_7_166,
input [18:0] Wgt_7_167,
input [18:0] Wgt_7_168,
input [18:0] Wgt_7_169,
input [18:0] Wgt_7_170,
input [18:0] Wgt_7_171,
input [18:0] Wgt_7_172,
input [18:0] Wgt_7_173,
input [18:0] Wgt_7_174,
input [18:0] Wgt_7_175,
input [18:0] Wgt_7_176,
input [18:0] Wgt_7_177,
input [18:0] Wgt_7_178,
input [18:0] Wgt_7_179,
input [18:0] Wgt_7_180,
input [18:0] Wgt_7_181,
input [18:0] Wgt_7_182,
input [18:0] Wgt_7_183,
input [18:0] Wgt_7_184,
input [18:0] Wgt_7_185,
input [18:0] Wgt_7_186,
input [18:0] Wgt_7_187,
input [18:0] Wgt_7_188,
input [18:0] Wgt_7_189,
input [18:0] Wgt_7_190,
input [18:0] Wgt_7_191,
input [18:0] Wgt_7_192,
input [18:0] Wgt_7_193,
input [18:0] Wgt_7_194,
input [18:0] Wgt_7_195,
input [18:0] Wgt_7_196,
input [18:0] Wgt_7_197,
input [18:0] Wgt_7_198,
input [18:0] Wgt_7_199,
input [18:0] Wgt_7_200,
input [18:0] Wgt_7_201,
input [18:0] Wgt_7_202,
input [18:0] Wgt_7_203,
input [18:0] Wgt_7_204,
input [18:0] Wgt_7_205,
input [18:0] Wgt_7_206,
input [18:0] Wgt_7_207,
input [18:0] Wgt_7_208,
input [18:0] Wgt_7_209,
input [18:0] Wgt_7_210,
input [18:0] Wgt_7_211,
input [18:0] Wgt_7_212,
input [18:0] Wgt_7_213,
input [18:0] Wgt_7_214,
input [18:0] Wgt_7_215,
input [18:0] Wgt_7_216,
input [18:0] Wgt_7_217,
input [18:0] Wgt_7_218,
input [18:0] Wgt_7_219,
input [18:0] Wgt_7_220,
input [18:0] Wgt_7_221,
input [18:0] Wgt_7_222,
input [18:0] Wgt_7_223,
input [18:0] Wgt_7_224,
input [18:0] Wgt_7_225,
input [18:0] Wgt_7_226,
input [18:0] Wgt_7_227,
input [18:0] Wgt_7_228,
input [18:0] Wgt_7_229,
input [18:0] Wgt_7_230,
input [18:0] Wgt_7_231,
input [18:0] Wgt_7_232,
input [18:0] Wgt_7_233,
input [18:0] Wgt_7_234,
input [18:0] Wgt_7_235,
input [18:0] Wgt_7_236,
input [18:0] Wgt_7_237,
input [18:0] Wgt_7_238,
input [18:0] Wgt_7_239,
input [18:0] Wgt_7_240,
input [18:0] Wgt_7_241,
input [18:0] Wgt_7_242,
input [18:0] Wgt_7_243,
input [18:0] Wgt_7_244,
input [18:0] Wgt_7_245,
input [18:0] Wgt_7_246,
input [18:0] Wgt_7_247,
input [18:0] Wgt_7_248,
input [18:0] Wgt_7_249,
input [18:0] Wgt_7_250,
input [18:0] Wgt_7_251,
input [18:0] Wgt_7_252,
input [18:0] Wgt_7_253,
input [18:0] Wgt_7_254,
input [18:0] Wgt_7_255,
input [18:0] Wgt_7_256,
input [18:0] Wgt_7_257,
input [18:0] Wgt_7_258,
input [18:0] Wgt_7_259,
input [18:0] Wgt_7_260,
input [18:0] Wgt_7_261,
input [18:0] Wgt_7_262,
input [18:0] Wgt_7_263,
input [18:0] Wgt_7_264,
input [18:0] Wgt_7_265,
input [18:0] Wgt_7_266,
input [18:0] Wgt_7_267,
input [18:0] Wgt_7_268,
input [18:0] Wgt_7_269,
input [18:0] Wgt_7_270,
input [18:0] Wgt_7_271,
input [18:0] Wgt_7_272,
input [18:0] Wgt_7_273,
input [18:0] Wgt_7_274,
input [18:0] Wgt_7_275,
input [18:0] Wgt_7_276,
input [18:0] Wgt_7_277,
input [18:0] Wgt_7_278,
input [18:0] Wgt_7_279,
input [18:0] Wgt_7_280,
input [18:0] Wgt_7_281,
input [18:0] Wgt_7_282,
input [18:0] Wgt_7_283,
input [18:0] Wgt_7_284,
input [18:0] Wgt_7_285,
input [18:0] Wgt_7_286,
input [18:0] Wgt_7_287,
input [18:0] Wgt_7_288,
input [18:0] Wgt_7_289,
input [18:0] Wgt_7_290,
input [18:0] Wgt_7_291,
input [18:0] Wgt_7_292,
input [18:0] Wgt_7_293,
input [18:0] Wgt_7_294,
input [18:0] Wgt_7_295,
input [18:0] Wgt_7_296,
input [18:0] Wgt_7_297,
input [18:0] Wgt_7_298,
input [18:0] Wgt_7_299,
input [18:0] Wgt_7_300,
input [18:0] Wgt_7_301,
input [18:0] Wgt_7_302,
input [18:0] Wgt_7_303,
input [18:0] Wgt_7_304,
input [18:0] Wgt_7_305,
input [18:0] Wgt_7_306,
input [18:0] Wgt_7_307,
input [18:0] Wgt_7_308,
input [18:0] Wgt_7_309,
input [18:0] Wgt_7_310,
input [18:0] Wgt_7_311,
input [18:0] Wgt_7_312,
input [18:0] Wgt_7_313,
input [18:0] Wgt_7_314,
input [18:0] Wgt_7_315,
input [18:0] Wgt_7_316,
input [18:0] Wgt_7_317,
input [18:0] Wgt_7_318,
input [18:0] Wgt_7_319,
input [18:0] Wgt_7_320,
input [18:0] Wgt_7_321,
input [18:0] Wgt_7_322,
input [18:0] Wgt_7_323,
input [18:0] Wgt_7_324,
input [18:0] Wgt_7_325,
input [18:0] Wgt_7_326,
input [18:0] Wgt_7_327,
input [18:0] Wgt_7_328,
input [18:0] Wgt_7_329,
input [18:0] Wgt_7_330,
input [18:0] Wgt_7_331,
input [18:0] Wgt_7_332,
input [18:0] Wgt_7_333,
input [18:0] Wgt_7_334,
input [18:0] Wgt_7_335,
input [18:0] Wgt_7_336,
input [18:0] Wgt_7_337,
input [18:0] Wgt_7_338,
input [18:0] Wgt_7_339,
input [18:0] Wgt_7_340,
input [18:0] Wgt_7_341,
input [18:0] Wgt_7_342,
input [18:0] Wgt_7_343,
input [18:0] Wgt_7_344,
input [18:0] Wgt_7_345,
input [18:0] Wgt_7_346,
input [18:0] Wgt_7_347,
input [18:0] Wgt_7_348,
input [18:0] Wgt_7_349,
input [18:0] Wgt_7_350,
input [18:0] Wgt_7_351,
input [18:0] Wgt_7_352,
input [18:0] Wgt_7_353,
input [18:0] Wgt_7_354,
input [18:0] Wgt_7_355,
input [18:0] Wgt_7_356,
input [18:0] Wgt_7_357,
input [18:0] Wgt_7_358,
input [18:0] Wgt_7_359,
input [18:0] Wgt_7_360,
input [18:0] Wgt_7_361,
input [18:0] Wgt_7_362,
input [18:0] Wgt_7_363,
input [18:0] Wgt_7_364,
input [18:0] Wgt_7_365,
input [18:0] Wgt_7_366,
input [18:0] Wgt_7_367,
input [18:0] Wgt_7_368,
input [18:0] Wgt_7_369,
input [18:0] Wgt_7_370,
input [18:0] Wgt_7_371,
input [18:0] Wgt_7_372,
input [18:0] Wgt_7_373,
input [18:0] Wgt_7_374,
input [18:0] Wgt_7_375,
input [18:0] Wgt_7_376,
input [18:0] Wgt_7_377,
input [18:0] Wgt_7_378,
input [18:0] Wgt_7_379,
input [18:0] Wgt_7_380,
input [18:0] Wgt_7_381,
input [18:0] Wgt_7_382,
input [18:0] Wgt_7_383,
input [18:0] Wgt_7_384,
input [18:0] Wgt_7_385,
input [18:0] Wgt_7_386,
input [18:0] Wgt_7_387,
input [18:0] Wgt_7_388,
input [18:0] Wgt_7_389,
input [18:0] Wgt_7_390,
input [18:0] Wgt_7_391,
input [18:0] Wgt_7_392,
input [18:0] Wgt_7_393,
input [18:0] Wgt_7_394,
input [18:0] Wgt_7_395,
input [18:0] Wgt_7_396,
input [18:0] Wgt_7_397,
input [18:0] Wgt_7_398,
input [18:0] Wgt_7_399,
input [18:0] Wgt_7_400,
input [18:0] Wgt_7_401,
input [18:0] Wgt_7_402,
input [18:0] Wgt_7_403,
input [18:0] Wgt_7_404,
input [18:0] Wgt_7_405,
input [18:0] Wgt_7_406,
input [18:0] Wgt_7_407,
input [18:0] Wgt_7_408,
input [18:0] Wgt_7_409,
input [18:0] Wgt_7_410,
input [18:0] Wgt_7_411,
input [18:0] Wgt_7_412,
input [18:0] Wgt_7_413,
input [18:0] Wgt_7_414,
input [18:0] Wgt_7_415,
input [18:0] Wgt_7_416,
input [18:0] Wgt_7_417,
input [18:0] Wgt_7_418,
input [18:0] Wgt_7_419,
input [18:0] Wgt_7_420,
input [18:0] Wgt_7_421,
input [18:0] Wgt_7_422,
input [18:0] Wgt_7_423,
input [18:0] Wgt_7_424,
input [18:0] Wgt_7_425,
input [18:0] Wgt_7_426,
input [18:0] Wgt_7_427,
input [18:0] Wgt_7_428,
input [18:0] Wgt_7_429,
input [18:0] Wgt_7_430,
input [18:0] Wgt_7_431,
input [18:0] Wgt_7_432,
input [18:0] Wgt_7_433,
input [18:0] Wgt_7_434,
input [18:0] Wgt_7_435,
input [18:0] Wgt_7_436,
input [18:0] Wgt_7_437,
input [18:0] Wgt_7_438,
input [18:0] Wgt_7_439,
input [18:0] Wgt_7_440,
input [18:0] Wgt_7_441,
input [18:0] Wgt_7_442,
input [18:0] Wgt_7_443,
input [18:0] Wgt_7_444,
input [18:0] Wgt_7_445,
input [18:0] Wgt_7_446,
input [18:0] Wgt_7_447,
input [18:0] Wgt_7_448,
input [18:0] Wgt_7_449,
input [18:0] Wgt_7_450,
input [18:0] Wgt_7_451,
input [18:0] Wgt_7_452,
input [18:0] Wgt_7_453,
input [18:0] Wgt_7_454,
input [18:0] Wgt_7_455,
input [18:0] Wgt_7_456,
input [18:0] Wgt_7_457,
input [18:0] Wgt_7_458,
input [18:0] Wgt_7_459,
input [18:0] Wgt_7_460,
input [18:0] Wgt_7_461,
input [18:0] Wgt_7_462,
input [18:0] Wgt_7_463,
input [18:0] Wgt_7_464,
input [18:0] Wgt_7_465,
input [18:0] Wgt_7_466,
input [18:0] Wgt_7_467,
input [18:0] Wgt_7_468,
input [18:0] Wgt_7_469,
input [18:0] Wgt_7_470,
input [18:0] Wgt_7_471,
input [18:0] Wgt_7_472,
input [18:0] Wgt_7_473,
input [18:0] Wgt_7_474,
input [18:0] Wgt_7_475,
input [18:0] Wgt_7_476,
input [18:0] Wgt_7_477,
input [18:0] Wgt_7_478,
input [18:0] Wgt_7_479,
input [18:0] Wgt_7_480,
input [18:0] Wgt_7_481,
input [18:0] Wgt_7_482,
input [18:0] Wgt_7_483,
input [18:0] Wgt_7_484,
input [18:0] Wgt_7_485,
input [18:0] Wgt_7_486,
input [18:0] Wgt_7_487,
input [18:0] Wgt_7_488,
input [18:0] Wgt_7_489,
input [18:0] Wgt_7_490,
input [18:0] Wgt_7_491,
input [18:0] Wgt_7_492,
input [18:0] Wgt_7_493,
input [18:0] Wgt_7_494,
input [18:0] Wgt_7_495,
input [18:0] Wgt_7_496,
input [18:0] Wgt_7_497,
input [18:0] Wgt_7_498,
input [18:0] Wgt_7_499,
input [18:0] Wgt_7_500,
input [18:0] Wgt_7_501,
input [18:0] Wgt_7_502,
input [18:0] Wgt_7_503,
input [18:0] Wgt_7_504,
input [18:0] Wgt_7_505,
input [18:0] Wgt_7_506,
input [18:0] Wgt_7_507,
input [18:0] Wgt_7_508,
input [18:0] Wgt_7_509,
input [18:0] Wgt_7_510,
input [18:0] Wgt_7_511,
input [18:0] Wgt_7_512,
input [18:0] Wgt_7_513,
input [18:0] Wgt_7_514,
input [18:0] Wgt_7_515,
input [18:0] Wgt_7_516,
input [18:0] Wgt_7_517,
input [18:0] Wgt_7_518,
input [18:0] Wgt_7_519,
input [18:0] Wgt_7_520,
input [18:0] Wgt_7_521,
input [18:0] Wgt_7_522,
input [18:0] Wgt_7_523,
input [18:0] Wgt_7_524,
input [18:0] Wgt_7_525,
input [18:0] Wgt_7_526,
input [18:0] Wgt_7_527,
input [18:0] Wgt_7_528,
input [18:0] Wgt_7_529,
input [18:0] Wgt_7_530,
input [18:0] Wgt_7_531,
input [18:0] Wgt_7_532,
input [18:0] Wgt_7_533,
input [18:0] Wgt_7_534,
input [18:0] Wgt_7_535,
input [18:0] Wgt_7_536,
input [18:0] Wgt_7_537,
input [18:0] Wgt_7_538,
input [18:0] Wgt_7_539,
input [18:0] Wgt_7_540,
input [18:0] Wgt_7_541,
input [18:0] Wgt_7_542,
input [18:0] Wgt_7_543,
input [18:0] Wgt_7_544,
input [18:0] Wgt_7_545,
input [18:0] Wgt_7_546,
input [18:0] Wgt_7_547,
input [18:0] Wgt_7_548,
input [18:0] Wgt_7_549,
input [18:0] Wgt_7_550,
input [18:0] Wgt_7_551,
input [18:0] Wgt_7_552,
input [18:0] Wgt_7_553,
input [18:0] Wgt_7_554,
input [18:0] Wgt_7_555,
input [18:0] Wgt_7_556,
input [18:0] Wgt_7_557,
input [18:0] Wgt_7_558,
input [18:0] Wgt_7_559,
input [18:0] Wgt_7_560,
input [18:0] Wgt_7_561,
input [18:0] Wgt_7_562,
input [18:0] Wgt_7_563,
input [18:0] Wgt_7_564,
input [18:0] Wgt_7_565,
input [18:0] Wgt_7_566,
input [18:0] Wgt_7_567,
input [18:0] Wgt_7_568,
input [18:0] Wgt_7_569,
input [18:0] Wgt_7_570,
input [18:0] Wgt_7_571,
input [18:0] Wgt_7_572,
input [18:0] Wgt_7_573,
input [18:0] Wgt_7_574,
input [18:0] Wgt_7_575,
input [18:0] Wgt_7_576,
input [18:0] Wgt_7_577,
input [18:0] Wgt_7_578,
input [18:0] Wgt_7_579,
input [18:0] Wgt_7_580,
input [18:0] Wgt_7_581,
input [18:0] Wgt_7_582,
input [18:0] Wgt_7_583,
input [18:0] Wgt_7_584,
input [18:0] Wgt_7_585,
input [18:0] Wgt_7_586,
input [18:0] Wgt_7_587,
input [18:0] Wgt_7_588,
input [18:0] Wgt_7_589,
input [18:0] Wgt_7_590,
input [18:0] Wgt_7_591,
input [18:0] Wgt_7_592,
input [18:0] Wgt_7_593,
input [18:0] Wgt_7_594,
input [18:0] Wgt_7_595,
input [18:0] Wgt_7_596,
input [18:0] Wgt_7_597,
input [18:0] Wgt_7_598,
input [18:0] Wgt_7_599,
input [18:0] Wgt_7_600,
input [18:0] Wgt_7_601,
input [18:0] Wgt_7_602,
input [18:0] Wgt_7_603,
input [18:0] Wgt_7_604,
input [18:0] Wgt_7_605,
input [18:0] Wgt_7_606,
input [18:0] Wgt_7_607,
input [18:0] Wgt_7_608,
input [18:0] Wgt_7_609,
input [18:0] Wgt_7_610,
input [18:0] Wgt_7_611,
input [18:0] Wgt_7_612,
input [18:0] Wgt_7_613,
input [18:0] Wgt_7_614,
input [18:0] Wgt_7_615,
input [18:0] Wgt_7_616,
input [18:0] Wgt_7_617,
input [18:0] Wgt_7_618,
input [18:0] Wgt_7_619,
input [18:0] Wgt_7_620,
input [18:0] Wgt_7_621,
input [18:0] Wgt_7_622,
input [18:0] Wgt_7_623,
input [18:0] Wgt_7_624,
input [18:0] Wgt_7_625,
input [18:0] Wgt_7_626,
input [18:0] Wgt_7_627,
input [18:0] Wgt_7_628,
input [18:0] Wgt_7_629,
input [18:0] Wgt_7_630,
input [18:0] Wgt_7_631,
input [18:0] Wgt_7_632,
input [18:0] Wgt_7_633,
input [18:0] Wgt_7_634,
input [18:0] Wgt_7_635,
input [18:0] Wgt_7_636,
input [18:0] Wgt_7_637,
input [18:0] Wgt_7_638,
input [18:0] Wgt_7_639,
input [18:0] Wgt_7_640,
input [18:0] Wgt_7_641,
input [18:0] Wgt_7_642,
input [18:0] Wgt_7_643,
input [18:0] Wgt_7_644,
input [18:0] Wgt_7_645,
input [18:0] Wgt_7_646,
input [18:0] Wgt_7_647,
input [18:0] Wgt_7_648,
input [18:0] Wgt_7_649,
input [18:0] Wgt_7_650,
input [18:0] Wgt_7_651,
input [18:0] Wgt_7_652,
input [18:0] Wgt_7_653,
input [18:0] Wgt_7_654,
input [18:0] Wgt_7_655,
input [18:0] Wgt_7_656,
input [18:0] Wgt_7_657,
input [18:0] Wgt_7_658,
input [18:0] Wgt_7_659,
input [18:0] Wgt_7_660,
input [18:0] Wgt_7_661,
input [18:0] Wgt_7_662,
input [18:0] Wgt_7_663,
input [18:0] Wgt_7_664,
input [18:0] Wgt_7_665,
input [18:0] Wgt_7_666,
input [18:0] Wgt_7_667,
input [18:0] Wgt_7_668,
input [18:0] Wgt_7_669,
input [18:0] Wgt_7_670,
input [18:0] Wgt_7_671,
input [18:0] Wgt_7_672,
input [18:0] Wgt_7_673,
input [18:0] Wgt_7_674,
input [18:0] Wgt_7_675,
input [18:0] Wgt_7_676,
input [18:0] Wgt_7_677,
input [18:0] Wgt_7_678,
input [18:0] Wgt_7_679,
input [18:0] Wgt_7_680,
input [18:0] Wgt_7_681,
input [18:0] Wgt_7_682,
input [18:0] Wgt_7_683,
input [18:0] Wgt_7_684,
input [18:0] Wgt_7_685,
input [18:0] Wgt_7_686,
input [18:0] Wgt_7_687,
input [18:0] Wgt_7_688,
input [18:0] Wgt_7_689,
input [18:0] Wgt_7_690,
input [18:0] Wgt_7_691,
input [18:0] Wgt_7_692,
input [18:0] Wgt_7_693,
input [18:0] Wgt_7_694,
input [18:0] Wgt_7_695,
input [18:0] Wgt_7_696,
input [18:0] Wgt_7_697,
input [18:0] Wgt_7_698,
input [18:0] Wgt_7_699,
input [18:0] Wgt_7_700,
input [18:0] Wgt_7_701,
input [18:0] Wgt_7_702,
input [18:0] Wgt_7_703,
input [18:0] Wgt_7_704,
input [18:0] Wgt_7_705,
input [18:0] Wgt_7_706,
input [18:0] Wgt_7_707,
input [18:0] Wgt_7_708,
input [18:0] Wgt_7_709,
input [18:0] Wgt_7_710,
input [18:0] Wgt_7_711,
input [18:0] Wgt_7_712,
input [18:0] Wgt_7_713,
input [18:0] Wgt_7_714,
input [18:0] Wgt_7_715,
input [18:0] Wgt_7_716,
input [18:0] Wgt_7_717,
input [18:0] Wgt_7_718,
input [18:0] Wgt_7_719,
input [18:0] Wgt_7_720,
input [18:0] Wgt_7_721,
input [18:0] Wgt_7_722,
input [18:0] Wgt_7_723,
input [18:0] Wgt_7_724,
input [18:0] Wgt_7_725,
input [18:0] Wgt_7_726,
input [18:0] Wgt_7_727,
input [18:0] Wgt_7_728,
input [18:0] Wgt_7_729,
input [18:0] Wgt_7_730,
input [18:0] Wgt_7_731,
input [18:0] Wgt_7_732,
input [18:0] Wgt_7_733,
input [18:0] Wgt_7_734,
input [18:0] Wgt_7_735,
input [18:0] Wgt_7_736,
input [18:0] Wgt_7_737,
input [18:0] Wgt_7_738,
input [18:0] Wgt_7_739,
input [18:0] Wgt_7_740,
input [18:0] Wgt_7_741,
input [18:0] Wgt_7_742,
input [18:0] Wgt_7_743,
input [18:0] Wgt_7_744,
input [18:0] Wgt_7_745,
input [18:0] Wgt_7_746,
input [18:0] Wgt_7_747,
input [18:0] Wgt_7_748,
input [18:0] Wgt_7_749,
input [18:0] Wgt_7_750,
input [18:0] Wgt_7_751,
input [18:0] Wgt_7_752,
input [18:0] Wgt_7_753,
input [18:0] Wgt_7_754,
input [18:0] Wgt_7_755,
input [18:0] Wgt_7_756,
input [18:0] Wgt_7_757,
input [18:0] Wgt_7_758,
input [18:0] Wgt_7_759,
input [18:0] Wgt_7_760,
input [18:0] Wgt_7_761,
input [18:0] Wgt_7_762,
input [18:0] Wgt_7_763,
input [18:0] Wgt_7_764,
input [18:0] Wgt_7_765,
input [18:0] Wgt_7_766,
input [18:0] Wgt_7_767,
input [18:0] Wgt_7_768,
input [18:0] Wgt_7_769,
input [18:0] Wgt_7_770,
input [18:0] Wgt_7_771,
input [18:0] Wgt_7_772,
input [18:0] Wgt_7_773,
input [18:0] Wgt_7_774,
input [18:0] Wgt_7_775,
input [18:0] Wgt_7_776,
input [18:0] Wgt_7_777,
input [18:0] Wgt_7_778,
input [18:0] Wgt_7_779,
input [18:0] Wgt_7_780,
input [18:0] Wgt_7_781,
input [18:0] Wgt_7_782,
input [18:0] Wgt_7_783,
input [18:0] Wgt_7_784,
input [18:0] Wgt_8_0,
input [18:0] Wgt_8_1,
input [18:0] Wgt_8_2,
input [18:0] Wgt_8_3,
input [18:0] Wgt_8_4,
input [18:0] Wgt_8_5,
input [18:0] Wgt_8_6,
input [18:0] Wgt_8_7,
input [18:0] Wgt_8_8,
input [18:0] Wgt_8_9,
input [18:0] Wgt_8_10,
input [18:0] Wgt_8_11,
input [18:0] Wgt_8_12,
input [18:0] Wgt_8_13,
input [18:0] Wgt_8_14,
input [18:0] Wgt_8_15,
input [18:0] Wgt_8_16,
input [18:0] Wgt_8_17,
input [18:0] Wgt_8_18,
input [18:0] Wgt_8_19,
input [18:0] Wgt_8_20,
input [18:0] Wgt_8_21,
input [18:0] Wgt_8_22,
input [18:0] Wgt_8_23,
input [18:0] Wgt_8_24,
input [18:0] Wgt_8_25,
input [18:0] Wgt_8_26,
input [18:0] Wgt_8_27,
input [18:0] Wgt_8_28,
input [18:0] Wgt_8_29,
input [18:0] Wgt_8_30,
input [18:0] Wgt_8_31,
input [18:0] Wgt_8_32,
input [18:0] Wgt_8_33,
input [18:0] Wgt_8_34,
input [18:0] Wgt_8_35,
input [18:0] Wgt_8_36,
input [18:0] Wgt_8_37,
input [18:0] Wgt_8_38,
input [18:0] Wgt_8_39,
input [18:0] Wgt_8_40,
input [18:0] Wgt_8_41,
input [18:0] Wgt_8_42,
input [18:0] Wgt_8_43,
input [18:0] Wgt_8_44,
input [18:0] Wgt_8_45,
input [18:0] Wgt_8_46,
input [18:0] Wgt_8_47,
input [18:0] Wgt_8_48,
input [18:0] Wgt_8_49,
input [18:0] Wgt_8_50,
input [18:0] Wgt_8_51,
input [18:0] Wgt_8_52,
input [18:0] Wgt_8_53,
input [18:0] Wgt_8_54,
input [18:0] Wgt_8_55,
input [18:0] Wgt_8_56,
input [18:0] Wgt_8_57,
input [18:0] Wgt_8_58,
input [18:0] Wgt_8_59,
input [18:0] Wgt_8_60,
input [18:0] Wgt_8_61,
input [18:0] Wgt_8_62,
input [18:0] Wgt_8_63,
input [18:0] Wgt_8_64,
input [18:0] Wgt_8_65,
input [18:0] Wgt_8_66,
input [18:0] Wgt_8_67,
input [18:0] Wgt_8_68,
input [18:0] Wgt_8_69,
input [18:0] Wgt_8_70,
input [18:0] Wgt_8_71,
input [18:0] Wgt_8_72,
input [18:0] Wgt_8_73,
input [18:0] Wgt_8_74,
input [18:0] Wgt_8_75,
input [18:0] Wgt_8_76,
input [18:0] Wgt_8_77,
input [18:0] Wgt_8_78,
input [18:0] Wgt_8_79,
input [18:0] Wgt_8_80,
input [18:0] Wgt_8_81,
input [18:0] Wgt_8_82,
input [18:0] Wgt_8_83,
input [18:0] Wgt_8_84,
input [18:0] Wgt_8_85,
input [18:0] Wgt_8_86,
input [18:0] Wgt_8_87,
input [18:0] Wgt_8_88,
input [18:0] Wgt_8_89,
input [18:0] Wgt_8_90,
input [18:0] Wgt_8_91,
input [18:0] Wgt_8_92,
input [18:0] Wgt_8_93,
input [18:0] Wgt_8_94,
input [18:0] Wgt_8_95,
input [18:0] Wgt_8_96,
input [18:0] Wgt_8_97,
input [18:0] Wgt_8_98,
input [18:0] Wgt_8_99,
input [18:0] Wgt_8_100,
input [18:0] Wgt_8_101,
input [18:0] Wgt_8_102,
input [18:0] Wgt_8_103,
input [18:0] Wgt_8_104,
input [18:0] Wgt_8_105,
input [18:0] Wgt_8_106,
input [18:0] Wgt_8_107,
input [18:0] Wgt_8_108,
input [18:0] Wgt_8_109,
input [18:0] Wgt_8_110,
input [18:0] Wgt_8_111,
input [18:0] Wgt_8_112,
input [18:0] Wgt_8_113,
input [18:0] Wgt_8_114,
input [18:0] Wgt_8_115,
input [18:0] Wgt_8_116,
input [18:0] Wgt_8_117,
input [18:0] Wgt_8_118,
input [18:0] Wgt_8_119,
input [18:0] Wgt_8_120,
input [18:0] Wgt_8_121,
input [18:0] Wgt_8_122,
input [18:0] Wgt_8_123,
input [18:0] Wgt_8_124,
input [18:0] Wgt_8_125,
input [18:0] Wgt_8_126,
input [18:0] Wgt_8_127,
input [18:0] Wgt_8_128,
input [18:0] Wgt_8_129,
input [18:0] Wgt_8_130,
input [18:0] Wgt_8_131,
input [18:0] Wgt_8_132,
input [18:0] Wgt_8_133,
input [18:0] Wgt_8_134,
input [18:0] Wgt_8_135,
input [18:0] Wgt_8_136,
input [18:0] Wgt_8_137,
input [18:0] Wgt_8_138,
input [18:0] Wgt_8_139,
input [18:0] Wgt_8_140,
input [18:0] Wgt_8_141,
input [18:0] Wgt_8_142,
input [18:0] Wgt_8_143,
input [18:0] Wgt_8_144,
input [18:0] Wgt_8_145,
input [18:0] Wgt_8_146,
input [18:0] Wgt_8_147,
input [18:0] Wgt_8_148,
input [18:0] Wgt_8_149,
input [18:0] Wgt_8_150,
input [18:0] Wgt_8_151,
input [18:0] Wgt_8_152,
input [18:0] Wgt_8_153,
input [18:0] Wgt_8_154,
input [18:0] Wgt_8_155,
input [18:0] Wgt_8_156,
input [18:0] Wgt_8_157,
input [18:0] Wgt_8_158,
input [18:0] Wgt_8_159,
input [18:0] Wgt_8_160,
input [18:0] Wgt_8_161,
input [18:0] Wgt_8_162,
input [18:0] Wgt_8_163,
input [18:0] Wgt_8_164,
input [18:0] Wgt_8_165,
input [18:0] Wgt_8_166,
input [18:0] Wgt_8_167,
input [18:0] Wgt_8_168,
input [18:0] Wgt_8_169,
input [18:0] Wgt_8_170,
input [18:0] Wgt_8_171,
input [18:0] Wgt_8_172,
input [18:0] Wgt_8_173,
input [18:0] Wgt_8_174,
input [18:0] Wgt_8_175,
input [18:0] Wgt_8_176,
input [18:0] Wgt_8_177,
input [18:0] Wgt_8_178,
input [18:0] Wgt_8_179,
input [18:0] Wgt_8_180,
input [18:0] Wgt_8_181,
input [18:0] Wgt_8_182,
input [18:0] Wgt_8_183,
input [18:0] Wgt_8_184,
input [18:0] Wgt_8_185,
input [18:0] Wgt_8_186,
input [18:0] Wgt_8_187,
input [18:0] Wgt_8_188,
input [18:0] Wgt_8_189,
input [18:0] Wgt_8_190,
input [18:0] Wgt_8_191,
input [18:0] Wgt_8_192,
input [18:0] Wgt_8_193,
input [18:0] Wgt_8_194,
input [18:0] Wgt_8_195,
input [18:0] Wgt_8_196,
input [18:0] Wgt_8_197,
input [18:0] Wgt_8_198,
input [18:0] Wgt_8_199,
input [18:0] Wgt_8_200,
input [18:0] Wgt_8_201,
input [18:0] Wgt_8_202,
input [18:0] Wgt_8_203,
input [18:0] Wgt_8_204,
input [18:0] Wgt_8_205,
input [18:0] Wgt_8_206,
input [18:0] Wgt_8_207,
input [18:0] Wgt_8_208,
input [18:0] Wgt_8_209,
input [18:0] Wgt_8_210,
input [18:0] Wgt_8_211,
input [18:0] Wgt_8_212,
input [18:0] Wgt_8_213,
input [18:0] Wgt_8_214,
input [18:0] Wgt_8_215,
input [18:0] Wgt_8_216,
input [18:0] Wgt_8_217,
input [18:0] Wgt_8_218,
input [18:0] Wgt_8_219,
input [18:0] Wgt_8_220,
input [18:0] Wgt_8_221,
input [18:0] Wgt_8_222,
input [18:0] Wgt_8_223,
input [18:0] Wgt_8_224,
input [18:0] Wgt_8_225,
input [18:0] Wgt_8_226,
input [18:0] Wgt_8_227,
input [18:0] Wgt_8_228,
input [18:0] Wgt_8_229,
input [18:0] Wgt_8_230,
input [18:0] Wgt_8_231,
input [18:0] Wgt_8_232,
input [18:0] Wgt_8_233,
input [18:0] Wgt_8_234,
input [18:0] Wgt_8_235,
input [18:0] Wgt_8_236,
input [18:0] Wgt_8_237,
input [18:0] Wgt_8_238,
input [18:0] Wgt_8_239,
input [18:0] Wgt_8_240,
input [18:0] Wgt_8_241,
input [18:0] Wgt_8_242,
input [18:0] Wgt_8_243,
input [18:0] Wgt_8_244,
input [18:0] Wgt_8_245,
input [18:0] Wgt_8_246,
input [18:0] Wgt_8_247,
input [18:0] Wgt_8_248,
input [18:0] Wgt_8_249,
input [18:0] Wgt_8_250,
input [18:0] Wgt_8_251,
input [18:0] Wgt_8_252,
input [18:0] Wgt_8_253,
input [18:0] Wgt_8_254,
input [18:0] Wgt_8_255,
input [18:0] Wgt_8_256,
input [18:0] Wgt_8_257,
input [18:0] Wgt_8_258,
input [18:0] Wgt_8_259,
input [18:0] Wgt_8_260,
input [18:0] Wgt_8_261,
input [18:0] Wgt_8_262,
input [18:0] Wgt_8_263,
input [18:0] Wgt_8_264,
input [18:0] Wgt_8_265,
input [18:0] Wgt_8_266,
input [18:0] Wgt_8_267,
input [18:0] Wgt_8_268,
input [18:0] Wgt_8_269,
input [18:0] Wgt_8_270,
input [18:0] Wgt_8_271,
input [18:0] Wgt_8_272,
input [18:0] Wgt_8_273,
input [18:0] Wgt_8_274,
input [18:0] Wgt_8_275,
input [18:0] Wgt_8_276,
input [18:0] Wgt_8_277,
input [18:0] Wgt_8_278,
input [18:0] Wgt_8_279,
input [18:0] Wgt_8_280,
input [18:0] Wgt_8_281,
input [18:0] Wgt_8_282,
input [18:0] Wgt_8_283,
input [18:0] Wgt_8_284,
input [18:0] Wgt_8_285,
input [18:0] Wgt_8_286,
input [18:0] Wgt_8_287,
input [18:0] Wgt_8_288,
input [18:0] Wgt_8_289,
input [18:0] Wgt_8_290,
input [18:0] Wgt_8_291,
input [18:0] Wgt_8_292,
input [18:0] Wgt_8_293,
input [18:0] Wgt_8_294,
input [18:0] Wgt_8_295,
input [18:0] Wgt_8_296,
input [18:0] Wgt_8_297,
input [18:0] Wgt_8_298,
input [18:0] Wgt_8_299,
input [18:0] Wgt_8_300,
input [18:0] Wgt_8_301,
input [18:0] Wgt_8_302,
input [18:0] Wgt_8_303,
input [18:0] Wgt_8_304,
input [18:0] Wgt_8_305,
input [18:0] Wgt_8_306,
input [18:0] Wgt_8_307,
input [18:0] Wgt_8_308,
input [18:0] Wgt_8_309,
input [18:0] Wgt_8_310,
input [18:0] Wgt_8_311,
input [18:0] Wgt_8_312,
input [18:0] Wgt_8_313,
input [18:0] Wgt_8_314,
input [18:0] Wgt_8_315,
input [18:0] Wgt_8_316,
input [18:0] Wgt_8_317,
input [18:0] Wgt_8_318,
input [18:0] Wgt_8_319,
input [18:0] Wgt_8_320,
input [18:0] Wgt_8_321,
input [18:0] Wgt_8_322,
input [18:0] Wgt_8_323,
input [18:0] Wgt_8_324,
input [18:0] Wgt_8_325,
input [18:0] Wgt_8_326,
input [18:0] Wgt_8_327,
input [18:0] Wgt_8_328,
input [18:0] Wgt_8_329,
input [18:0] Wgt_8_330,
input [18:0] Wgt_8_331,
input [18:0] Wgt_8_332,
input [18:0] Wgt_8_333,
input [18:0] Wgt_8_334,
input [18:0] Wgt_8_335,
input [18:0] Wgt_8_336,
input [18:0] Wgt_8_337,
input [18:0] Wgt_8_338,
input [18:0] Wgt_8_339,
input [18:0] Wgt_8_340,
input [18:0] Wgt_8_341,
input [18:0] Wgt_8_342,
input [18:0] Wgt_8_343,
input [18:0] Wgt_8_344,
input [18:0] Wgt_8_345,
input [18:0] Wgt_8_346,
input [18:0] Wgt_8_347,
input [18:0] Wgt_8_348,
input [18:0] Wgt_8_349,
input [18:0] Wgt_8_350,
input [18:0] Wgt_8_351,
input [18:0] Wgt_8_352,
input [18:0] Wgt_8_353,
input [18:0] Wgt_8_354,
input [18:0] Wgt_8_355,
input [18:0] Wgt_8_356,
input [18:0] Wgt_8_357,
input [18:0] Wgt_8_358,
input [18:0] Wgt_8_359,
input [18:0] Wgt_8_360,
input [18:0] Wgt_8_361,
input [18:0] Wgt_8_362,
input [18:0] Wgt_8_363,
input [18:0] Wgt_8_364,
input [18:0] Wgt_8_365,
input [18:0] Wgt_8_366,
input [18:0] Wgt_8_367,
input [18:0] Wgt_8_368,
input [18:0] Wgt_8_369,
input [18:0] Wgt_8_370,
input [18:0] Wgt_8_371,
input [18:0] Wgt_8_372,
input [18:0] Wgt_8_373,
input [18:0] Wgt_8_374,
input [18:0] Wgt_8_375,
input [18:0] Wgt_8_376,
input [18:0] Wgt_8_377,
input [18:0] Wgt_8_378,
input [18:0] Wgt_8_379,
input [18:0] Wgt_8_380,
input [18:0] Wgt_8_381,
input [18:0] Wgt_8_382,
input [18:0] Wgt_8_383,
input [18:0] Wgt_8_384,
input [18:0] Wgt_8_385,
input [18:0] Wgt_8_386,
input [18:0] Wgt_8_387,
input [18:0] Wgt_8_388,
input [18:0] Wgt_8_389,
input [18:0] Wgt_8_390,
input [18:0] Wgt_8_391,
input [18:0] Wgt_8_392,
input [18:0] Wgt_8_393,
input [18:0] Wgt_8_394,
input [18:0] Wgt_8_395,
input [18:0] Wgt_8_396,
input [18:0] Wgt_8_397,
input [18:0] Wgt_8_398,
input [18:0] Wgt_8_399,
input [18:0] Wgt_8_400,
input [18:0] Wgt_8_401,
input [18:0] Wgt_8_402,
input [18:0] Wgt_8_403,
input [18:0] Wgt_8_404,
input [18:0] Wgt_8_405,
input [18:0] Wgt_8_406,
input [18:0] Wgt_8_407,
input [18:0] Wgt_8_408,
input [18:0] Wgt_8_409,
input [18:0] Wgt_8_410,
input [18:0] Wgt_8_411,
input [18:0] Wgt_8_412,
input [18:0] Wgt_8_413,
input [18:0] Wgt_8_414,
input [18:0] Wgt_8_415,
input [18:0] Wgt_8_416,
input [18:0] Wgt_8_417,
input [18:0] Wgt_8_418,
input [18:0] Wgt_8_419,
input [18:0] Wgt_8_420,
input [18:0] Wgt_8_421,
input [18:0] Wgt_8_422,
input [18:0] Wgt_8_423,
input [18:0] Wgt_8_424,
input [18:0] Wgt_8_425,
input [18:0] Wgt_8_426,
input [18:0] Wgt_8_427,
input [18:0] Wgt_8_428,
input [18:0] Wgt_8_429,
input [18:0] Wgt_8_430,
input [18:0] Wgt_8_431,
input [18:0] Wgt_8_432,
input [18:0] Wgt_8_433,
input [18:0] Wgt_8_434,
input [18:0] Wgt_8_435,
input [18:0] Wgt_8_436,
input [18:0] Wgt_8_437,
input [18:0] Wgt_8_438,
input [18:0] Wgt_8_439,
input [18:0] Wgt_8_440,
input [18:0] Wgt_8_441,
input [18:0] Wgt_8_442,
input [18:0] Wgt_8_443,
input [18:0] Wgt_8_444,
input [18:0] Wgt_8_445,
input [18:0] Wgt_8_446,
input [18:0] Wgt_8_447,
input [18:0] Wgt_8_448,
input [18:0] Wgt_8_449,
input [18:0] Wgt_8_450,
input [18:0] Wgt_8_451,
input [18:0] Wgt_8_452,
input [18:0] Wgt_8_453,
input [18:0] Wgt_8_454,
input [18:0] Wgt_8_455,
input [18:0] Wgt_8_456,
input [18:0] Wgt_8_457,
input [18:0] Wgt_8_458,
input [18:0] Wgt_8_459,
input [18:0] Wgt_8_460,
input [18:0] Wgt_8_461,
input [18:0] Wgt_8_462,
input [18:0] Wgt_8_463,
input [18:0] Wgt_8_464,
input [18:0] Wgt_8_465,
input [18:0] Wgt_8_466,
input [18:0] Wgt_8_467,
input [18:0] Wgt_8_468,
input [18:0] Wgt_8_469,
input [18:0] Wgt_8_470,
input [18:0] Wgt_8_471,
input [18:0] Wgt_8_472,
input [18:0] Wgt_8_473,
input [18:0] Wgt_8_474,
input [18:0] Wgt_8_475,
input [18:0] Wgt_8_476,
input [18:0] Wgt_8_477,
input [18:0] Wgt_8_478,
input [18:0] Wgt_8_479,
input [18:0] Wgt_8_480,
input [18:0] Wgt_8_481,
input [18:0] Wgt_8_482,
input [18:0] Wgt_8_483,
input [18:0] Wgt_8_484,
input [18:0] Wgt_8_485,
input [18:0] Wgt_8_486,
input [18:0] Wgt_8_487,
input [18:0] Wgt_8_488,
input [18:0] Wgt_8_489,
input [18:0] Wgt_8_490,
input [18:0] Wgt_8_491,
input [18:0] Wgt_8_492,
input [18:0] Wgt_8_493,
input [18:0] Wgt_8_494,
input [18:0] Wgt_8_495,
input [18:0] Wgt_8_496,
input [18:0] Wgt_8_497,
input [18:0] Wgt_8_498,
input [18:0] Wgt_8_499,
input [18:0] Wgt_8_500,
input [18:0] Wgt_8_501,
input [18:0] Wgt_8_502,
input [18:0] Wgt_8_503,
input [18:0] Wgt_8_504,
input [18:0] Wgt_8_505,
input [18:0] Wgt_8_506,
input [18:0] Wgt_8_507,
input [18:0] Wgt_8_508,
input [18:0] Wgt_8_509,
input [18:0] Wgt_8_510,
input [18:0] Wgt_8_511,
input [18:0] Wgt_8_512,
input [18:0] Wgt_8_513,
input [18:0] Wgt_8_514,
input [18:0] Wgt_8_515,
input [18:0] Wgt_8_516,
input [18:0] Wgt_8_517,
input [18:0] Wgt_8_518,
input [18:0] Wgt_8_519,
input [18:0] Wgt_8_520,
input [18:0] Wgt_8_521,
input [18:0] Wgt_8_522,
input [18:0] Wgt_8_523,
input [18:0] Wgt_8_524,
input [18:0] Wgt_8_525,
input [18:0] Wgt_8_526,
input [18:0] Wgt_8_527,
input [18:0] Wgt_8_528,
input [18:0] Wgt_8_529,
input [18:0] Wgt_8_530,
input [18:0] Wgt_8_531,
input [18:0] Wgt_8_532,
input [18:0] Wgt_8_533,
input [18:0] Wgt_8_534,
input [18:0] Wgt_8_535,
input [18:0] Wgt_8_536,
input [18:0] Wgt_8_537,
input [18:0] Wgt_8_538,
input [18:0] Wgt_8_539,
input [18:0] Wgt_8_540,
input [18:0] Wgt_8_541,
input [18:0] Wgt_8_542,
input [18:0] Wgt_8_543,
input [18:0] Wgt_8_544,
input [18:0] Wgt_8_545,
input [18:0] Wgt_8_546,
input [18:0] Wgt_8_547,
input [18:0] Wgt_8_548,
input [18:0] Wgt_8_549,
input [18:0] Wgt_8_550,
input [18:0] Wgt_8_551,
input [18:0] Wgt_8_552,
input [18:0] Wgt_8_553,
input [18:0] Wgt_8_554,
input [18:0] Wgt_8_555,
input [18:0] Wgt_8_556,
input [18:0] Wgt_8_557,
input [18:0] Wgt_8_558,
input [18:0] Wgt_8_559,
input [18:0] Wgt_8_560,
input [18:0] Wgt_8_561,
input [18:0] Wgt_8_562,
input [18:0] Wgt_8_563,
input [18:0] Wgt_8_564,
input [18:0] Wgt_8_565,
input [18:0] Wgt_8_566,
input [18:0] Wgt_8_567,
input [18:0] Wgt_8_568,
input [18:0] Wgt_8_569,
input [18:0] Wgt_8_570,
input [18:0] Wgt_8_571,
input [18:0] Wgt_8_572,
input [18:0] Wgt_8_573,
input [18:0] Wgt_8_574,
input [18:0] Wgt_8_575,
input [18:0] Wgt_8_576,
input [18:0] Wgt_8_577,
input [18:0] Wgt_8_578,
input [18:0] Wgt_8_579,
input [18:0] Wgt_8_580,
input [18:0] Wgt_8_581,
input [18:0] Wgt_8_582,
input [18:0] Wgt_8_583,
input [18:0] Wgt_8_584,
input [18:0] Wgt_8_585,
input [18:0] Wgt_8_586,
input [18:0] Wgt_8_587,
input [18:0] Wgt_8_588,
input [18:0] Wgt_8_589,
input [18:0] Wgt_8_590,
input [18:0] Wgt_8_591,
input [18:0] Wgt_8_592,
input [18:0] Wgt_8_593,
input [18:0] Wgt_8_594,
input [18:0] Wgt_8_595,
input [18:0] Wgt_8_596,
input [18:0] Wgt_8_597,
input [18:0] Wgt_8_598,
input [18:0] Wgt_8_599,
input [18:0] Wgt_8_600,
input [18:0] Wgt_8_601,
input [18:0] Wgt_8_602,
input [18:0] Wgt_8_603,
input [18:0] Wgt_8_604,
input [18:0] Wgt_8_605,
input [18:0] Wgt_8_606,
input [18:0] Wgt_8_607,
input [18:0] Wgt_8_608,
input [18:0] Wgt_8_609,
input [18:0] Wgt_8_610,
input [18:0] Wgt_8_611,
input [18:0] Wgt_8_612,
input [18:0] Wgt_8_613,
input [18:0] Wgt_8_614,
input [18:0] Wgt_8_615,
input [18:0] Wgt_8_616,
input [18:0] Wgt_8_617,
input [18:0] Wgt_8_618,
input [18:0] Wgt_8_619,
input [18:0] Wgt_8_620,
input [18:0] Wgt_8_621,
input [18:0] Wgt_8_622,
input [18:0] Wgt_8_623,
input [18:0] Wgt_8_624,
input [18:0] Wgt_8_625,
input [18:0] Wgt_8_626,
input [18:0] Wgt_8_627,
input [18:0] Wgt_8_628,
input [18:0] Wgt_8_629,
input [18:0] Wgt_8_630,
input [18:0] Wgt_8_631,
input [18:0] Wgt_8_632,
input [18:0] Wgt_8_633,
input [18:0] Wgt_8_634,
input [18:0] Wgt_8_635,
input [18:0] Wgt_8_636,
input [18:0] Wgt_8_637,
input [18:0] Wgt_8_638,
input [18:0] Wgt_8_639,
input [18:0] Wgt_8_640,
input [18:0] Wgt_8_641,
input [18:0] Wgt_8_642,
input [18:0] Wgt_8_643,
input [18:0] Wgt_8_644,
input [18:0] Wgt_8_645,
input [18:0] Wgt_8_646,
input [18:0] Wgt_8_647,
input [18:0] Wgt_8_648,
input [18:0] Wgt_8_649,
input [18:0] Wgt_8_650,
input [18:0] Wgt_8_651,
input [18:0] Wgt_8_652,
input [18:0] Wgt_8_653,
input [18:0] Wgt_8_654,
input [18:0] Wgt_8_655,
input [18:0] Wgt_8_656,
input [18:0] Wgt_8_657,
input [18:0] Wgt_8_658,
input [18:0] Wgt_8_659,
input [18:0] Wgt_8_660,
input [18:0] Wgt_8_661,
input [18:0] Wgt_8_662,
input [18:0] Wgt_8_663,
input [18:0] Wgt_8_664,
input [18:0] Wgt_8_665,
input [18:0] Wgt_8_666,
input [18:0] Wgt_8_667,
input [18:0] Wgt_8_668,
input [18:0] Wgt_8_669,
input [18:0] Wgt_8_670,
input [18:0] Wgt_8_671,
input [18:0] Wgt_8_672,
input [18:0] Wgt_8_673,
input [18:0] Wgt_8_674,
input [18:0] Wgt_8_675,
input [18:0] Wgt_8_676,
input [18:0] Wgt_8_677,
input [18:0] Wgt_8_678,
input [18:0] Wgt_8_679,
input [18:0] Wgt_8_680,
input [18:0] Wgt_8_681,
input [18:0] Wgt_8_682,
input [18:0] Wgt_8_683,
input [18:0] Wgt_8_684,
input [18:0] Wgt_8_685,
input [18:0] Wgt_8_686,
input [18:0] Wgt_8_687,
input [18:0] Wgt_8_688,
input [18:0] Wgt_8_689,
input [18:0] Wgt_8_690,
input [18:0] Wgt_8_691,
input [18:0] Wgt_8_692,
input [18:0] Wgt_8_693,
input [18:0] Wgt_8_694,
input [18:0] Wgt_8_695,
input [18:0] Wgt_8_696,
input [18:0] Wgt_8_697,
input [18:0] Wgt_8_698,
input [18:0] Wgt_8_699,
input [18:0] Wgt_8_700,
input [18:0] Wgt_8_701,
input [18:0] Wgt_8_702,
input [18:0] Wgt_8_703,
input [18:0] Wgt_8_704,
input [18:0] Wgt_8_705,
input [18:0] Wgt_8_706,
input [18:0] Wgt_8_707,
input [18:0] Wgt_8_708,
input [18:0] Wgt_8_709,
input [18:0] Wgt_8_710,
input [18:0] Wgt_8_711,
input [18:0] Wgt_8_712,
input [18:0] Wgt_8_713,
input [18:0] Wgt_8_714,
input [18:0] Wgt_8_715,
input [18:0] Wgt_8_716,
input [18:0] Wgt_8_717,
input [18:0] Wgt_8_718,
input [18:0] Wgt_8_719,
input [18:0] Wgt_8_720,
input [18:0] Wgt_8_721,
input [18:0] Wgt_8_722,
input [18:0] Wgt_8_723,
input [18:0] Wgt_8_724,
input [18:0] Wgt_8_725,
input [18:0] Wgt_8_726,
input [18:0] Wgt_8_727,
input [18:0] Wgt_8_728,
input [18:0] Wgt_8_729,
input [18:0] Wgt_8_730,
input [18:0] Wgt_8_731,
input [18:0] Wgt_8_732,
input [18:0] Wgt_8_733,
input [18:0] Wgt_8_734,
input [18:0] Wgt_8_735,
input [18:0] Wgt_8_736,
input [18:0] Wgt_8_737,
input [18:0] Wgt_8_738,
input [18:0] Wgt_8_739,
input [18:0] Wgt_8_740,
input [18:0] Wgt_8_741,
input [18:0] Wgt_8_742,
input [18:0] Wgt_8_743,
input [18:0] Wgt_8_744,
input [18:0] Wgt_8_745,
input [18:0] Wgt_8_746,
input [18:0] Wgt_8_747,
input [18:0] Wgt_8_748,
input [18:0] Wgt_8_749,
input [18:0] Wgt_8_750,
input [18:0] Wgt_8_751,
input [18:0] Wgt_8_752,
input [18:0] Wgt_8_753,
input [18:0] Wgt_8_754,
input [18:0] Wgt_8_755,
input [18:0] Wgt_8_756,
input [18:0] Wgt_8_757,
input [18:0] Wgt_8_758,
input [18:0] Wgt_8_759,
input [18:0] Wgt_8_760,
input [18:0] Wgt_8_761,
input [18:0] Wgt_8_762,
input [18:0] Wgt_8_763,
input [18:0] Wgt_8_764,
input [18:0] Wgt_8_765,
input [18:0] Wgt_8_766,
input [18:0] Wgt_8_767,
input [18:0] Wgt_8_768,
input [18:0] Wgt_8_769,
input [18:0] Wgt_8_770,
input [18:0] Wgt_8_771,
input [18:0] Wgt_8_772,
input [18:0] Wgt_8_773,
input [18:0] Wgt_8_774,
input [18:0] Wgt_8_775,
input [18:0] Wgt_8_776,
input [18:0] Wgt_8_777,
input [18:0] Wgt_8_778,
input [18:0] Wgt_8_779,
input [18:0] Wgt_8_780,
input [18:0] Wgt_8_781,
input [18:0] Wgt_8_782,
input [18:0] Wgt_8_783,
input [18:0] Wgt_8_784,
input [18:0] Wgt_9_0,
input [18:0] Wgt_9_1,
input [18:0] Wgt_9_2,
input [18:0] Wgt_9_3,
input [18:0] Wgt_9_4,
input [18:0] Wgt_9_5,
input [18:0] Wgt_9_6,
input [18:0] Wgt_9_7,
input [18:0] Wgt_9_8,
input [18:0] Wgt_9_9,
input [18:0] Wgt_9_10,
input [18:0] Wgt_9_11,
input [18:0] Wgt_9_12,
input [18:0] Wgt_9_13,
input [18:0] Wgt_9_14,
input [18:0] Wgt_9_15,
input [18:0] Wgt_9_16,
input [18:0] Wgt_9_17,
input [18:0] Wgt_9_18,
input [18:0] Wgt_9_19,
input [18:0] Wgt_9_20,
input [18:0] Wgt_9_21,
input [18:0] Wgt_9_22,
input [18:0] Wgt_9_23,
input [18:0] Wgt_9_24,
input [18:0] Wgt_9_25,
input [18:0] Wgt_9_26,
input [18:0] Wgt_9_27,
input [18:0] Wgt_9_28,
input [18:0] Wgt_9_29,
input [18:0] Wgt_9_30,
input [18:0] Wgt_9_31,
input [18:0] Wgt_9_32,
input [18:0] Wgt_9_33,
input [18:0] Wgt_9_34,
input [18:0] Wgt_9_35,
input [18:0] Wgt_9_36,
input [18:0] Wgt_9_37,
input [18:0] Wgt_9_38,
input [18:0] Wgt_9_39,
input [18:0] Wgt_9_40,
input [18:0] Wgt_9_41,
input [18:0] Wgt_9_42,
input [18:0] Wgt_9_43,
input [18:0] Wgt_9_44,
input [18:0] Wgt_9_45,
input [18:0] Wgt_9_46,
input [18:0] Wgt_9_47,
input [18:0] Wgt_9_48,
input [18:0] Wgt_9_49,
input [18:0] Wgt_9_50,
input [18:0] Wgt_9_51,
input [18:0] Wgt_9_52,
input [18:0] Wgt_9_53,
input [18:0] Wgt_9_54,
input [18:0] Wgt_9_55,
input [18:0] Wgt_9_56,
input [18:0] Wgt_9_57,
input [18:0] Wgt_9_58,
input [18:0] Wgt_9_59,
input [18:0] Wgt_9_60,
input [18:0] Wgt_9_61,
input [18:0] Wgt_9_62,
input [18:0] Wgt_9_63,
input [18:0] Wgt_9_64,
input [18:0] Wgt_9_65,
input [18:0] Wgt_9_66,
input [18:0] Wgt_9_67,
input [18:0] Wgt_9_68,
input [18:0] Wgt_9_69,
input [18:0] Wgt_9_70,
input [18:0] Wgt_9_71,
input [18:0] Wgt_9_72,
input [18:0] Wgt_9_73,
input [18:0] Wgt_9_74,
input [18:0] Wgt_9_75,
input [18:0] Wgt_9_76,
input [18:0] Wgt_9_77,
input [18:0] Wgt_9_78,
input [18:0] Wgt_9_79,
input [18:0] Wgt_9_80,
input [18:0] Wgt_9_81,
input [18:0] Wgt_9_82,
input [18:0] Wgt_9_83,
input [18:0] Wgt_9_84,
input [18:0] Wgt_9_85,
input [18:0] Wgt_9_86,
input [18:0] Wgt_9_87,
input [18:0] Wgt_9_88,
input [18:0] Wgt_9_89,
input [18:0] Wgt_9_90,
input [18:0] Wgt_9_91,
input [18:0] Wgt_9_92,
input [18:0] Wgt_9_93,
input [18:0] Wgt_9_94,
input [18:0] Wgt_9_95,
input [18:0] Wgt_9_96,
input [18:0] Wgt_9_97,
input [18:0] Wgt_9_98,
input [18:0] Wgt_9_99,
input [18:0] Wgt_9_100,
input [18:0] Wgt_9_101,
input [18:0] Wgt_9_102,
input [18:0] Wgt_9_103,
input [18:0] Wgt_9_104,
input [18:0] Wgt_9_105,
input [18:0] Wgt_9_106,
input [18:0] Wgt_9_107,
input [18:0] Wgt_9_108,
input [18:0] Wgt_9_109,
input [18:0] Wgt_9_110,
input [18:0] Wgt_9_111,
input [18:0] Wgt_9_112,
input [18:0] Wgt_9_113,
input [18:0] Wgt_9_114,
input [18:0] Wgt_9_115,
input [18:0] Wgt_9_116,
input [18:0] Wgt_9_117,
input [18:0] Wgt_9_118,
input [18:0] Wgt_9_119,
input [18:0] Wgt_9_120,
input [18:0] Wgt_9_121,
input [18:0] Wgt_9_122,
input [18:0] Wgt_9_123,
input [18:0] Wgt_9_124,
input [18:0] Wgt_9_125,
input [18:0] Wgt_9_126,
input [18:0] Wgt_9_127,
input [18:0] Wgt_9_128,
input [18:0] Wgt_9_129,
input [18:0] Wgt_9_130,
input [18:0] Wgt_9_131,
input [18:0] Wgt_9_132,
input [18:0] Wgt_9_133,
input [18:0] Wgt_9_134,
input [18:0] Wgt_9_135,
input [18:0] Wgt_9_136,
input [18:0] Wgt_9_137,
input [18:0] Wgt_9_138,
input [18:0] Wgt_9_139,
input [18:0] Wgt_9_140,
input [18:0] Wgt_9_141,
input [18:0] Wgt_9_142,
input [18:0] Wgt_9_143,
input [18:0] Wgt_9_144,
input [18:0] Wgt_9_145,
input [18:0] Wgt_9_146,
input [18:0] Wgt_9_147,
input [18:0] Wgt_9_148,
input [18:0] Wgt_9_149,
input [18:0] Wgt_9_150,
input [18:0] Wgt_9_151,
input [18:0] Wgt_9_152,
input [18:0] Wgt_9_153,
input [18:0] Wgt_9_154,
input [18:0] Wgt_9_155,
input [18:0] Wgt_9_156,
input [18:0] Wgt_9_157,
input [18:0] Wgt_9_158,
input [18:0] Wgt_9_159,
input [18:0] Wgt_9_160,
input [18:0] Wgt_9_161,
input [18:0] Wgt_9_162,
input [18:0] Wgt_9_163,
input [18:0] Wgt_9_164,
input [18:0] Wgt_9_165,
input [18:0] Wgt_9_166,
input [18:0] Wgt_9_167,
input [18:0] Wgt_9_168,
input [18:0] Wgt_9_169,
input [18:0] Wgt_9_170,
input [18:0] Wgt_9_171,
input [18:0] Wgt_9_172,
input [18:0] Wgt_9_173,
input [18:0] Wgt_9_174,
input [18:0] Wgt_9_175,
input [18:0] Wgt_9_176,
input [18:0] Wgt_9_177,
input [18:0] Wgt_9_178,
input [18:0] Wgt_9_179,
input [18:0] Wgt_9_180,
input [18:0] Wgt_9_181,
input [18:0] Wgt_9_182,
input [18:0] Wgt_9_183,
input [18:0] Wgt_9_184,
input [18:0] Wgt_9_185,
input [18:0] Wgt_9_186,
input [18:0] Wgt_9_187,
input [18:0] Wgt_9_188,
input [18:0] Wgt_9_189,
input [18:0] Wgt_9_190,
input [18:0] Wgt_9_191,
input [18:0] Wgt_9_192,
input [18:0] Wgt_9_193,
input [18:0] Wgt_9_194,
input [18:0] Wgt_9_195,
input [18:0] Wgt_9_196,
input [18:0] Wgt_9_197,
input [18:0] Wgt_9_198,
input [18:0] Wgt_9_199,
input [18:0] Wgt_9_200,
input [18:0] Wgt_9_201,
input [18:0] Wgt_9_202,
input [18:0] Wgt_9_203,
input [18:0] Wgt_9_204,
input [18:0] Wgt_9_205,
input [18:0] Wgt_9_206,
input [18:0] Wgt_9_207,
input [18:0] Wgt_9_208,
input [18:0] Wgt_9_209,
input [18:0] Wgt_9_210,
input [18:0] Wgt_9_211,
input [18:0] Wgt_9_212,
input [18:0] Wgt_9_213,
input [18:0] Wgt_9_214,
input [18:0] Wgt_9_215,
input [18:0] Wgt_9_216,
input [18:0] Wgt_9_217,
input [18:0] Wgt_9_218,
input [18:0] Wgt_9_219,
input [18:0] Wgt_9_220,
input [18:0] Wgt_9_221,
input [18:0] Wgt_9_222,
input [18:0] Wgt_9_223,
input [18:0] Wgt_9_224,
input [18:0] Wgt_9_225,
input [18:0] Wgt_9_226,
input [18:0] Wgt_9_227,
input [18:0] Wgt_9_228,
input [18:0] Wgt_9_229,
input [18:0] Wgt_9_230,
input [18:0] Wgt_9_231,
input [18:0] Wgt_9_232,
input [18:0] Wgt_9_233,
input [18:0] Wgt_9_234,
input [18:0] Wgt_9_235,
input [18:0] Wgt_9_236,
input [18:0] Wgt_9_237,
input [18:0] Wgt_9_238,
input [18:0] Wgt_9_239,
input [18:0] Wgt_9_240,
input [18:0] Wgt_9_241,
input [18:0] Wgt_9_242,
input [18:0] Wgt_9_243,
input [18:0] Wgt_9_244,
input [18:0] Wgt_9_245,
input [18:0] Wgt_9_246,
input [18:0] Wgt_9_247,
input [18:0] Wgt_9_248,
input [18:0] Wgt_9_249,
input [18:0] Wgt_9_250,
input [18:0] Wgt_9_251,
input [18:0] Wgt_9_252,
input [18:0] Wgt_9_253,
input [18:0] Wgt_9_254,
input [18:0] Wgt_9_255,
input [18:0] Wgt_9_256,
input [18:0] Wgt_9_257,
input [18:0] Wgt_9_258,
input [18:0] Wgt_9_259,
input [18:0] Wgt_9_260,
input [18:0] Wgt_9_261,
input [18:0] Wgt_9_262,
input [18:0] Wgt_9_263,
input [18:0] Wgt_9_264,
input [18:0] Wgt_9_265,
input [18:0] Wgt_9_266,
input [18:0] Wgt_9_267,
input [18:0] Wgt_9_268,
input [18:0] Wgt_9_269,
input [18:0] Wgt_9_270,
input [18:0] Wgt_9_271,
input [18:0] Wgt_9_272,
input [18:0] Wgt_9_273,
input [18:0] Wgt_9_274,
input [18:0] Wgt_9_275,
input [18:0] Wgt_9_276,
input [18:0] Wgt_9_277,
input [18:0] Wgt_9_278,
input [18:0] Wgt_9_279,
input [18:0] Wgt_9_280,
input [18:0] Wgt_9_281,
input [18:0] Wgt_9_282,
input [18:0] Wgt_9_283,
input [18:0] Wgt_9_284,
input [18:0] Wgt_9_285,
input [18:0] Wgt_9_286,
input [18:0] Wgt_9_287,
input [18:0] Wgt_9_288,
input [18:0] Wgt_9_289,
input [18:0] Wgt_9_290,
input [18:0] Wgt_9_291,
input [18:0] Wgt_9_292,
input [18:0] Wgt_9_293,
input [18:0] Wgt_9_294,
input [18:0] Wgt_9_295,
input [18:0] Wgt_9_296,
input [18:0] Wgt_9_297,
input [18:0] Wgt_9_298,
input [18:0] Wgt_9_299,
input [18:0] Wgt_9_300,
input [18:0] Wgt_9_301,
input [18:0] Wgt_9_302,
input [18:0] Wgt_9_303,
input [18:0] Wgt_9_304,
input [18:0] Wgt_9_305,
input [18:0] Wgt_9_306,
input [18:0] Wgt_9_307,
input [18:0] Wgt_9_308,
input [18:0] Wgt_9_309,
input [18:0] Wgt_9_310,
input [18:0] Wgt_9_311,
input [18:0] Wgt_9_312,
input [18:0] Wgt_9_313,
input [18:0] Wgt_9_314,
input [18:0] Wgt_9_315,
input [18:0] Wgt_9_316,
input [18:0] Wgt_9_317,
input [18:0] Wgt_9_318,
input [18:0] Wgt_9_319,
input [18:0] Wgt_9_320,
input [18:0] Wgt_9_321,
input [18:0] Wgt_9_322,
input [18:0] Wgt_9_323,
input [18:0] Wgt_9_324,
input [18:0] Wgt_9_325,
input [18:0] Wgt_9_326,
input [18:0] Wgt_9_327,
input [18:0] Wgt_9_328,
input [18:0] Wgt_9_329,
input [18:0] Wgt_9_330,
input [18:0] Wgt_9_331,
input [18:0] Wgt_9_332,
input [18:0] Wgt_9_333,
input [18:0] Wgt_9_334,
input [18:0] Wgt_9_335,
input [18:0] Wgt_9_336,
input [18:0] Wgt_9_337,
input [18:0] Wgt_9_338,
input [18:0] Wgt_9_339,
input [18:0] Wgt_9_340,
input [18:0] Wgt_9_341,
input [18:0] Wgt_9_342,
input [18:0] Wgt_9_343,
input [18:0] Wgt_9_344,
input [18:0] Wgt_9_345,
input [18:0] Wgt_9_346,
input [18:0] Wgt_9_347,
input [18:0] Wgt_9_348,
input [18:0] Wgt_9_349,
input [18:0] Wgt_9_350,
input [18:0] Wgt_9_351,
input [18:0] Wgt_9_352,
input [18:0] Wgt_9_353,
input [18:0] Wgt_9_354,
input [18:0] Wgt_9_355,
input [18:0] Wgt_9_356,
input [18:0] Wgt_9_357,
input [18:0] Wgt_9_358,
input [18:0] Wgt_9_359,
input [18:0] Wgt_9_360,
input [18:0] Wgt_9_361,
input [18:0] Wgt_9_362,
input [18:0] Wgt_9_363,
input [18:0] Wgt_9_364,
input [18:0] Wgt_9_365,
input [18:0] Wgt_9_366,
input [18:0] Wgt_9_367,
input [18:0] Wgt_9_368,
input [18:0] Wgt_9_369,
input [18:0] Wgt_9_370,
input [18:0] Wgt_9_371,
input [18:0] Wgt_9_372,
input [18:0] Wgt_9_373,
input [18:0] Wgt_9_374,
input [18:0] Wgt_9_375,
input [18:0] Wgt_9_376,
input [18:0] Wgt_9_377,
input [18:0] Wgt_9_378,
input [18:0] Wgt_9_379,
input [18:0] Wgt_9_380,
input [18:0] Wgt_9_381,
input [18:0] Wgt_9_382,
input [18:0] Wgt_9_383,
input [18:0] Wgt_9_384,
input [18:0] Wgt_9_385,
input [18:0] Wgt_9_386,
input [18:0] Wgt_9_387,
input [18:0] Wgt_9_388,
input [18:0] Wgt_9_389,
input [18:0] Wgt_9_390,
input [18:0] Wgt_9_391,
input [18:0] Wgt_9_392,
input [18:0] Wgt_9_393,
input [18:0] Wgt_9_394,
input [18:0] Wgt_9_395,
input [18:0] Wgt_9_396,
input [18:0] Wgt_9_397,
input [18:0] Wgt_9_398,
input [18:0] Wgt_9_399,
input [18:0] Wgt_9_400,
input [18:0] Wgt_9_401,
input [18:0] Wgt_9_402,
input [18:0] Wgt_9_403,
input [18:0] Wgt_9_404,
input [18:0] Wgt_9_405,
input [18:0] Wgt_9_406,
input [18:0] Wgt_9_407,
input [18:0] Wgt_9_408,
input [18:0] Wgt_9_409,
input [18:0] Wgt_9_410,
input [18:0] Wgt_9_411,
input [18:0] Wgt_9_412,
input [18:0] Wgt_9_413,
input [18:0] Wgt_9_414,
input [18:0] Wgt_9_415,
input [18:0] Wgt_9_416,
input [18:0] Wgt_9_417,
input [18:0] Wgt_9_418,
input [18:0] Wgt_9_419,
input [18:0] Wgt_9_420,
input [18:0] Wgt_9_421,
input [18:0] Wgt_9_422,
input [18:0] Wgt_9_423,
input [18:0] Wgt_9_424,
input [18:0] Wgt_9_425,
input [18:0] Wgt_9_426,
input [18:0] Wgt_9_427,
input [18:0] Wgt_9_428,
input [18:0] Wgt_9_429,
input [18:0] Wgt_9_430,
input [18:0] Wgt_9_431,
input [18:0] Wgt_9_432,
input [18:0] Wgt_9_433,
input [18:0] Wgt_9_434,
input [18:0] Wgt_9_435,
input [18:0] Wgt_9_436,
input [18:0] Wgt_9_437,
input [18:0] Wgt_9_438,
input [18:0] Wgt_9_439,
input [18:0] Wgt_9_440,
input [18:0] Wgt_9_441,
input [18:0] Wgt_9_442,
input [18:0] Wgt_9_443,
input [18:0] Wgt_9_444,
input [18:0] Wgt_9_445,
input [18:0] Wgt_9_446,
input [18:0] Wgt_9_447,
input [18:0] Wgt_9_448,
input [18:0] Wgt_9_449,
input [18:0] Wgt_9_450,
input [18:0] Wgt_9_451,
input [18:0] Wgt_9_452,
input [18:0] Wgt_9_453,
input [18:0] Wgt_9_454,
input [18:0] Wgt_9_455,
input [18:0] Wgt_9_456,
input [18:0] Wgt_9_457,
input [18:0] Wgt_9_458,
input [18:0] Wgt_9_459,
input [18:0] Wgt_9_460,
input [18:0] Wgt_9_461,
input [18:0] Wgt_9_462,
input [18:0] Wgt_9_463,
input [18:0] Wgt_9_464,
input [18:0] Wgt_9_465,
input [18:0] Wgt_9_466,
input [18:0] Wgt_9_467,
input [18:0] Wgt_9_468,
input [18:0] Wgt_9_469,
input [18:0] Wgt_9_470,
input [18:0] Wgt_9_471,
input [18:0] Wgt_9_472,
input [18:0] Wgt_9_473,
input [18:0] Wgt_9_474,
input [18:0] Wgt_9_475,
input [18:0] Wgt_9_476,
input [18:0] Wgt_9_477,
input [18:0] Wgt_9_478,
input [18:0] Wgt_9_479,
input [18:0] Wgt_9_480,
input [18:0] Wgt_9_481,
input [18:0] Wgt_9_482,
input [18:0] Wgt_9_483,
input [18:0] Wgt_9_484,
input [18:0] Wgt_9_485,
input [18:0] Wgt_9_486,
input [18:0] Wgt_9_487,
input [18:0] Wgt_9_488,
input [18:0] Wgt_9_489,
input [18:0] Wgt_9_490,
input [18:0] Wgt_9_491,
input [18:0] Wgt_9_492,
input [18:0] Wgt_9_493,
input [18:0] Wgt_9_494,
input [18:0] Wgt_9_495,
input [18:0] Wgt_9_496,
input [18:0] Wgt_9_497,
input [18:0] Wgt_9_498,
input [18:0] Wgt_9_499,
input [18:0] Wgt_9_500,
input [18:0] Wgt_9_501,
input [18:0] Wgt_9_502,
input [18:0] Wgt_9_503,
input [18:0] Wgt_9_504,
input [18:0] Wgt_9_505,
input [18:0] Wgt_9_506,
input [18:0] Wgt_9_507,
input [18:0] Wgt_9_508,
input [18:0] Wgt_9_509,
input [18:0] Wgt_9_510,
input [18:0] Wgt_9_511,
input [18:0] Wgt_9_512,
input [18:0] Wgt_9_513,
input [18:0] Wgt_9_514,
input [18:0] Wgt_9_515,
input [18:0] Wgt_9_516,
input [18:0] Wgt_9_517,
input [18:0] Wgt_9_518,
input [18:0] Wgt_9_519,
input [18:0] Wgt_9_520,
input [18:0] Wgt_9_521,
input [18:0] Wgt_9_522,
input [18:0] Wgt_9_523,
input [18:0] Wgt_9_524,
input [18:0] Wgt_9_525,
input [18:0] Wgt_9_526,
input [18:0] Wgt_9_527,
input [18:0] Wgt_9_528,
input [18:0] Wgt_9_529,
input [18:0] Wgt_9_530,
input [18:0] Wgt_9_531,
input [18:0] Wgt_9_532,
input [18:0] Wgt_9_533,
input [18:0] Wgt_9_534,
input [18:0] Wgt_9_535,
input [18:0] Wgt_9_536,
input [18:0] Wgt_9_537,
input [18:0] Wgt_9_538,
input [18:0] Wgt_9_539,
input [18:0] Wgt_9_540,
input [18:0] Wgt_9_541,
input [18:0] Wgt_9_542,
input [18:0] Wgt_9_543,
input [18:0] Wgt_9_544,
input [18:0] Wgt_9_545,
input [18:0] Wgt_9_546,
input [18:0] Wgt_9_547,
input [18:0] Wgt_9_548,
input [18:0] Wgt_9_549,
input [18:0] Wgt_9_550,
input [18:0] Wgt_9_551,
input [18:0] Wgt_9_552,
input [18:0] Wgt_9_553,
input [18:0] Wgt_9_554,
input [18:0] Wgt_9_555,
input [18:0] Wgt_9_556,
input [18:0] Wgt_9_557,
input [18:0] Wgt_9_558,
input [18:0] Wgt_9_559,
input [18:0] Wgt_9_560,
input [18:0] Wgt_9_561,
input [18:0] Wgt_9_562,
input [18:0] Wgt_9_563,
input [18:0] Wgt_9_564,
input [18:0] Wgt_9_565,
input [18:0] Wgt_9_566,
input [18:0] Wgt_9_567,
input [18:0] Wgt_9_568,
input [18:0] Wgt_9_569,
input [18:0] Wgt_9_570,
input [18:0] Wgt_9_571,
input [18:0] Wgt_9_572,
input [18:0] Wgt_9_573,
input [18:0] Wgt_9_574,
input [18:0] Wgt_9_575,
input [18:0] Wgt_9_576,
input [18:0] Wgt_9_577,
input [18:0] Wgt_9_578,
input [18:0] Wgt_9_579,
input [18:0] Wgt_9_580,
input [18:0] Wgt_9_581,
input [18:0] Wgt_9_582,
input [18:0] Wgt_9_583,
input [18:0] Wgt_9_584,
input [18:0] Wgt_9_585,
input [18:0] Wgt_9_586,
input [18:0] Wgt_9_587,
input [18:0] Wgt_9_588,
input [18:0] Wgt_9_589,
input [18:0] Wgt_9_590,
input [18:0] Wgt_9_591,
input [18:0] Wgt_9_592,
input [18:0] Wgt_9_593,
input [18:0] Wgt_9_594,
input [18:0] Wgt_9_595,
input [18:0] Wgt_9_596,
input [18:0] Wgt_9_597,
input [18:0] Wgt_9_598,
input [18:0] Wgt_9_599,
input [18:0] Wgt_9_600,
input [18:0] Wgt_9_601,
input [18:0] Wgt_9_602,
input [18:0] Wgt_9_603,
input [18:0] Wgt_9_604,
input [18:0] Wgt_9_605,
input [18:0] Wgt_9_606,
input [18:0] Wgt_9_607,
input [18:0] Wgt_9_608,
input [18:0] Wgt_9_609,
input [18:0] Wgt_9_610,
input [18:0] Wgt_9_611,
input [18:0] Wgt_9_612,
input [18:0] Wgt_9_613,
input [18:0] Wgt_9_614,
input [18:0] Wgt_9_615,
input [18:0] Wgt_9_616,
input [18:0] Wgt_9_617,
input [18:0] Wgt_9_618,
input [18:0] Wgt_9_619,
input [18:0] Wgt_9_620,
input [18:0] Wgt_9_621,
input [18:0] Wgt_9_622,
input [18:0] Wgt_9_623,
input [18:0] Wgt_9_624,
input [18:0] Wgt_9_625,
input [18:0] Wgt_9_626,
input [18:0] Wgt_9_627,
input [18:0] Wgt_9_628,
input [18:0] Wgt_9_629,
input [18:0] Wgt_9_630,
input [18:0] Wgt_9_631,
input [18:0] Wgt_9_632,
input [18:0] Wgt_9_633,
input [18:0] Wgt_9_634,
input [18:0] Wgt_9_635,
input [18:0] Wgt_9_636,
input [18:0] Wgt_9_637,
input [18:0] Wgt_9_638,
input [18:0] Wgt_9_639,
input [18:0] Wgt_9_640,
input [18:0] Wgt_9_641,
input [18:0] Wgt_9_642,
input [18:0] Wgt_9_643,
input [18:0] Wgt_9_644,
input [18:0] Wgt_9_645,
input [18:0] Wgt_9_646,
input [18:0] Wgt_9_647,
input [18:0] Wgt_9_648,
input [18:0] Wgt_9_649,
input [18:0] Wgt_9_650,
input [18:0] Wgt_9_651,
input [18:0] Wgt_9_652,
input [18:0] Wgt_9_653,
input [18:0] Wgt_9_654,
input [18:0] Wgt_9_655,
input [18:0] Wgt_9_656,
input [18:0] Wgt_9_657,
input [18:0] Wgt_9_658,
input [18:0] Wgt_9_659,
input [18:0] Wgt_9_660,
input [18:0] Wgt_9_661,
input [18:0] Wgt_9_662,
input [18:0] Wgt_9_663,
input [18:0] Wgt_9_664,
input [18:0] Wgt_9_665,
input [18:0] Wgt_9_666,
input [18:0] Wgt_9_667,
input [18:0] Wgt_9_668,
input [18:0] Wgt_9_669,
input [18:0] Wgt_9_670,
input [18:0] Wgt_9_671,
input [18:0] Wgt_9_672,
input [18:0] Wgt_9_673,
input [18:0] Wgt_9_674,
input [18:0] Wgt_9_675,
input [18:0] Wgt_9_676,
input [18:0] Wgt_9_677,
input [18:0] Wgt_9_678,
input [18:0] Wgt_9_679,
input [18:0] Wgt_9_680,
input [18:0] Wgt_9_681,
input [18:0] Wgt_9_682,
input [18:0] Wgt_9_683,
input [18:0] Wgt_9_684,
input [18:0] Wgt_9_685,
input [18:0] Wgt_9_686,
input [18:0] Wgt_9_687,
input [18:0] Wgt_9_688,
input [18:0] Wgt_9_689,
input [18:0] Wgt_9_690,
input [18:0] Wgt_9_691,
input [18:0] Wgt_9_692,
input [18:0] Wgt_9_693,
input [18:0] Wgt_9_694,
input [18:0] Wgt_9_695,
input [18:0] Wgt_9_696,
input [18:0] Wgt_9_697,
input [18:0] Wgt_9_698,
input [18:0] Wgt_9_699,
input [18:0] Wgt_9_700,
input [18:0] Wgt_9_701,
input [18:0] Wgt_9_702,
input [18:0] Wgt_9_703,
input [18:0] Wgt_9_704,
input [18:0] Wgt_9_705,
input [18:0] Wgt_9_706,
input [18:0] Wgt_9_707,
input [18:0] Wgt_9_708,
input [18:0] Wgt_9_709,
input [18:0] Wgt_9_710,
input [18:0] Wgt_9_711,
input [18:0] Wgt_9_712,
input [18:0] Wgt_9_713,
input [18:0] Wgt_9_714,
input [18:0] Wgt_9_715,
input [18:0] Wgt_9_716,
input [18:0] Wgt_9_717,
input [18:0] Wgt_9_718,
input [18:0] Wgt_9_719,
input [18:0] Wgt_9_720,
input [18:0] Wgt_9_721,
input [18:0] Wgt_9_722,
input [18:0] Wgt_9_723,
input [18:0] Wgt_9_724,
input [18:0] Wgt_9_725,
input [18:0] Wgt_9_726,
input [18:0] Wgt_9_727,
input [18:0] Wgt_9_728,
input [18:0] Wgt_9_729,
input [18:0] Wgt_9_730,
input [18:0] Wgt_9_731,
input [18:0] Wgt_9_732,
input [18:0] Wgt_9_733,
input [18:0] Wgt_9_734,
input [18:0] Wgt_9_735,
input [18:0] Wgt_9_736,
input [18:0] Wgt_9_737,
input [18:0] Wgt_9_738,
input [18:0] Wgt_9_739,
input [18:0] Wgt_9_740,
input [18:0] Wgt_9_741,
input [18:0] Wgt_9_742,
input [18:0] Wgt_9_743,
input [18:0] Wgt_9_744,
input [18:0] Wgt_9_745,
input [18:0] Wgt_9_746,
input [18:0] Wgt_9_747,
input [18:0] Wgt_9_748,
input [18:0] Wgt_9_749,
input [18:0] Wgt_9_750,
input [18:0] Wgt_9_751,
input [18:0] Wgt_9_752,
input [18:0] Wgt_9_753,
input [18:0] Wgt_9_754,
input [18:0] Wgt_9_755,
input [18:0] Wgt_9_756,
input [18:0] Wgt_9_757,
input [18:0] Wgt_9_758,
input [18:0] Wgt_9_759,
input [18:0] Wgt_9_760,
input [18:0] Wgt_9_761,
input [18:0] Wgt_9_762,
input [18:0] Wgt_9_763,
input [18:0] Wgt_9_764,
input [18:0] Wgt_9_765,
input [18:0] Wgt_9_766,
input [18:0] Wgt_9_767,
input [18:0] Wgt_9_768,
input [18:0] Wgt_9_769,
input [18:0] Wgt_9_770,
input [18:0] Wgt_9_771,
input [18:0] Wgt_9_772,
input [18:0] Wgt_9_773,
input [18:0] Wgt_9_774,
input [18:0] Wgt_9_775,
input [18:0] Wgt_9_776,
input [18:0] Wgt_9_777,
input [18:0] Wgt_9_778,
input [18:0] Wgt_9_779,
input [18:0] Wgt_9_780,
input [18:0] Wgt_9_781,
input [18:0] Wgt_9_782,
input [18:0] Wgt_9_783,
input [18:0] Wgt_9_784,
input [9:0] Pix_0,
input [9:0] Pix_1,
input [9:0] Pix_2,
input [9:0] Pix_3,
input [9:0] Pix_4,
input [9:0] Pix_5,
input [9:0] Pix_6,
input [9:0] Pix_7,
input [9:0] Pix_8,
input [9:0] Pix_9,
input [9:0] Pix_10,
input [9:0] Pix_11,
input [9:0] Pix_12,
input [9:0] Pix_13,
input [9:0] Pix_14,
input [9:0] Pix_15,
input [9:0] Pix_16,
input [9:0] Pix_17,
input [9:0] Pix_18,
input [9:0] Pix_19,
input [9:0] Pix_20,
input [9:0] Pix_21,
input [9:0] Pix_22,
input [9:0] Pix_23,
input [9:0] Pix_24,
input [9:0] Pix_25,
input [9:0] Pix_26,
input [9:0] Pix_27,
input [9:0] Pix_28,
input [9:0] Pix_29,
input [9:0] Pix_30,
input [9:0] Pix_31,
input [9:0] Pix_32,
input [9:0] Pix_33,
input [9:0] Pix_34,
input [9:0] Pix_35,
input [9:0] Pix_36,
input [9:0] Pix_37,
input [9:0] Pix_38,
input [9:0] Pix_39,
input [9:0] Pix_40,
input [9:0] Pix_41,
input [9:0] Pix_42,
input [9:0] Pix_43,
input [9:0] Pix_44,
input [9:0] Pix_45,
input [9:0] Pix_46,
input [9:0] Pix_47,
input [9:0] Pix_48,
input [9:0] Pix_49,
input [9:0] Pix_50,
input [9:0] Pix_51,
input [9:0] Pix_52,
input [9:0] Pix_53,
input [9:0] Pix_54,
input [9:0] Pix_55,
input [9:0] Pix_56,
input [9:0] Pix_57,
input [9:0] Pix_58,
input [9:0] Pix_59,
input [9:0] Pix_60,
input [9:0] Pix_61,
input [9:0] Pix_62,
input [9:0] Pix_63,
input [9:0] Pix_64,
input [9:0] Pix_65,
input [9:0] Pix_66,
input [9:0] Pix_67,
input [9:0] Pix_68,
input [9:0] Pix_69,
input [9:0] Pix_70,
input [9:0] Pix_71,
input [9:0] Pix_72,
input [9:0] Pix_73,
input [9:0] Pix_74,
input [9:0] Pix_75,
input [9:0] Pix_76,
input [9:0] Pix_77,
input [9:0] Pix_78,
input [9:0] Pix_79,
input [9:0] Pix_80,
input [9:0] Pix_81,
input [9:0] Pix_82,
input [9:0] Pix_83,
input [9:0] Pix_84,
input [9:0] Pix_85,
input [9:0] Pix_86,
input [9:0] Pix_87,
input [9:0] Pix_88,
input [9:0] Pix_89,
input [9:0] Pix_90,
input [9:0] Pix_91,
input [9:0] Pix_92,
input [9:0] Pix_93,
input [9:0] Pix_94,
input [9:0] Pix_95,
input [9:0] Pix_96,
input [9:0] Pix_97,
input [9:0] Pix_98,
input [9:0] Pix_99,
input [9:0] Pix_100,
input [9:0] Pix_101,
input [9:0] Pix_102,
input [9:0] Pix_103,
input [9:0] Pix_104,
input [9:0] Pix_105,
input [9:0] Pix_106,
input [9:0] Pix_107,
input [9:0] Pix_108,
input [9:0] Pix_109,
input [9:0] Pix_110,
input [9:0] Pix_111,
input [9:0] Pix_112,
input [9:0] Pix_113,
input [9:0] Pix_114,
input [9:0] Pix_115,
input [9:0] Pix_116,
input [9:0] Pix_117,
input [9:0] Pix_118,
input [9:0] Pix_119,
input [9:0] Pix_120,
input [9:0] Pix_121,
input [9:0] Pix_122,
input [9:0] Pix_123,
input [9:0] Pix_124,
input [9:0] Pix_125,
input [9:0] Pix_126,
input [9:0] Pix_127,
input [9:0] Pix_128,
input [9:0] Pix_129,
input [9:0] Pix_130,
input [9:0] Pix_131,
input [9:0] Pix_132,
input [9:0] Pix_133,
input [9:0] Pix_134,
input [9:0] Pix_135,
input [9:0] Pix_136,
input [9:0] Pix_137,
input [9:0] Pix_138,
input [9:0] Pix_139,
input [9:0] Pix_140,
input [9:0] Pix_141,
input [9:0] Pix_142,
input [9:0] Pix_143,
input [9:0] Pix_144,
input [9:0] Pix_145,
input [9:0] Pix_146,
input [9:0] Pix_147,
input [9:0] Pix_148,
input [9:0] Pix_149,
input [9:0] Pix_150,
input [9:0] Pix_151,
input [9:0] Pix_152,
input [9:0] Pix_153,
input [9:0] Pix_154,
input [9:0] Pix_155,
input [9:0] Pix_156,
input [9:0] Pix_157,
input [9:0] Pix_158,
input [9:0] Pix_159,
input [9:0] Pix_160,
input [9:0] Pix_161,
input [9:0] Pix_162,
input [9:0] Pix_163,
input [9:0] Pix_164,
input [9:0] Pix_165,
input [9:0] Pix_166,
input [9:0] Pix_167,
input [9:0] Pix_168,
input [9:0] Pix_169,
input [9:0] Pix_170,
input [9:0] Pix_171,
input [9:0] Pix_172,
input [9:0] Pix_173,
input [9:0] Pix_174,
input [9:0] Pix_175,
input [9:0] Pix_176,
input [9:0] Pix_177,
input [9:0] Pix_178,
input [9:0] Pix_179,
input [9:0] Pix_180,
input [9:0] Pix_181,
input [9:0] Pix_182,
input [9:0] Pix_183,
input [9:0] Pix_184,
input [9:0] Pix_185,
input [9:0] Pix_186,
input [9:0] Pix_187,
input [9:0] Pix_188,
input [9:0] Pix_189,
input [9:0] Pix_190,
input [9:0] Pix_191,
input [9:0] Pix_192,
input [9:0] Pix_193,
input [9:0] Pix_194,
input [9:0] Pix_195,
input [9:0] Pix_196,
input [9:0] Pix_197,
input [9:0] Pix_198,
input [9:0] Pix_199,
input [9:0] Pix_200,
input [9:0] Pix_201,
input [9:0] Pix_202,
input [9:0] Pix_203,
input [9:0] Pix_204,
input [9:0] Pix_205,
input [9:0] Pix_206,
input [9:0] Pix_207,
input [9:0] Pix_208,
input [9:0] Pix_209,
input [9:0] Pix_210,
input [9:0] Pix_211,
input [9:0] Pix_212,
input [9:0] Pix_213,
input [9:0] Pix_214,
input [9:0] Pix_215,
input [9:0] Pix_216,
input [9:0] Pix_217,
input [9:0] Pix_218,
input [9:0] Pix_219,
input [9:0] Pix_220,
input [9:0] Pix_221,
input [9:0] Pix_222,
input [9:0] Pix_223,
input [9:0] Pix_224,
input [9:0] Pix_225,
input [9:0] Pix_226,
input [9:0] Pix_227,
input [9:0] Pix_228,
input [9:0] Pix_229,
input [9:0] Pix_230,
input [9:0] Pix_231,
input [9:0] Pix_232,
input [9:0] Pix_233,
input [9:0] Pix_234,
input [9:0] Pix_235,
input [9:0] Pix_236,
input [9:0] Pix_237,
input [9:0] Pix_238,
input [9:0] Pix_239,
input [9:0] Pix_240,
input [9:0] Pix_241,
input [9:0] Pix_242,
input [9:0] Pix_243,
input [9:0] Pix_244,
input [9:0] Pix_245,
input [9:0] Pix_246,
input [9:0] Pix_247,
input [9:0] Pix_248,
input [9:0] Pix_249,
input [9:0] Pix_250,
input [9:0] Pix_251,
input [9:0] Pix_252,
input [9:0] Pix_253,
input [9:0] Pix_254,
input [9:0] Pix_255,
input [9:0] Pix_256,
input [9:0] Pix_257,
input [9:0] Pix_258,
input [9:0] Pix_259,
input [9:0] Pix_260,
input [9:0] Pix_261,
input [9:0] Pix_262,
input [9:0] Pix_263,
input [9:0] Pix_264,
input [9:0] Pix_265,
input [9:0] Pix_266,
input [9:0] Pix_267,
input [9:0] Pix_268,
input [9:0] Pix_269,
input [9:0] Pix_270,
input [9:0] Pix_271,
input [9:0] Pix_272,
input [9:0] Pix_273,
input [9:0] Pix_274,
input [9:0] Pix_275,
input [9:0] Pix_276,
input [9:0] Pix_277,
input [9:0] Pix_278,
input [9:0] Pix_279,
input [9:0] Pix_280,
input [9:0] Pix_281,
input [9:0] Pix_282,
input [9:0] Pix_283,
input [9:0] Pix_284,
input [9:0] Pix_285,
input [9:0] Pix_286,
input [9:0] Pix_287,
input [9:0] Pix_288,
input [9:0] Pix_289,
input [9:0] Pix_290,
input [9:0] Pix_291,
input [9:0] Pix_292,
input [9:0] Pix_293,
input [9:0] Pix_294,
input [9:0] Pix_295,
input [9:0] Pix_296,
input [9:0] Pix_297,
input [9:0] Pix_298,
input [9:0] Pix_299,
input [9:0] Pix_300,
input [9:0] Pix_301,
input [9:0] Pix_302,
input [9:0] Pix_303,
input [9:0] Pix_304,
input [9:0] Pix_305,
input [9:0] Pix_306,
input [9:0] Pix_307,
input [9:0] Pix_308,
input [9:0] Pix_309,
input [9:0] Pix_310,
input [9:0] Pix_311,
input [9:0] Pix_312,
input [9:0] Pix_313,
input [9:0] Pix_314,
input [9:0] Pix_315,
input [9:0] Pix_316,
input [9:0] Pix_317,
input [9:0] Pix_318,
input [9:0] Pix_319,
input [9:0] Pix_320,
input [9:0] Pix_321,
input [9:0] Pix_322,
input [9:0] Pix_323,
input [9:0] Pix_324,
input [9:0] Pix_325,
input [9:0] Pix_326,
input [9:0] Pix_327,
input [9:0] Pix_328,
input [9:0] Pix_329,
input [9:0] Pix_330,
input [9:0] Pix_331,
input [9:0] Pix_332,
input [9:0] Pix_333,
input [9:0] Pix_334,
input [9:0] Pix_335,
input [9:0] Pix_336,
input [9:0] Pix_337,
input [9:0] Pix_338,
input [9:0] Pix_339,
input [9:0] Pix_340,
input [9:0] Pix_341,
input [9:0] Pix_342,
input [9:0] Pix_343,
input [9:0] Pix_344,
input [9:0] Pix_345,
input [9:0] Pix_346,
input [9:0] Pix_347,
input [9:0] Pix_348,
input [9:0] Pix_349,
input [9:0] Pix_350,
input [9:0] Pix_351,
input [9:0] Pix_352,
input [9:0] Pix_353,
input [9:0] Pix_354,
input [9:0] Pix_355,
input [9:0] Pix_356,
input [9:0] Pix_357,
input [9:0] Pix_358,
input [9:0] Pix_359,
input [9:0] Pix_360,
input [9:0] Pix_361,
input [9:0] Pix_362,
input [9:0] Pix_363,
input [9:0] Pix_364,
input [9:0] Pix_365,
input [9:0] Pix_366,
input [9:0] Pix_367,
input [9:0] Pix_368,
input [9:0] Pix_369,
input [9:0] Pix_370,
input [9:0] Pix_371,
input [9:0] Pix_372,
input [9:0] Pix_373,
input [9:0] Pix_374,
input [9:0] Pix_375,
input [9:0] Pix_376,
input [9:0] Pix_377,
input [9:0] Pix_378,
input [9:0] Pix_379,
input [9:0] Pix_380,
input [9:0] Pix_381,
input [9:0] Pix_382,
input [9:0] Pix_383,
input [9:0] Pix_384,
input [9:0] Pix_385,
input [9:0] Pix_386,
input [9:0] Pix_387,
input [9:0] Pix_388,
input [9:0] Pix_389,
input [9:0] Pix_390,
input [9:0] Pix_391,
input [9:0] Pix_392,
input [9:0] Pix_393,
input [9:0] Pix_394,
input [9:0] Pix_395,
input [9:0] Pix_396,
input [9:0] Pix_397,
input [9:0] Pix_398,
input [9:0] Pix_399,
input [9:0] Pix_400,
input [9:0] Pix_401,
input [9:0] Pix_402,
input [9:0] Pix_403,
input [9:0] Pix_404,
input [9:0] Pix_405,
input [9:0] Pix_406,
input [9:0] Pix_407,
input [9:0] Pix_408,
input [9:0] Pix_409,
input [9:0] Pix_410,
input [9:0] Pix_411,
input [9:0] Pix_412,
input [9:0] Pix_413,
input [9:0] Pix_414,
input [9:0] Pix_415,
input [9:0] Pix_416,
input [9:0] Pix_417,
input [9:0] Pix_418,
input [9:0] Pix_419,
input [9:0] Pix_420,
input [9:0] Pix_421,
input [9:0] Pix_422,
input [9:0] Pix_423,
input [9:0] Pix_424,
input [9:0] Pix_425,
input [9:0] Pix_426,
input [9:0] Pix_427,
input [9:0] Pix_428,
input [9:0] Pix_429,
input [9:0] Pix_430,
input [9:0] Pix_431,
input [9:0] Pix_432,
input [9:0] Pix_433,
input [9:0] Pix_434,
input [9:0] Pix_435,
input [9:0] Pix_436,
input [9:0] Pix_437,
input [9:0] Pix_438,
input [9:0] Pix_439,
input [9:0] Pix_440,
input [9:0] Pix_441,
input [9:0] Pix_442,
input [9:0] Pix_443,
input [9:0] Pix_444,
input [9:0] Pix_445,
input [9:0] Pix_446,
input [9:0] Pix_447,
input [9:0] Pix_448,
input [9:0] Pix_449,
input [9:0] Pix_450,
input [9:0] Pix_451,
input [9:0] Pix_452,
input [9:0] Pix_453,
input [9:0] Pix_454,
input [9:0] Pix_455,
input [9:0] Pix_456,
input [9:0] Pix_457,
input [9:0] Pix_458,
input [9:0] Pix_459,
input [9:0] Pix_460,
input [9:0] Pix_461,
input [9:0] Pix_462,
input [9:0] Pix_463,
input [9:0] Pix_464,
input [9:0] Pix_465,
input [9:0] Pix_466,
input [9:0] Pix_467,
input [9:0] Pix_468,
input [9:0] Pix_469,
input [9:0] Pix_470,
input [9:0] Pix_471,
input [9:0] Pix_472,
input [9:0] Pix_473,
input [9:0] Pix_474,
input [9:0] Pix_475,
input [9:0] Pix_476,
input [9:0] Pix_477,
input [9:0] Pix_478,
input [9:0] Pix_479,
input [9:0] Pix_480,
input [9:0] Pix_481,
input [9:0] Pix_482,
input [9:0] Pix_483,
input [9:0] Pix_484,
input [9:0] Pix_485,
input [9:0] Pix_486,
input [9:0] Pix_487,
input [9:0] Pix_488,
input [9:0] Pix_489,
input [9:0] Pix_490,
input [9:0] Pix_491,
input [9:0] Pix_492,
input [9:0] Pix_493,
input [9:0] Pix_494,
input [9:0] Pix_495,
input [9:0] Pix_496,
input [9:0] Pix_497,
input [9:0] Pix_498,
input [9:0] Pix_499,
input [9:0] Pix_500,
input [9:0] Pix_501,
input [9:0] Pix_502,
input [9:0] Pix_503,
input [9:0] Pix_504,
input [9:0] Pix_505,
input [9:0] Pix_506,
input [9:0] Pix_507,
input [9:0] Pix_508,
input [9:0] Pix_509,
input [9:0] Pix_510,
input [9:0] Pix_511,
input [9:0] Pix_512,
input [9:0] Pix_513,
input [9:0] Pix_514,
input [9:0] Pix_515,
input [9:0] Pix_516,
input [9:0] Pix_517,
input [9:0] Pix_518,
input [9:0] Pix_519,
input [9:0] Pix_520,
input [9:0] Pix_521,
input [9:0] Pix_522,
input [9:0] Pix_523,
input [9:0] Pix_524,
input [9:0] Pix_525,
input [9:0] Pix_526,
input [9:0] Pix_527,
input [9:0] Pix_528,
input [9:0] Pix_529,
input [9:0] Pix_530,
input [9:0] Pix_531,
input [9:0] Pix_532,
input [9:0] Pix_533,
input [9:0] Pix_534,
input [9:0] Pix_535,
input [9:0] Pix_536,
input [9:0] Pix_537,
input [9:0] Pix_538,
input [9:0] Pix_539,
input [9:0] Pix_540,
input [9:0] Pix_541,
input [9:0] Pix_542,
input [9:0] Pix_543,
input [9:0] Pix_544,
input [9:0] Pix_545,
input [9:0] Pix_546,
input [9:0] Pix_547,
input [9:0] Pix_548,
input [9:0] Pix_549,
input [9:0] Pix_550,
input [9:0] Pix_551,
input [9:0] Pix_552,
input [9:0] Pix_553,
input [9:0] Pix_554,
input [9:0] Pix_555,
input [9:0] Pix_556,
input [9:0] Pix_557,
input [9:0] Pix_558,
input [9:0] Pix_559,
input [9:0] Pix_560,
input [9:0] Pix_561,
input [9:0] Pix_562,
input [9:0] Pix_563,
input [9:0] Pix_564,
input [9:0] Pix_565,
input [9:0] Pix_566,
input [9:0] Pix_567,
input [9:0] Pix_568,
input [9:0] Pix_569,
input [9:0] Pix_570,
input [9:0] Pix_571,
input [9:0] Pix_572,
input [9:0] Pix_573,
input [9:0] Pix_574,
input [9:0] Pix_575,
input [9:0] Pix_576,
input [9:0] Pix_577,
input [9:0] Pix_578,
input [9:0] Pix_579,
input [9:0] Pix_580,
input [9:0] Pix_581,
input [9:0] Pix_582,
input [9:0] Pix_583,
input [9:0] Pix_584,
input [9:0] Pix_585,
input [9:0] Pix_586,
input [9:0] Pix_587,
input [9:0] Pix_588,
input [9:0] Pix_589,
input [9:0] Pix_590,
input [9:0] Pix_591,
input [9:0] Pix_592,
input [9:0] Pix_593,
input [9:0] Pix_594,
input [9:0] Pix_595,
input [9:0] Pix_596,
input [9:0] Pix_597,
input [9:0] Pix_598,
input [9:0] Pix_599,
input [9:0] Pix_600,
input [9:0] Pix_601,
input [9:0] Pix_602,
input [9:0] Pix_603,
input [9:0] Pix_604,
input [9:0] Pix_605,
input [9:0] Pix_606,
input [9:0] Pix_607,
input [9:0] Pix_608,
input [9:0] Pix_609,
input [9:0] Pix_610,
input [9:0] Pix_611,
input [9:0] Pix_612,
input [9:0] Pix_613,
input [9:0] Pix_614,
input [9:0] Pix_615,
input [9:0] Pix_616,
input [9:0] Pix_617,
input [9:0] Pix_618,
input [9:0] Pix_619,
input [9:0] Pix_620,
input [9:0] Pix_621,
input [9:0] Pix_622,
input [9:0] Pix_623,
input [9:0] Pix_624,
input [9:0] Pix_625,
input [9:0] Pix_626,
input [9:0] Pix_627,
input [9:0] Pix_628,
input [9:0] Pix_629,
input [9:0] Pix_630,
input [9:0] Pix_631,
input [9:0] Pix_632,
input [9:0] Pix_633,
input [9:0] Pix_634,
input [9:0] Pix_635,
input [9:0] Pix_636,
input [9:0] Pix_637,
input [9:0] Pix_638,
input [9:0] Pix_639,
input [9:0] Pix_640,
input [9:0] Pix_641,
input [9:0] Pix_642,
input [9:0] Pix_643,
input [9:0] Pix_644,
input [9:0] Pix_645,
input [9:0] Pix_646,
input [9:0] Pix_647,
input [9:0] Pix_648,
input [9:0] Pix_649,
input [9:0] Pix_650,
input [9:0] Pix_651,
input [9:0] Pix_652,
input [9:0] Pix_653,
input [9:0] Pix_654,
input [9:0] Pix_655,
input [9:0] Pix_656,
input [9:0] Pix_657,
input [9:0] Pix_658,
input [9:0] Pix_659,
input [9:0] Pix_660,
input [9:0] Pix_661,
input [9:0] Pix_662,
input [9:0] Pix_663,
input [9:0] Pix_664,
input [9:0] Pix_665,
input [9:0] Pix_666,
input [9:0] Pix_667,
input [9:0] Pix_668,
input [9:0] Pix_669,
input [9:0] Pix_670,
input [9:0] Pix_671,
input [9:0] Pix_672,
input [9:0] Pix_673,
input [9:0] Pix_674,
input [9:0] Pix_675,
input [9:0] Pix_676,
input [9:0] Pix_677,
input [9:0] Pix_678,
input [9:0] Pix_679,
input [9:0] Pix_680,
input [9:0] Pix_681,
input [9:0] Pix_682,
input [9:0] Pix_683,
input [9:0] Pix_684,
input [9:0] Pix_685,
input [9:0] Pix_686,
input [9:0] Pix_687,
input [9:0] Pix_688,
input [9:0] Pix_689,
input [9:0] Pix_690,
input [9:0] Pix_691,
input [9:0] Pix_692,
input [9:0] Pix_693,
input [9:0] Pix_694,
input [9:0] Pix_695,
input [9:0] Pix_696,
input [9:0] Pix_697,
input [9:0] Pix_698,
input [9:0] Pix_699,
input [9:0] Pix_700,
input [9:0] Pix_701,
input [9:0] Pix_702,
input [9:0] Pix_703,
input [9:0] Pix_704,
input [9:0] Pix_705,
input [9:0] Pix_706,
input [9:0] Pix_707,
input [9:0] Pix_708,
input [9:0] Pix_709,
input [9:0] Pix_710,
input [9:0] Pix_711,
input [9:0] Pix_712,
input [9:0] Pix_713,
input [9:0] Pix_714,
input [9:0] Pix_715,
input [9:0] Pix_716,
input [9:0] Pix_717,
input [9:0] Pix_718,
input [9:0] Pix_719,
input [9:0] Pix_720,
input [9:0] Pix_721,
input [9:0] Pix_722,
input [9:0] Pix_723,
input [9:0] Pix_724,
input [9:0] Pix_725,
input [9:0] Pix_726,
input [9:0] Pix_727,
input [9:0] Pix_728,
input [9:0] Pix_729,
input [9:0] Pix_730,
input [9:0] Pix_731,
input [9:0] Pix_732,
input [9:0] Pix_733,
input [9:0] Pix_734,
input [9:0] Pix_735,
input [9:0] Pix_736,
input [9:0] Pix_737,
input [9:0] Pix_738,
input [9:0] Pix_739,
input [9:0] Pix_740,
input [9:0] Pix_741,
input [9:0] Pix_742,
input [9:0] Pix_743,
input [9:0] Pix_744,
input [9:0] Pix_745,
input [9:0] Pix_746,
input [9:0] Pix_747,
input [9:0] Pix_748,
input [9:0] Pix_749,
input [9:0] Pix_750,
input [9:0] Pix_751,
input [9:0] Pix_752,
input [9:0] Pix_753,
input [9:0] Pix_754,
input [9:0] Pix_755,
input [9:0] Pix_756,
input [9:0] Pix_757,
input [9:0] Pix_758,
input [9:0] Pix_759,
input [9:0] Pix_760,
input [9:0] Pix_761,
input [9:0] Pix_762,
input [9:0] Pix_763,
input [9:0] Pix_764,
input [9:0] Pix_765,
input [9:0] Pix_766,
input [9:0] Pix_767,
input [9:0] Pix_768,
input [9:0] Pix_769,
input [9:0] Pix_770,
input [9:0] Pix_771,
input [9:0] Pix_772,
input [9:0] Pix_773,
input [9:0] Pix_774,
input [9:0] Pix_775,
input [9:0] Pix_776,
input [9:0] Pix_777,
input [9:0] Pix_778,
input [9:0] Pix_779,
input [9:0] Pix_780,
input [9:0] Pix_781,
input [9:0] Pix_782,
input [9:0] Pix_783,
input [9:0] Pix_784,
output [3:0] Image_Number,
output Output_Valid
);

reg[9:0] PixelsStore[0:784];
reg[18:0] WeightsStore0[0:784];
reg[18:0] WeightsStore1[0:784];
reg[18:0] WeightsStore2[0:784];
reg[18:0] WeightsStore3[0:784];
reg[18:0] WeightsStore4[0:784];
reg[18:0] WeightsStore5[0:784];
reg[18:0] WeightsStore6[0:784];
reg[18:0] WeightsStore7[0:784];
reg[18:0] WeightsStore8[0:784];
reg[18:0] WeightsStore9[0:784];
reg[31:0] switchCounter;
reg ready;
reg internalReset
;wire[259:0] value;

assign Output_Valid = ready;

DotProduct784 DP0(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore0[0]),
	.Weight1(WeightsStore0[1]),
	.Weight2(WeightsStore0[2]),
	.Weight3(WeightsStore0[3]),
	.Weight4(WeightsStore0[4]),
	.Weight5(WeightsStore0[5]),
	.Weight6(WeightsStore0[6]),
	.Weight7(WeightsStore0[7]),
	.Weight8(WeightsStore0[8]),
	.Weight9(WeightsStore0[9]),
	.Weight10(WeightsStore0[10]),
	.Weight11(WeightsStore0[11]),
	.Weight12(WeightsStore0[12]),
	.Weight13(WeightsStore0[13]),
	.Weight14(WeightsStore0[14]),
	.Weight15(WeightsStore0[15]),
	.Weight16(WeightsStore0[16]),
	.Weight17(WeightsStore0[17]),
	.Weight18(WeightsStore0[18]),
	.Weight19(WeightsStore0[19]),
	.Weight20(WeightsStore0[20]),
	.Weight21(WeightsStore0[21]),
	.Weight22(WeightsStore0[22]),
	.Weight23(WeightsStore0[23]),
	.Weight24(WeightsStore0[24]),
	.Weight25(WeightsStore0[25]),
	.Weight26(WeightsStore0[26]),
	.Weight27(WeightsStore0[27]),
	.WeightBias(WeightsStore0[784]),
	.value(value[25:0])
	);
DotProduct784 DP1(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore1[0]),
	.Weight1(WeightsStore1[1]),
	.Weight2(WeightsStore1[2]),
	.Weight3(WeightsStore1[3]),
	.Weight4(WeightsStore1[4]),
	.Weight5(WeightsStore1[5]),
	.Weight6(WeightsStore1[6]),
	.Weight7(WeightsStore1[7]),
	.Weight8(WeightsStore1[8]),
	.Weight9(WeightsStore1[9]),
	.Weight10(WeightsStore1[10]),
	.Weight11(WeightsStore1[11]),
	.Weight12(WeightsStore1[12]),
	.Weight13(WeightsStore1[13]),
	.Weight14(WeightsStore1[14]),
	.Weight15(WeightsStore1[15]),
	.Weight16(WeightsStore1[16]),
	.Weight17(WeightsStore1[17]),
	.Weight18(WeightsStore1[18]),
	.Weight19(WeightsStore1[19]),
	.Weight20(WeightsStore1[20]),
	.Weight21(WeightsStore1[21]),
	.Weight22(WeightsStore1[22]),
	.Weight23(WeightsStore1[23]),
	.Weight24(WeightsStore1[24]),
	.Weight25(WeightsStore1[25]),
	.Weight26(WeightsStore1[26]),
	.Weight27(WeightsStore1[27]),
	.WeightBias(WeightsStore1[784]),
	.value(value[51:26])
	);
DotProduct784 DP2(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore2[0]),
	.Weight1(WeightsStore2[1]),
	.Weight2(WeightsStore2[2]),
	.Weight3(WeightsStore2[3]),
	.Weight4(WeightsStore2[4]),
	.Weight5(WeightsStore2[5]),
	.Weight6(WeightsStore2[6]),
	.Weight7(WeightsStore2[7]),
	.Weight8(WeightsStore2[8]),
	.Weight9(WeightsStore2[9]),
	.Weight10(WeightsStore2[10]),
	.Weight11(WeightsStore2[11]),
	.Weight12(WeightsStore2[12]),
	.Weight13(WeightsStore2[13]),
	.Weight14(WeightsStore2[14]),
	.Weight15(WeightsStore2[15]),
	.Weight16(WeightsStore2[16]),
	.Weight17(WeightsStore2[17]),
	.Weight18(WeightsStore2[18]),
	.Weight19(WeightsStore2[19]),
	.Weight20(WeightsStore2[20]),
	.Weight21(WeightsStore2[21]),
	.Weight22(WeightsStore2[22]),
	.Weight23(WeightsStore2[23]),
	.Weight24(WeightsStore2[24]),
	.Weight25(WeightsStore2[25]),
	.Weight26(WeightsStore2[26]),
	.Weight27(WeightsStore2[27]),
	.WeightBias(WeightsStore2[784]),
	.value(value[77:52])
	);
DotProduct784 DP3(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore3[0]),
	.Weight1(WeightsStore3[1]),
	.Weight2(WeightsStore3[2]),
	.Weight3(WeightsStore3[3]),
	.Weight4(WeightsStore3[4]),
	.Weight5(WeightsStore3[5]),
	.Weight6(WeightsStore3[6]),
	.Weight7(WeightsStore3[7]),
	.Weight8(WeightsStore3[8]),
	.Weight9(WeightsStore3[9]),
	.Weight10(WeightsStore3[10]),
	.Weight11(WeightsStore3[11]),
	.Weight12(WeightsStore3[12]),
	.Weight13(WeightsStore3[13]),
	.Weight14(WeightsStore3[14]),
	.Weight15(WeightsStore3[15]),
	.Weight16(WeightsStore3[16]),
	.Weight17(WeightsStore3[17]),
	.Weight18(WeightsStore3[18]),
	.Weight19(WeightsStore3[19]),
	.Weight20(WeightsStore3[20]),
	.Weight21(WeightsStore3[21]),
	.Weight22(WeightsStore3[22]),
	.Weight23(WeightsStore3[23]),
	.Weight24(WeightsStore3[24]),
	.Weight25(WeightsStore3[25]),
	.Weight26(WeightsStore3[26]),
	.Weight27(WeightsStore3[27]),
	.WeightBias(WeightsStore3[784]),
	.value(value[103:78])
	);
DotProduct784 DP4(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore4[0]),
	.Weight1(WeightsStore4[1]),
	.Weight2(WeightsStore4[2]),
	.Weight3(WeightsStore4[3]),
	.Weight4(WeightsStore4[4]),
	.Weight5(WeightsStore4[5]),
	.Weight6(WeightsStore4[6]),
	.Weight7(WeightsStore4[7]),
	.Weight8(WeightsStore4[8]),
	.Weight9(WeightsStore4[9]),
	.Weight10(WeightsStore4[10]),
	.Weight11(WeightsStore4[11]),
	.Weight12(WeightsStore4[12]),
	.Weight13(WeightsStore4[13]),
	.Weight14(WeightsStore4[14]),
	.Weight15(WeightsStore4[15]),
	.Weight16(WeightsStore4[16]),
	.Weight17(WeightsStore4[17]),
	.Weight18(WeightsStore4[18]),
	.Weight19(WeightsStore4[19]),
	.Weight20(WeightsStore4[20]),
	.Weight21(WeightsStore4[21]),
	.Weight22(WeightsStore4[22]),
	.Weight23(WeightsStore4[23]),
	.Weight24(WeightsStore4[24]),
	.Weight25(WeightsStore4[25]),
	.Weight26(WeightsStore4[26]),
	.Weight27(WeightsStore4[27]),
	.WeightBias(WeightsStore4[784]),
	.value(value[129:104])
	);
DotProduct784 DP5(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore5[0]),
	.Weight1(WeightsStore5[1]),
	.Weight2(WeightsStore5[2]),
	.Weight3(WeightsStore5[3]),
	.Weight4(WeightsStore5[4]),
	.Weight5(WeightsStore5[5]),
	.Weight6(WeightsStore5[6]),
	.Weight7(WeightsStore5[7]),
	.Weight8(WeightsStore5[8]),
	.Weight9(WeightsStore5[9]),
	.Weight10(WeightsStore5[10]),
	.Weight11(WeightsStore5[11]),
	.Weight12(WeightsStore5[12]),
	.Weight13(WeightsStore5[13]),
	.Weight14(WeightsStore5[14]),
	.Weight15(WeightsStore5[15]),
	.Weight16(WeightsStore5[16]),
	.Weight17(WeightsStore5[17]),
	.Weight18(WeightsStore5[18]),
	.Weight19(WeightsStore5[19]),
	.Weight20(WeightsStore5[20]),
	.Weight21(WeightsStore5[21]),
	.Weight22(WeightsStore5[22]),
	.Weight23(WeightsStore5[23]),
	.Weight24(WeightsStore5[24]),
	.Weight25(WeightsStore5[25]),
	.Weight26(WeightsStore5[26]),
	.Weight27(WeightsStore5[27]),
	.WeightBias(WeightsStore5[784]),
	.value(value[155:130])
	);
DotProduct784 DP6(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore6[0]),
	.Weight1(WeightsStore6[1]),
	.Weight2(WeightsStore6[2]),
	.Weight3(WeightsStore6[3]),
	.Weight4(WeightsStore6[4]),
	.Weight5(WeightsStore6[5]),
	.Weight6(WeightsStore6[6]),
	.Weight7(WeightsStore6[7]),
	.Weight8(WeightsStore6[8]),
	.Weight9(WeightsStore6[9]),
	.Weight10(WeightsStore6[10]),
	.Weight11(WeightsStore6[11]),
	.Weight12(WeightsStore6[12]),
	.Weight13(WeightsStore6[13]),
	.Weight14(WeightsStore6[14]),
	.Weight15(WeightsStore6[15]),
	.Weight16(WeightsStore6[16]),
	.Weight17(WeightsStore6[17]),
	.Weight18(WeightsStore6[18]),
	.Weight19(WeightsStore6[19]),
	.Weight20(WeightsStore6[20]),
	.Weight21(WeightsStore6[21]),
	.Weight22(WeightsStore6[22]),
	.Weight23(WeightsStore6[23]),
	.Weight24(WeightsStore6[24]),
	.Weight25(WeightsStore6[25]),
	.Weight26(WeightsStore6[26]),
	.Weight27(WeightsStore6[27]),
	.WeightBias(WeightsStore6[784]),
	.value(value[181:156])
	);
DotProduct784 DP7(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore7[0]),
	.Weight1(WeightsStore7[1]),
	.Weight2(WeightsStore7[2]),
	.Weight3(WeightsStore7[3]),
	.Weight4(WeightsStore7[4]),
	.Weight5(WeightsStore7[5]),
	.Weight6(WeightsStore7[6]),
	.Weight7(WeightsStore7[7]),
	.Weight8(WeightsStore7[8]),
	.Weight9(WeightsStore7[9]),
	.Weight10(WeightsStore7[10]),
	.Weight11(WeightsStore7[11]),
	.Weight12(WeightsStore7[12]),
	.Weight13(WeightsStore7[13]),
	.Weight14(WeightsStore7[14]),
	.Weight15(WeightsStore7[15]),
	.Weight16(WeightsStore7[16]),
	.Weight17(WeightsStore7[17]),
	.Weight18(WeightsStore7[18]),
	.Weight19(WeightsStore7[19]),
	.Weight20(WeightsStore7[20]),
	.Weight21(WeightsStore7[21]),
	.Weight22(WeightsStore7[22]),
	.Weight23(WeightsStore7[23]),
	.Weight24(WeightsStore7[24]),
	.Weight25(WeightsStore7[25]),
	.Weight26(WeightsStore7[26]),
	.Weight27(WeightsStore7[27]),
	.WeightBias(WeightsStore7[784]),
	.value(value[207:182])
	);
DotProduct784 DP8(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore8[0]),
	.Weight1(WeightsStore8[1]),
	.Weight2(WeightsStore8[2]),
	.Weight3(WeightsStore8[3]),
	.Weight4(WeightsStore8[4]),
	.Weight5(WeightsStore8[5]),
	.Weight6(WeightsStore8[6]),
	.Weight7(WeightsStore8[7]),
	.Weight8(WeightsStore8[8]),
	.Weight9(WeightsStore8[9]),
	.Weight10(WeightsStore8[10]),
	.Weight11(WeightsStore8[11]),
	.Weight12(WeightsStore8[12]),
	.Weight13(WeightsStore8[13]),
	.Weight14(WeightsStore8[14]),
	.Weight15(WeightsStore8[15]),
	.Weight16(WeightsStore8[16]),
	.Weight17(WeightsStore8[17]),
	.Weight18(WeightsStore8[18]),
	.Weight19(WeightsStore8[19]),
	.Weight20(WeightsStore8[20]),
	.Weight21(WeightsStore8[21]),
	.Weight22(WeightsStore8[22]),
	.Weight23(WeightsStore8[23]),
	.Weight24(WeightsStore8[24]),
	.Weight25(WeightsStore8[25]),
	.Weight26(WeightsStore8[26]),
	.Weight27(WeightsStore8[27]),
	.WeightBias(WeightsStore8[784]),
	.value(value[233:208])
	);
DotProduct784 DP9(.clk(clk),
	.GlobalReset(internalReset),
	.Pixel0(PixelsStore[0]),
	.Pixel1(PixelsStore[1]),
	.Pixel2(PixelsStore[2]),
	.Pixel3(PixelsStore[3]),
	.Pixel4(PixelsStore[4]),
	.Pixel5(PixelsStore[5]),
	.Pixel6(PixelsStore[6]),
	.Pixel7(PixelsStore[7]),
	.Pixel8(PixelsStore[8]),
	.Pixel9(PixelsStore[9]),
	.Pixel10(PixelsStore[10]),
	.Pixel11(PixelsStore[11]),
	.Pixel12(PixelsStore[12]),
	.Pixel13(PixelsStore[13]),
	.Pixel14(PixelsStore[14]),
	.Pixel15(PixelsStore[15]),
	.Pixel16(PixelsStore[16]),
	.Pixel17(PixelsStore[17]),
	.Pixel18(PixelsStore[18]),
	.Pixel19(PixelsStore[19]),
	.Pixel20(PixelsStore[20]),
	.Pixel21(PixelsStore[21]),
	.Pixel22(PixelsStore[22]),
	.Pixel23(PixelsStore[23]),
	.Pixel24(PixelsStore[24]),
	.Pixel25(PixelsStore[25]),
	.Pixel26(PixelsStore[26]),
	.Pixel27(PixelsStore[27]),
	.Weight0(WeightsStore9[0]),
	.Weight1(WeightsStore9[1]),
	.Weight2(WeightsStore9[2]),
	.Weight3(WeightsStore9[3]),
	.Weight4(WeightsStore9[4]),
	.Weight5(WeightsStore9[5]),
	.Weight6(WeightsStore9[6]),
	.Weight7(WeightsStore9[7]),
	.Weight8(WeightsStore9[8]),
	.Weight9(WeightsStore9[9]),
	.Weight10(WeightsStore9[10]),
	.Weight11(WeightsStore9[11]),
	.Weight12(WeightsStore9[12]),
	.Weight13(WeightsStore9[13]),
	.Weight14(WeightsStore9[14]),
	.Weight15(WeightsStore9[15]),
	.Weight16(WeightsStore9[16]),
	.Weight17(WeightsStore9[17]),
	.Weight18(WeightsStore9[18]),
	.Weight19(WeightsStore9[19]),
	.Weight20(WeightsStore9[20]),
	.Weight21(WeightsStore9[21]),
	.Weight22(WeightsStore9[22]),
	.Weight23(WeightsStore9[23]),
	.Weight24(WeightsStore9[24]),
	.Weight25(WeightsStore9[25]),
	.Weight26(WeightsStore9[26]),
	.Weight27(WeightsStore9[27]),
	.WeightBias(WeightsStore9[784]),
	.value(value[259:234])
	);
Max max(.GlobalReset(internalReset),
	.Num(value),
	.Index(Image_Number)
	);

always@(posedge clk)begin
	if(GlobalReset == 1'b0)begin
		switchCounter <= 32'd0;
		ready <= 1'b0;
		internalReset = 1'b0;
	end
	if(Input_Valid == 1'b1)begin
		switchCounter <= 32'd0;
		ready <= 1'b0;
		internalReset = 1'b0;
	end else begin
		internalReset = 1'b1;
		switchCounter <= switchCounter + 32'd1;
		if(switchCounter == 32'd0)begin
		end else if(switchCounter == 32'd6)begin
		end else if(switchCounter == 32'd13)begin
		end else if(switchCounter == 32'd20)begin
		end else if(switchCounter == 32'd27)begin
		end else if(switchCounter == 32'd34)begin
		end else if(switchCounter == 32'd41)begin
		end else if(switchCounter == 32'd48)begin
		end else if(switchCounter == 32'd55)begin
		end else if(switchCounter == 32'd62)begin
		end else if(switchCounter == 32'd69)begin
		end else if(switchCounter == 32'd76)begin
		end else if(switchCounter == 32'd83)begin
		end else if(switchCounter == 32'd90)begin
		end else if(switchCounter == 32'd97)begin
		end else if(switchCounter == 32'd104)begin
		end else if(switchCounter == 32'd111)begin
		end else if(switchCounter == 32'd118)begin
		end else if(switchCounter == 32'd125)begin
		end else if(switchCounter == 32'd132)begin
		end else if(switchCounter == 32'd139)begin
		end else if(switchCounter == 32'd146)begin
		end else if(switchCounter == 32'd153)begin
		end else if(switchCounter == 32'd160)begin
		end else if(switchCounter == 32'd167)begin
		end else if(switchCounter == 32'd174)begin
		end else if(switchCounter == 32'd181)begin
		end else if(switchCounter == 32'd188)begin
		end else if(switchCounter == 32'd299) begin
			ready <= 1'b1;
			$display("%d %b.%b", switchCounter, value[259:252],value[251:234]);
			$display("%d %b.%b", switchCounter, value[233:226],value[225:208]);
			$display("%d %b.%b", switchCounter, value[207:200],value[199:182]);
			$display("%d %b.%b", switchCounter, value[181:174],value[173:156]);
			$display("%d %b.%b", switchCounter, value[155:148],value[147:130]);
			$display("%d %b.%b", switchCounter, value[129:122],value[121:104]);
			$display("%d %b.%b", switchCounter, value[103:96],value[95:78]);
			$display("%d %b.%b", switchCounter, value[77:70],value[69:52]);
			$display("%d %b.%b", switchCounter, value[51:44],value[43:26]);
			$display("%d %b.%b", switchCounter, value[25:18],value[17:0]);
		end
	end
end
endmodule
